PK   �X�X�,�-�  [    cirkitFile.json�]ێ�6��#�yK%x'�o;�]�k7ƃ���FBʝ���ڬ,�x�������*��P��Pf5�ƌ�$*ƍT���6�կ��f뗿���j����z>��m����U6�=����f��6{�8{�{�;����b��q���ݲ��,��2OSi�da�\�Z��;U�%��y��0Ӻ�\�D�L&J�,�*^&6+r+�-���{;�Zk���>K�si���L2[���)˖��>�?�a�S���m�m)�V������&Yae���Yʘ<*��W�0��0f�4���%9cy^�2���ؖ%/��E�3�Ne�'iZ�ċBƼs9��	\Ǆ����E��<c��&^)�,�K����f̖FXK����36f$�#3�[S��c�F
��c+�Bs�%λ"QRB�EV%�e�^q�KY̩.����p�Uy��>sI�	_qSy�E���p�\*YI�(!E���3��`���,AZ1� Uvo�<��+�Id�t�
W&Ϊ2�l�������uL{�VTD{	˜� \嬀y�0OEY���R��k>�'8L����g��U�}�Z��2+ڈUd�i�rE��E	�"/�k�?��4�`��5�gM�9�������a%k
�$����b�FG��I=��tc�{FMs3�qN{\����c��� ��!Tφ&2}����[y�le���B��v���LTL���<�R���8ȑ~3a�NRIHiGT%�A�7Rb�c��Α�wB�1��4��=#�*�g���nP�J�f����x�(�=�0���%�gE��+p\�B�f	=�0���c�	�HL��(�gb�@�9�{���I<�%xd�'��A�%�ޱ�L���s)%��=H�D,&�����\�Y"A��7	f++E�h��]f��Ҹ���R8i�H ��v#�yRe�v���.�����<_HNT�d=�$�S�/��y�R#U7С�!�zF�+����&h����M�k�3E�ȇ#��6`�I��$��Ai�X�ȇ	���xo�W�v�|gԆ��G=Uަy
��Ka�����Ll��<�,���&�h�
�s������Q���M����&���xJ+�D�s"�yܣ�=?���'b����k{��_�j���3�����8����� M�y�l�if�r�E<}乖ٷ�g��r�@�dN����*���5��T�*���Ț��S���.�����1�`����,c���y�(��=^t%�~*���a�`����ݞ^ح��Ո�6��>	1	9	5��ۣè�nuN0";F��9b���"��vpxDؽ��a���G�ݾ�ح�a]��V��-�a����#��T3���f�ndk)��#ңk�E5�:�v��`R8��@66G�m��a�t����������8pCTF��y���R�S�#��1t�UY�0v�axD��	���a�PᣨC&�/L�%a��MBet`�#�����ʨ��f�g�fV[E�Rc7uU�c�d�x��z���T�$T�iP7x�A/��|�ʢ��S���܌&"���\25<���iޓ�9�l�v��SS�k���fĔ� tʖNe^�$T�tʖNetD�-���L�S�t*z�
:eK�2:��-��(/�-��4��� tʖNe��-�����՘ؔ-�ʸ��l��S�t*�#B�l��S�t*�#B�l�T��.6eK�2/�3�N�ҩ��:t�vxMcS�t*�s�N�ҩL��(^�)�A*�-�ʨ\�)[:�Q��S�t*����S����S�6e;H���S�$ؔ-��4��[5lʖNe|aS�t*�<:eK��&��N����;z�4�����O`>��4�F�l�T.Q�e��s�?c�\����|>�������CV�r�Z/7��ogo�M_�{�z��rسד׮A��O�oDI_Rz��u�$iG���5y�,t�"�;��M ʘ)g�E�gR�Bl��<bk�L_�[�d�:;��/��+7�g$�7�g�zF��cc�Gu��5	�gd���ȼ�<#��7�I�)��]�s����'�6�:f����b�2�:,���	/��+
^f�y�2WE���ke\��R���P"%�=���9*m$�7�g$߷�6a�����'#���sEI>FzF&@))�Hϔ5��%��'�t|��&�AWM��\�l�Pz�h��)���_���NJ�Ŵ.�FI�Sz�0�ᘥ��O�_}���e_����ji��s���bo��{���Sz�) f��G��.b��.b�o��{d�����#Hg��
d�A:����� 6?8,�;�	k^�����i«$c�Y˛�����K��a�L�t��2�CF�fS�MlK��M:�4��}��� 1����#��i�[���%�<��R�w��-�/�|�{����i����1��c`��{l2p�� ����;�K��t�{�Sp�-:ԝ�aO�t��a'!ۖϫ��n���MU��ϫ�Zҁ�~H��9Z��C.RP]�EΒR�r�����M�"Ą������Je^�%��@W�h���It���u$p�C�h��,2te���
@��X�����yI|���2�8(��KPFg�ϣJ����,Aa�G�F���nt�*�ѡ�K�F�.4�"G�L5V+�KO��E,
�E�\�{i�b��D���<�J9d�'�.IA�P�28(��Q4��*֡S��]�7Xt�����E*"ϣ�S��MI��]��E����]w�-��q�E���\w������%�׃;J�g��\4v��kb���������G��G��h��glM��Bt���|JE�T|r*@����W� ����h�Z?�,::���q�[��b��e>;�Y�!���Bv�{_�"��̇I���ς�?������k"���^g��[�UL�� &�ۑ��,(o[	��h��0�}�!L��#&nJ�Ņ���=b^�a\���9s0U�WA�Ux�"q%xUU!��~�9N�?��K ��6��y`���"t�8ԡc�_Jk?��k_�v�kG��f�[S��4�h�NAu=�5����Z�硣�	_���oAya���ܑB��wx�-�I��Ú��$%�B�*"0�0��S�&P	�P+,u�&h�^L�l.QrG����>,My��.�S�{"���,���kQ��E�W�(�m�m�҈�RV������ߔ �2�$�ܥ�D7�����'��*��D7��'� *�HD7�M�nD7��
�QT���!0C<y�v�P�C���w�4fH[��w߄�����-޽%�D��<ܒ�[�pKuo��-ݽe�L��=ܲ�[�p�uo��[i�?J�w��O��ʃ����G��D�Q"�+~	�ʄe��	f�|�2�d�PE��,VO�}��s��_�]�~�/��n�v��!����yZ�V�540J-�6Kc��r:uL� ���p7�֬�'��g����0��4�,�=u�w�}�i��l�~�e�bO�М�6�P���͞�նx��!�S�.t�����|aE��9ȱ���~����s�ڜ8��\H�X,�P��}���Zh���4�S2��T٤�\�(bV��X�2?�@I��mKg����# ���0rnD��N(�~@f&���o[�o�Zz�{�.x#ՂIA�~BŜ˅P�IyZ*��w^WUT�m1�)��V����aU��W��%T'� ���{�Y��D^\pya.�����͇�$b�q��6נ�҅�mZZ/Zf�v�/h��n����Kj���TO���Y-a4�D-�Ҝ�:����	Sl+p4LZB�$��1�&-�Q�
�3��9v�sXC�`��zѢ��K�5����	���O��j�3p��>���������9��m0$��h����q����w@s����<�|�ۿ��V��?]���~^m=�g�}�0C���3����m(����ٙ�+�j���}���|��@�\5�8	�[؆�����QY1����LTnM%�\��Np#�fG
��`� �sq���`L�?X-�����ZS���k��l���U��I
� �' �ե?�g�z�A�?⬃p J�~��ց�|I���3�̾���ܾ�u5�η�}sc��� ����hb�|P��	���%���2}y�n`Ap.A�ϭt�kNY
>P�A����PI**��*����L+�s�0;��][�9�#�P�����q�ZN $T�^HGʷj�;�p|�9ȪQ����]� �q�ȅ��,�s�gA~��PG'�"�S2�����2��=KX��(KPz
!�i���rK@�*�����W������x��;2V4B����'Z"Qi��"1)�T�O��.�C�@ɨ����j��Tl������k�����,��s����:�k��;�x�(���æ�%�K�9�LD��� S�3^P�{x�`ζcB�� 8	��}��Mh��I_���� �^��$��j��b�ǰ�&����
������[�K�5I�Y ]#����s|+���$�2C�푂q5K!rv�D��G �P`�!��9ġ�d�o��Z�f2�k�ZR��.�7_�o����+e����l��<�o���.�JyB�T{]{��4�����:&l�@�h��ę�L9�Q;N� A�C�Ձ�k�#L������oI=0n��?�Kkg)7F��N&X�J�E�����N���1�i��*c
gK����'�Uy�i�c��F�ҧ�S ZS�:����:�.��i�m�~�8��^a[�4��^�`�|��,�c��j̊o���������Y����l���vA�t���ŕCa_cp�7;�Ϫ���w��~�*���}|{�~�K8�\���v�.�_�`��L��y��V����Ϗ���͑�urlu����q��w/��Ci��j�������z�y"
��(�־�<���~��<�^[Y�࠲Rc5x4.�KpuB�!eHh��]�
��0*��-S��y�� ;	�U�A$d�@ne�N%��	ԥ��������;%��]�2Bg	@��C�����TJ�$� L+��K�*+q@��nK��W�|Xb�hm��Kȋ�4S�r
�v���>�  �xi���Г	u+P��GI	T�+M�v�)�N����Ԛ����K�������g���Z#��WR[_��,�<J[@�P��g�)*�4�%dP/+`�#z��:�3!	��4�u�O��G_����i���D���0���ht��������Ӛؽ���&��U��l�spE�<��f��U,d�a���y��6?�r���>stnu����0�A�O�� �p	"�����E�����O�dҨ'����)��c�͟�u�4�_���&�l������xa.�)��i}�w��j���a��D�L��#D	�+t�Z
�Wp^���� F*;y�n���Ve��K�*�x��vЪf�_0%�h�WS�`�A�r����'�n��fX��*�kZ�dn��q)�w����n?w�.j�q~ޕ;�ػ@��c�|��� �U��n/�㹋#!�u�C�d���W����H3mքLG�n�xz��zɍI���[����e[ :� ���i�2]0���Sއ��)M,)6�%���!�!�;tl#��C5�А��A��:\s��l��������d3�J	��q���EȲ�Oh`�p"j����%�iXA��Ur�;�79f�zǲ�5v�u� ,�y�O���}��hH5�]�n��D~���4YP�5��n>�V�>�e ?�\����@����"\�g��ߚ��ݳ�/�|:��v�w������>"���߃$6���7�g�r�����n����j�}Y�z�[�51�.I�^�Im��?M�����{ܬֻ���cM�����������O�Z|
W߼��<��<����yO#0(�ͩ�j�;a[q��ʌ������@��@���B���=���b�]�,��W�_E�\�۫�����ky��\Nh�մ� �ᥐ)��n�����O:��E���8u�n5��	�_Ҫ=��Fn�d��W��5��*~�R�V\a��k5-��W`_�T?�\�������
�U?��d���d���(���=�k[�v�	`����*����W���R��3���}�ИPc��꼖Ƹ��{h׋������^ɯ��G���+��2�c��9Ϋ�%�eT��lҤ�B!W�jbd(,2���jd\��2�<+���i�"6G4�׌[�
�����acj{�'����I����Gm�Z�^} �EO�Ȕ��o�)8C���6����sw��_��l��1�FB���s��+Z�2���z���+��.N/���V�5�n��k�q_kƯ����?��|�
�����׉\�����ܽ".�ä�;͐�bU��z$2puF��L]J\��T�����K{��1��V��'�Z[d�V8��*\����
.�`�Uq�6���vh.q���H�?��\�^��;�&��⹻�F4��c���&h���`�W%:O9���S@U�\Y�+��g�+���D�.�ҝ�V+�z�\7�?�U�ǯKg\7���Wpw��r|F���9a�)��ۻ��!�轋+��֭<�F�U�Jp.0Ƥ�kL�����t��?��T��e~F���O=�ZE�A� �U�ǯKg\7���Wpw�3(��B1�ed��>1]V�
/�
֦�j����Xp���f3�,�U[
ݬQ~j QQ0)Vk�>�1]j�O��T��y��T�Y�Y��5��!�YK\+�=&q4p�Zyh\���B��^�R�#�ժ����gO������8�������@[�+���eQ��a�ZENc^����A��R�H�t�B��Gx]�AWpGDPw� �f�JC�V͒D�V_4pߵz-h\��W�fi�Kl\VW�i�<VeԇŦ�5z��T�x��hMgW���z�RV|�;;�Y�}!�f�
��3�?7�h�f���eT:�"o&�yl,���t����M屾,�i�(�N�"�"��J�O𣾄�3�#��
�0f �ݵ�+��2�O4�[����K��u�m�#��*��먯RN�kN��Y�
/��ib�h��L��Z���U��������?��߮���ٛ�����տ|����9{�����;��)�C���v�_����?��������PK   ��X �x  ��  /   images/0edaf19c-8cfa-4246-aa67-58db36a161f7.png�{y<����3��ڂ"Kڕ%%e/[�P����ن�eʉ�H����K�Xg�l��C��;Ì��=�9����>9�^�?z�纯��~_�}��˺<ۄ� �s�� � ![���[ҫ�?[�.X� ����?Ȯg�� @��u�$ q����.Ӯ����~�~-��RF猴vAX#��i}��y��sl��wwR��/�o�};����H� �;F9�duyZ�/C	l��u��`2�;�r�������?�:��W޻
�Mwu,Mv��.�Z̲��2yQ�M��$����(1;�uw�!����ٮ�a��k3$�j����y����������W�����*~"�-����7���-�|�c�_�#)w�]y�Vc�U߄�<شck����w�cgK�T,��_����/c6�\�.����݋<�G���׷/�aR`;��L>&�c'H'Ä7�zOzY'���B�JcP�j��U��=��l+~���X�~י#A�݋�� �i>�'jcM�W��f�$�2S�<mg�?��[��x|������:.j�2&����om�q5���=:�s-��t	%m��|u�Y���}�V��Ձm����#L2--r3,-B��ݻT���c(GqNEH���H�ރ���w�3?�c�ؗ}�ؓn�};��b�]��"�b�!�®�I���p�<$\u[�`��'E뵲�΅�㑖<H�%ƷQ]6(��[�@��S��9D	U�W	Q	�~�*���ip�J&���qI�CZ?�0;YM즒c�ϑ�,풓��~�H�2s�;�6����o���,�癦J���MF��-��Z׍�k�V`*H�qt/zn2��go�9	�fXQ���mBfz�d2�q��bt�#�h�l�d^x'�f_u�#a�V+@]�\ ��˒�e-d�)5�l����*q�Y7�
��7����^�[\q�1���*l�u����]��H��v�q��GθI|w6�k�3%Kaˊ��!F�K=��K� �}4��%/���f�-c�M�o�9yxU�9Q���y��۹������:h<�����;��}q��n��[��ݓ�j=UT^�=2��z;��& �o�J����ݢ`jcUdK��?G��>خ��-i�h!i|�`�Z��h�+�bg�[㟏S���~_��<�� R���<���ˌ���0���.X��4Y`
z߂M��UrI公�	�y6�3�S?W5�1�N��{���p���S�,�+T�dS��y��;{e*͟���޷	"}m�HH^ЮR/�f�)G���~���g7��+U0P6wN��Ҧ�������wJDZ����)�/^&U��1{�.�6HY ��(ЖDk�����hA0϶��l�V��\��(���]����3���"�@Y�_���'�ۏ{C�㸚?�^�=VH@y�_L5���r0����@��d��x@�C�GG�>�tI�l�V��U��X�ș�"��i�+b�r�4����-�~Q�A�S�������F�[��
�iI
w�J��hҗb�m�5��%�%�4W�,�(O/m^Z������cl���@��>�ο2�e�����sY�@FWN��F���%�h�	2(���X%��2U�Zo]�����'��+�O��Bۯ,��!��wR-{�	�e�0�N]3��9P��i�0�e�oM���xr�Oh>�g}$ҝ'.�*E����yJ�:,��ۤ����g�����p���F���+.��{%�p��� �����cu�3�"����|�b��c�0�e��7�W�eA�	�:,
ց��9|�z��͘U�d�[e���نD�矊[��m��lv+�ocV����/��妰�˪!������vF9O˗�j1w��;��`L<��&�(pL^���m]]L��0�������abd��bA�R�� �������סeR3�@�GV6�$I*�����V_���4���dk��d3_�V,KvCCe��LA�öA!�rz���~镼#�D�3���5��ܩ��*2o4�r���ɓcr�ð6�v@�5��8�=�8i��k<XQ�߾t"dm%�JF�w�����ʃ��vS�{�MR�J�6Hyt��9����!ҩ:h�i��t��,/ ��-ā��k��5~��W��v�4Q>A��w��d�c�%�])I����4��lm9�^�I0C���
�{p$����_q;���Zd�"�VG�E
/o9����q0+�¾��� �*���CF�, {�f�0+3B�=쁷*OF���Ѥ���_*V����<�ٲ!�gjBxʒ��뷷�X��x�b~/�ʁ�d�(�%-�K	�ɰ���l �Tl���u�^�L��(�0.��AgPb�Ө�9x-�ڀ:*���}UmZ&�Rϩ��Lˆ����c8W�XN.>�M��ײŲ[��֡K����g�������eu�
�1<0b��H��Ԓ] $̌V�m�t��5�ؾM!�$��_�y�x�S~"��� ��.�=]�?� �H����͐�W�I@X���o���x�LTO>�5T
�|�����<����T	�g$X��^���ȴ]N�e�971ɣ���:����a.�3{�A����=��(�ҡ��@r珖ձ&g.	Z���׫�5k�M���f��D�(�_i�� �mU+V� �k+��������[ ^7��T�9�pح�&��p�6k��p�05H�`���ȅT��eT����xci{  �k1��>^�֝ĪT��c��6�N�����1�e�g-\Mlf��c��2|; ��0@�E�e3����y�e�{��&�tl� ˧�+@��؅�7�=��O�s�m����s/ii+�!UM�h]����&=�F7ʒ���B����v`�.� ��R�6a���G��r�N����k��:��K�Oe\o�a�s3�:w�B�1[7A��
�
�H�Ꮽ;O[
�x1���������meI`��s�﹜���=\�����DYlQ��!�E!��	�[�/�4�d+�����'DrP&OT�ven�W���N��~�����_$�Ǣ����^��TY�d(AqP�1������ZP؄[�7����-Oѷ.���񛃒�����q�*Ѽ2��n}��?V�l�Ώ��o>�⮹��E,��,�]/�ia����A򯞐�mft�����y�%lK�&����6H��V�ks��%p;h}�i�����:ƅ�\�����nU�o0H�F&�$��@+���ߩY��<�l���O�eh7տ3���G]_�LF6v��|
���w;Q��,[^3�p'����|�/�-�l��'؀�%�675�X�hӈq`�2;f�V\��c�5�9ub	z��k�@g�`���L�ǀ�¿Y�[d{��ؓG��[�k�������n�Q�
;�7�b�ԅ�ũ�ԥY.�*DC�k|�<���
��%W�>_���ۏ�oOuX���;�}=�*�*��g���&t���~�A{ _��)&�:KX�tpD�[q�ݕ�Vp�f�a��Al��*��{��r�3�T�v�[Ti1vi֪�r'�xuI-��'C���HQ>��� ﲐٯ���/������	m`V��%L�]���{�"����z��ďX y�,�Y��hh1�]:d�t�}�W	��|�� �`��f��{����	�+>���.���C��s6��I�T�}���<I��#�x{F�S����� �u���U���\�������f��l���(�#-�OkĪ3L���F� ���@�ǜؤV<���3%�q�§\R},{��,�2����s=�7d`0���V@��~����Z�/�p�=3
�E5���ŧDK��"�ɧ��\v?��Y�XTM|�dY9�W��i >���0�p����'�j��$�F�U �;������s &���"8륭�Ž�@%��qU0�.��]�d?jF��(��$�Q�[��C��ǩ_$��܀gٜYF%����.��W����˺��e<�ħ�3�Y�@�Jq�e�=����5.+�����{�r �M�!���W}�B�������9_�� *-�T�yH���ҳ x�ˀ�Ͷwc�[�O���  ��X����h>��\��e�(�؄"`=ˇ$���Jq�6@x���?�$�5��yE'hi�4̎Z�r�K��[� ��hu-�׭�w� 
$�O��)t���C����-��^{��<�� ��N���UB���Ruc� ��n�\�mro�3H���YJ���~�a�J:�|p];��kR_X�Nw��M=���,��P}
H�M�9:�K�ݞ�4� .}7���I��*%�_��y ���7��j
Oe[,�2��[��ˠ�l˱R�iL3^ƆA��WŃ�
Z
H��j�at��aF�5�K�!�g�!U���v��r�f�=������lאJ~�P���<?l�п�5�[�w�0�fҳl�Ǳ]���3�u���C��ztl���QE_g��A�d��<�6��=�)���J���5d�����v���S��6����tΉ�Z?�\�0UR�p����ﻞ*s�.�F���l�%�a󺜻ъI��W�0̥�o�:s�P���z�5���o�5���4ay�" G��=�4>��T
��}�:�l:��ƳlȔT�h+�X�K}����,..��톫1먽ىt�	�����B���8H;1�⿲:�M���b���s
{U;h����?[-�G�Keԩ?x���l��
��B�\ב�6�NW�;K��Ƹ����H7���Ye���%��W�`���eI���l��_�v�s��_	�䜶\������Q:U��[#O�0Avv�ͥ�������V�J�� +��hr���� `�t�^M|�� /���ȱ�F&��W���;��1�^o�H�u6��(3�q�����>�g顐Y:���]g�Sw�0Nq>�ߗeptA���!��&��v]&	��5�?��#���	-�(����i�K>KءGQ�I��8�d�%������zr��.��*�H� ��	$�4�AT��N���*��Xaz�Y��uW�������p���F����M�0i���Xg/�ۿ���:��/��|����5�F/��u��r.��jl@���f�Ws��|�/�#��m�v("����p6�+��q�U��l0������G�m�h�[��[�`ށ��9��QS���b_���W����S��`��a���x�ך@A�Y+��E� ��O����k@�}����<|��P6ؠp��&
�*fg�����a���-�9;��:m�<_��'z����w�� �Z�����,�<���(2oA&����mr}�������*�}���tf�e҄���%E���͇�
F��x�n�^Ie��g��~��EmP����w�z'F�~G��(�pi�+��uN NF��RF�/��t�p�ˮ��+�dH��r������u�I�U���c�p����X�T�����������w�_�d�ʋ�%6��+�H(øSح��
X�/�=^M���Q@���&�%N֦�ݲs�%kX+�%`o�tX�e��wTN�Y���MOG�`L\��8`Bp
(��-K��Q�0��ϗK<������ʙ�g�G�!d�*}���>n?3;�nHU3QtR{�8�����K��)��ȮT�7��b�*.�c��go\���x���d�n5c�˕?���;�^Ւ���Fw���R�c"SD�O��Mc=�$p�j���h��w	YfKE!��N��KDl���I˽P�U�/��ߡ��n��[�ދ�G�D$=)@���Xrd���X�̪���Ce��e�� "@�x{���h�H�c�g+�;k� �m��C^��**�v���~'��Ah���{�[�%��č?̭�J0��ȝ�	6��">W��j7�S�7㦾�������GV�Z!�]i��k.)�w�%	!��[#%�*��M��b��T-G��=L$�[�V�e
=�����9�J3[�H7/��_߾:��uz�=�j���}H�|pz�@|/�TBLn~���`j5� KF����*Z��؄�\���
�]�����#VΟZ�(9�s~�~�Ը��*��k�C�A��I���D�8'���)�SG�G�m��Ebn�����cy6	�`�
��j������0|xᒕ�qx��	4d_���6�0��S�/�Px߭���1�7Y�f��n���'J�'#��F1ϸEnٛ�����b�*� �-��x�������	"�"Oql8`%%J���9�j˽U���E�<O
S�|ɋ�E�1�g�*[�>
���8a����G�^�'d�~1[��ҕ���9�x����\��,�p�����R�nQ]86����6Vq6nx�y�gW��my� �a�Ş1!=��גΉ7�66c�3�|X@���^�n�\$���eAg�����W?�A�_Bo'����n0i��6��)E3�œ����Hi��4�;j9��dR*�!�Jk�����a�XP��Uy�h��BO�t_"lܶ��K������Ql�5�6�[�<o;�g�?m]s�+�r	���5��<G�j���a0+J�+d�~���?d4���8���{��V b�`��?�10���Bmܘ���-��Bt��q�{C��>�WYϠu��2�_�.����������k�=,�q;n��R<��A,�^�K���{�dʬdT`Jc�Pu��x����R�*qx8�r�i[x�|0��1�p����(w�S�����e��E���� �8y
̺uo��/����6Z�]�5V��#��ژ����ƒ-%�
�
N�I���-3��j�R��Ջ��2���|ܣ�	��X];��k�GQ���i���Hk#VQY��c��\=]n��e UӍ�&��O�� ���cB�>�κq��
�|�b?@Y�uE�V|��k�wS�⻺o�����yg�[P�j�&�mvɚCUEQ�p�_�����ݚ�^�7�$�-y��:�3	Ixu��Nˤ���V�l�C�(�T��U��&�h�`��k����z
c$ Mg�k]V��[l�S� 
��܊KK�v��W;����׳j~�����x�����q�V����xwB^��ꃦ�@	u[��y�K*.[����!�3�G�F��,u���a����*�W7�
�9�>�1�o
��0X�~^�����b����M���Y���v+X��&jzW�����콑ᇽ�%�����q�@�e��������	�gH�q���O���/�/���[�VRf� ?..�����Y�z��J����n9�m.��j�J����!�GPw�9��I>�FIC�\B�rѦѩȦ3�]�\W�XB �F��ɰN%)���z���5㳈v�37Hd����V��7'l���,������V�F��C�|����^�l@�:���mY�T70X�%9������l���h���ĕ���r&���Mc+��3�I4��
d�4���@K2��D80�����q�I�D��.n_���x�� 9y���iC92a��W���E�K=u�-I�!�g�������,�秐RB/�?E0E��{(mE���<"_����41�w�Fyg����2"�R�~�	ytu��H�,+�ԞYJ�CSS/IE�+2A��<)=�p'.�tx�If�4�t:�Ƅ���n(-��Z��}Ӹ�u�;�S"Yh%&�e�8�#F<Z�A-��>�ap�������'{���=����,�ދ����O�_�'��!�?l��H�?i��^ޥEV��
 �k�n���m�3�Qb��0�dVa��2Ϗ�;��eoi��%~�ظ�\
�[����$�?�<A:�6�3:��Y��B#~߾�S����_�8����=(��z"��x�-��YC�@2�����cڨЄ�[�D�[�%��_�deY����;�s��1F�:�����Ҽ���q�*dT���CF�{"��˾�m��ԧo�g�{|H���3�hx��s��#\[d�4ڧ��_�q%aq_A���ǇIh�O�n�G��9:e�K.�˻�|Iv�A�,gW��aZ����'��sT�kg�1���"��Hk�1��0}�����|�_� ���]��$��3Y�]^����C���;�u��_�{��[�N����AC�"P�q�ʞ�T�r?�1�<���2��c(��M��<ύEfuYڨ��1G��{b/��l��룃����"��q��ǖB��
��p$�86ί�x%+��$L����閄p4S�G�4u����ΞR���wx���
C���c��=I��N'Ɯ�~�߂�,�p!��'��`J�y��;�d�:�T�s�E���p��@l�;���x�GN~�yWFq:|�Xƅ�9!�������WY@�RT�X�C}�+�N\�tZTv�,y���:7c7�8��~���G�(
��w��<=�Eo��}��a�[rʟ� <��>�xX(P�QL^D�5,�X�>��S�������-��*t��q�����d0������,�IV��0�M1_�'.zX>4�����x�\��Vkr�%~�M�y'��,T�J�k�1S�W�yF��,)ڟc��iv�=� ��ӋF����rʹ��95��������5@i�!�5�����v#�W-R�K�K�j����w�����#gH�75�V��m4�3S�S�*u�ٰ6P�,��X�Lz$(�������/W���m�!��N+l�M��o��\�X"��TAA[��t'J��c�ʃ��xz~!Z���gF�~ŉ0��G�_��m[���R����˖~�FV#�iñ}yx��)���D�X.Tq<i�:�'������s6�k����#��ںA�ֺ���67RYSwc���j;�e�k���>���Ƙ ��6�v��g҄���	�}�_��k�&%���E��u�|Iՙ�%�d�ik�)�~)�jV�m����z�'��)!���tƂ����ݕ�~f��sm��X��P4�â_���u���;kN��oL�P� KQF��P=�r�@GpЃ��e�=�b���s(���3ز&��pU��ʇ�~�'ƹ�fkJ����OՎ@4���FaC���V��A|���ѴP��oh����gA.H�6Z�:��FCM�~o����2��)��L3��M@"�o�5����"���K�G����vS�څ�a5Dfo���Rz�2�v�����t@����c_ ���[%i��W_���_h��.Ế�㪉���P���D�4bFDs4�>��C��G��@������U�Ӄ٠�"�0��D|E�::����5���6`��Y7&7�w"��D6K�N���k <ߣ��^`Qv�$/VA�=PY�d�]<�0;)~���>���=�[��h	'ç�%���C�j/H"KX5Eg\x-��h��:
�b�u��/��9��FJ�=iyc�1M=���<�K��`��\N��\@�"�h����!��/r���Ov~&�X)ZP*�{f���SD�}i���n�YBo�Gs��g~��+��GިВJʌV��K�l�3T�b�X���_�x�89�'���.ʛ	U��:D�=NL�2pN��*J(J�W�&���w���PJ���7��
t�;ɕ5\N���1���b�
��o��ؓ�SV�����
${�����1Յ�����[��uJ{��.���'����6"k�e���7���Ewlq�{�<7U��~�6���=Sz�I+�J���(�]�Eܣ#Wק>%����#��\/�|�e�����i������˔j璥�[\��:[nw�[�@�{�6Q���:�cs+��iQ�Z����Z�~/�A�I��:�����짜������]�t���ʢ�m�u�Ӭ��ꛋ~��,b[��fs�E�gC#�Q���bϭ���@G�1��,W���~��OXq�P��Π������9W�F�N�t�1Y.�<� �"-K^��L]5O�������9�����ܓ�y+K�Mx7ug���]k�47217�@f��}�Q���8R��e��Ƿ��)�X��DĨꍬ:k�v�kzL['��.������4�"d�G�zp�:���H0U�LJ89O[`���U���LE�)���)�N�mO����ʬ�Ns|�fK���i��2ɲ/�jg���-�3�@��<�ea�hc]Vo�z���յ�J����1�J+goa�m��2,a�2�u��Eŏɨ�g�k��Q8��XY=�'ƇGq Ԣ���OI)V������)�?w.�J�]�����K}��G��H��>�GUX�Y��X��#�@�	��1�uc�eƛ�(���d"ɪ4d�R7с���i�XU^����p�n�՚��l}~�\]��)�șnk Y֩$��EC��B\���~���-��]�������&j
������K����L?������⥊��|j����Kd���� �����+�� �p
�C���oMC���2a���k��>���>s\�f�F�FU��iI*���gZ�F��[F���Y�8�D���4��`2� ���H������D�Ə�[DU-ab��߃=�g곧+Ҧ+w����b�w�]�$���mӀB���e+rӊ�O��&�)?	�=q��L����pC�?�)�����m�u�&���_�z�Gn�{ɧ-��1^LN~(v��90�	t����Ҹ��u!�[�%��bK�{<���׉�-�v�6xW�/tU����~�ڿP�Ǝ��`�.8Ў�4dE�a�G��ei�B��!O�9LH~R��F�6�K��J�%���Ք!�f�m����y��
;�^w�����ꙋ�S%�X9,an�T6���R�ļEc�]�(���
�V�n.���� ��|�j3��Hk=�\K5IJ�w�X�����	װ�7���Gp �4���re0i��Hk�վ��bC�w4H��(6xM:ᛏ����*Rlo_w�z+s�p�[>���_�;~MV6`"�um5_���������sudr���JV2��A���*]>���R��G'�}d-��JG�e����Վ2��m�i�H��^ڰ00ިlܽ��)%�M�r7m�܎B�D�����(PML���)���I D�zu�&:�		����y`*�+?�y������Hk^^���q��c���a;t2b��#Ď�T�<yOIl �JiMjoZ�x�3CU�z��|�6�a�"Q�.����S�<��=P�N���B���&�p�kP2R%���5�_�+���(����x�YP䌡;���U�]�b�i�?%��䟘9�ʸ��։�ݞ���PP�;C�zrF�P��|����8DS[��zo|C�΄����e����M�e�k���E6��b
���p��(�ϢW~���(j �{B�����s���iB�"h���If��9�S`���
%�vl��sW��"sd5j�a�ۗ6�_�q������s����OR����ʜՏ�:�.��/�9U�b�.� P~�1��Z�@"n��)n��Q8����!��k'�({o�Ӓ�--
��X�)]O��r]�

�C&�#]�`�VR��Lٷ*D����I7V�����MD��Wck�O*�Yo4�s>U\͘;�&jGٻ�z�v��>K�_���\M�7\��,M����𠄕}O�"�u} �b<�P]��N
T��݋�Ǉ�6�^��m�[�lǯ6a	������+/>�Y�t@���������A$�	�{0W�os���WG@�f��Rm��q�\��8�w��O�`2�o���nhiO#��;K�jqĤ�+��V�g��0�͂R���>�,�9ih��Ŝ���T�q�ˇ�1�-�n��J��u<=pl�����>���R��\â�i��7��"Y�S��TN��#5IF*�OY�⊨�2�/2��9�D�eć�8V ��pX� c9@]H�u�� F�
���.  ��X�¹�5�U3C�1�L�|Zd�(��NKh,C�2��0��Mz���>���,d�l��ѲL��m��T_�m)Ð��k��9�+�!������օ�z�ˡx�
�	�����w�
D_����w��E��.�@���7��%z����)�BG�p���&��T�D�ݟ�a��gj[�X9[B��be�Ig'��<��?��i�!`��s"�o55K�=�ɿ���DS�|�\|e�k�kO�w|��qh�-�u�e���П��d�z�"�M9�iN����luLɗ��/�Ӫ�ٺ����B�8׏6?���嵇
�!�ZN�N���]�X�gB�Ö�ӥ��q�=�n��o�e��K��duI�#�9 C��U\)�/��E�Z�f�ςlz}|V
X��x?�Cl�ʑ�����0w�;Ţ����v�MG��䞲�GE
��h��%��������|e�t���s���I��HeO�)ř��2�ÿ_��q\$6h��]"�e�Klc�i6���62���I�HT���P��L"!Qۄ�/�(���2��f^�2s
��;z�J��_�\,���:5�j��«����˕�vn$�xP���=�D���f�	������L�1��K���/eώ1�_)�9�$N8�27�}���OF�.[��Nj�ׁ��n39X�����
�����R�I�l�y��*�0y�>�ctj���BOȴ�ܕ1�7|�e��z�*�fg�{������,j�G`�\�J��q5ZDP',t��o#]y� '-0q����v��BHO���⺠ٗ-#C����x���u�$I� ̣mL̩��{Y��^�#��Hr5�ߌ��޳���W�@Xzr�����}��F�r�|���Q��"}�wh5���Dh�}G���CI�g�<�
 ��4�(M��d�Pr
�Ap��T� �'h��p�{Ѷ�[B�k�~�ٺ3%"� ����������@�г}�F����5�d*]ip�6"%���cfP���&_�w�<���%~0�t�x���� �H?���\�r�L?�'h��y��x�����v`�r÷��(�L��͗�!�p��0�P�g
�%�(��2�Ҍ`���v���@22�,�*�_�����얇xV)`�R9yL~���@�A\�Ѹ�;�a(��0��ڥ�^�j�d\�9sxef�R�036��j"��(�3�x�(�a�K��/���ͳ���B�mN魘{i��
��O(M�$�3Jϣ"z<��i����F�JG<��lNP�f����I)m���	~T6K���5�?��_@n�l5|/# �>XI���� `�P4���������� ��Y��]��O�֦ax&{���A3��")�?=ꪪ�h�-���ъ�=ؼ����ٮ=E��#[p q�X��'�r�u	3 ���p�\d�0��d�La�Ã A�]gG�]�d�K[p��54i�9�)��MH�f��cn����hc���5�'Uf6����ƛ�pj0WR�7X��l6GFYbm�!A���Ag�il�c�:D��7Qh�K���E߂E�7<^Y��s!h��s��wUc�wH��`��p���.zRy8�V�	�kU��֞�fˁۘM�o���X=E����L.+/~��b o��.LB���ݺjd<Y���Ԡ��_��,��Rb�I0{Y��ctk<���TA����7 Z�����v������m���Hu�L���117��5$��>�w�E���\�<���M�D`��Ư]��x�#߶��L|����uR`�9Vu�����]� ����P�J驪/�kI�X���K�'!�|�����L����&��3��U��7�;�6.��$�����GmhŇ�Ts�Y�Q炽z��U�N��������s�Pz���NW�8;�\쌧�̼�4�RWnr�iH�iW�'W�SknZ��G�G�c�n��W��G�e�B�fWыo+��I��s�,S@nD���e���q4ND�hq���V8�!�a_S>_�_%�m|�����"��˸�Y�X�d|&~�-z�T.����"��]�R~��7Q:����-�1*r����m��3�~do&>�4���&6����`��+`��oJ�hΖ�1�>J=���a�j1��m��Nja�H�t��T2U�V���f�c�޸�,���������虚�����q畲���=ꋃ�=h	���PhP�{�{}ma�|�?�I��Ny<3/���k7��nL�'V??��٧܅�Lx�A>W����W��6c�����N��N�dN#`=kB`�:
�=�)l@�֍�.�7�Q���(�β�ι�-RPw)��8��A!�o�n#��̟\�Ԓ?m�ԔB�F�,)�{VIx
�I�VEx��&!����5={��wН7;��m��[���������[���I�4܌���JM�Cy}AF.�Q��7Zhw��YY9�Lm�2��$�ql�%l����*=��M�~����·��:s!��?|T�R���P�NZ9��^����;)܅���M�	�
ݸM8���&��h[q��t�:���:���	K�>���t�'J�������EkL�����o-:�Oy#Ƴ��Co���-s�|����i���P�XK����6ㅺ8��@�����T�O#�kT7*Eش�y�7�/�=�d*�(���z�q�v礤��Μ�jdE4Q��'?*q+9�����"|�'�Z=lN���"CeVT�*<�����������.T�����9��}���Q��}*�f �VG��;M 20�AV�ݎ�a�Y����'Y���m���i�q��֎�l��'��(�����;��6?(��&���� �CdVQ��
<O*w��=�6s���i,mԮS�����Ǔ�w���r�ʮ���t�iz��;l�T8��f�Yζ�2��Ih{>��:�ښc��\)y����O+&�S�Ө�2�"����Xm3�;��e�nF��+��m�#�=7[��%����f�u�?�܆��ށ�4��lE�k��z)y�A7��F�Bζ�fӲe}�D�b^.Ud�is��1��� �p�9��y�s�dKX�?p
���P����8B\""�"�Z�s~O%\g���2���3�`���'?�&�|�J�>�}��kGrx�����'�[=騟�K��x|��ad�d�lg6���f�]^za�!�J�sNrh�a �d,�!V;��vo@�u= �0�u.!q$���u�|�"�f�N�.BO��yS�<���y�V��	mC��1�&�[��J�{L����*�N�I�'����'�[jܣ�}�mZ�����D�8N�(�w�%����W�Z>�j;�>܏9����Y��Cs��#�~}*�`Մ��l�M�p[��[8�[A���]�h�K �*Al~b�{��>�����<��5�#L够�� �f��_M�D�Q���ZX��]ˌ��k�f#�/�����W��x�Ւ-�+����m��2���|t��n�[��ќ���k�g	_o�:��`�w	��\m;���j���𘌫_|&�lR�S"��m��s)t!�$���E�>�*��;"�M���lh��{c�1o�\�'�C��!j��[���x�k �����O�ZP��U^�I�"n�M���Xۢ8p���m��fZq�;LFM�!�?�eF�YZ͍�}�������VN��C^��OD^o��w���%LZF-�4r����O�x�L4��ez�M+��I�¼,p�zYIe� Y�IV��4��=6ؘ����:�DEi��}*��tD������M�}��.�{�	s	�O�3�ӃtP�����~q�%]���(k����Hm���ilZ��]�cW��es���=���Ս>�x}�Nև�!y����I�Ƣ��t��U���\�����g�~��V��ye��(��o@������WB����p�zrQ[�����%����p��y@G,��RVQ��ꡄ���iz�D��:P��x^��m�J;T7���qq�̌���$��,)�j�B]�y��w����ߒ*���G�i��4`�%��ϚlC�:�/6��!s�A⫗j'P_�W8*m۸oJ����/�[5	�]ç^�d�|b�����w�����ś��nc$�1�����XY���Z��N6�'�X���e��\^�	��4K�
��&]�h@N�-`�H3p_��	��4'P�%hQf"߻\�C���w�~�0'EY9���>�r��?�vS=T<���	
D�5�az�^DM�g��CK֨���?���n�.�e�r5�HhDl����Sa+�ՅT)evX���<~K�Y���p�����Ҍ��kf�>���s���,+��!�Rڵ ��ƻ�bl���#���g���yN!;�+�>�lNf�@���(�8�\S��RvбŻ��i?o;3wK�Y�I���cԝ��,��:��� ��%��P�Twbndk��Ӭ��sh��*�ebo1���a	u�'��<���%{_fU�{�7=��N'r�� [�p]ѭ5��H������2�^T����Jl��7��躿�r�P�E�`7r"���3����)J��	�cV��_Óg�H�-��Fe�?�Y�{��¿.Έ0�m�]s����2����Q�ҝ�p���>��A���
�^{�$�	��r+3�5�~����k@��^�]�l(&IӞn]oj�����Ys�v��c�A*�隻H��@/�����ֺq^d�*�~O�Pi�P�&aa��V񩬠�a�}�J�&f ?�<֯�Ɠ2\4;��8��ŕ@(���:����ј�T�J����r�X:�(���Q'19�E�}�����YA���)x�1��v �ruz�����@ �(����G��bJ��ϝ-o�}a%葫�K�>,��/N
��Q�=٠MCɍ��i��9��5d��5�?gi;�����{��d�7�j��������$�R(sJ,�{2hu���l�i��i�-���8b����{�V�����e��`�ݣ��6d�A��T�Q�z�~�P�����rTx��8����S�����Tw�Y~:�Q��bn;����t�R:���(��!�\%Ռ����E�'m�ք##�J�0���_n�Y���3u�cv<��ũ��iEC+�,v��ܢ�_7}z�A�Пg��N�V����D�mwM���=�����=�=�6�����Wؕ�C���WNTb�!k:�d)ɾ��(�T(�P$�3:�J�9B�,ɞ%�:#
��C���3�̼�w���;��N����>���������<����=�?Lz��;T�}h�+���	��������adx>�$�7�_���u�+�Z�p��Ϻ`vXC:��	P��~ں�D���M*=�+�'��k�N��%�)j�2�ٔǽ*���~k�F��%̂\���3��7��t�	���ظ��o�8_YQ}ub�tk�i���+��(V
2����U��m��h�݀��q`x�	ul��RP���<*��R#;8]!�����~�q�%�/�D���{��n�%��k[�do�'�WRC�188} �p@��iS�������ʩ�a!����i�邱IuׅC��bbQ��ħ��`zI�D���f�T��K'm��Hz��T�|�?����=>C��ah�Pv�e��"���:��%�a�B�ьl�"O��=�^��V,Y������ J�&g�F/���E ���g�B�i1�iM�a0O �=�Ton �(��!Ȕc��]F����3�u��˲u���T� ��C�l��NPY'��,
�=<Ӫ��.Q���貴��;K��q�C�H�����p��E�f�Q?��}��+���A����a�F�D�5�yB��0�М�eaa[�\����S���{K��P�P��0��5����s<�����7}6���1�X��{90@�������?.�=�$~9�o*��_�JyΡ�J���p��@����K
���fg��º�"�楍G��8s��!���$�{k��PX��H���σ�#�7����Z��GG'��]�T�������@ppp����-c�؜Wߧ�Q���^���67��!o��ӛ���2�p�D��PV�U�g��yv��H%�iH��h�S��F>��V&��G���\�_ �I�DN�7)4��U*`��}���p�B�}��a��]>?��D+BՊ���a�5���W8Ч�z������N�����̞�Ӊ����d�>l͇.����%��o���a�ҜTf�8�OuZ>�BB.ωw�TkU(U1HhX(�N.���o���.snk��Z���*Qd�%�A�bs���Fɗ�qk��X-�v�l�h1*�؅_1�2�3���x� !�������mi�:��i*�CiQ���n�=��ź�Լ��Y���e쩏��_g{OR�)�6}S �؟W$��S)���j6��y��I��u;R��(�R�|�~,�q��V�Y��X�x*�Tߖ��pCH�@ĺ�T�0/]#�fa.M@c�R�_l/�}F.�����ڛ��#B�p�s1��"��>l��F�NS���Y�.VR�>�И�H*(�u�?-8�
!���$����q��څA��w(��'���W�v�D'�L�`5���L�s���%����=�|�{�-�.���u*|~��p�rp_��BU���G�(GS�)4�i+5��au���ɕ���	�e��z�x�ӌ���`A)�O�۾�66��ɹ��.�,��'�"���Lm��������ĩ~��5U1gk��̅��3��f����K���h�c��ء��|��sB�����<�����=��j8͝;J�C.�G0����ʒ��T��W����w���%�ď��9ddj�F.�&�W���*xF���
�F�0F���y[�����d?�{��gO^�Bx˔U��nEc�y�-"�=^��qh�O'D�ݓ�B1���wα�mjL^��/Mw�l삨 ���Zn�&���UL[T��5�<�ܗI��r���I�L�R�D�G����#mΔWäx�[�N����2�E$��!z�Q��#K�4T�(,�(c��<�������/�\�{D���-�5D��~��X#'Fb����z?�Ç ����;}�,�'=S�:˫i^�B�w����;�Y�b���⾄1/�=]�
�L�R�����!��U����vc��;]N���n���G�8-Ԉ���n_I�Bd�$]�8\�h��r��b�!_�O��p-ň�6B}L;q�o�rQ���#�Wﰨ�Y�'ď��l/�2j"��?_����%}iһᬓ����M��1Lex�1x_n
YV���gVZ�4�숇������u,'��_�-�"6%�
0s��0����G>�a��������<�&�no��b� ����e���r����k?�W��-|k�3�������_�Q�2��������9�����Nt9���Vk��H��4%���*-��4y��Qv�(�}�9��񤒲�u�t�f��N���ك�]�DE|�����9�����IY9ü��9s���;��pb_�A+Z'��՜��rŐ�gJ��/K
�f�d�u�S1F><�v�W<�b�Z<�g��	�x�ɼuP��q����X����$�3��*��,�;����q�vH+wqh� ~���u�8��U�͹��GjY�W�Õ�.��*�M*�Q�)'g��t�c|D�,�����[�>�5�Eym�'L�4M�s�Y��_ϖU�]�z�j3�>�2���5Z���{-%��f�ԅ�ط[�K?6/����TZ\:x���CZʂ�����\�*`�;o��N��,���H}|K��j3�f�U{��b5r�6Cyo������d����g���9�zU)X���Ûp��Is�֝>�$���P�����/bVF�W膳'�X����lf� wRP6�3���}`Yj]s���3>q��%ݹ�u����&'������U���o{@<滙4Z�>u��s.���;�~��/�Z���-T^�mH��z�K�ܽf��D�~raS���_֙5S�ܸ���҈��K�*�x#&����q�%�Ӽ��` ��E%�����zǭ�J��
�\Y���Q�-�o����E�1�xZ�������b����z���\oE�ϸ��H�@�4�L3�+���k����4M
E�J��3�R�
��RGJ��&	9�}k�Nj�����/����.���]��_��Pa/�p���C�z���-���xAe|����z3-����cf/9��ʓ<��2Oߺ{�]�W�?�Ic�(�?�Dڑ�u"u/��
��L�EA�kʻ^���3ҴG�.�N#n�(��2*�LC"59j�� ���E5�ED_�����Q+�Ք�����Z�e��5��]��+؛Gc�{�PZE�P���?��*���V��M��LV�n|ï�˒�	�kG*ޚ��;�e������Y�D/찞6a��*C�$�l� ����esN�x���T�a�wY5+Vz���HHꓼm���L"K��Ư��"�Oêq��L�T!SU������u�����>L�������Õ6V��� \��8�T�#;����c�Q��B��N�=�oV}`����
��L'@�<�N������B�7VfcJW�:���v����;v4��t@��Z@mk+��Ց�I��)%
0�8���P��.�m�z|*Td^��gX��<�$�Ø��W�'1���CS����*�4����_K�9��)���5�]��Z�>�F�u´�1�W���"��^�N* ڛ��0��c���>U�t��'���6�87�<��~[�iV�K��P#�J���s;�y�ƪt�����BMS�x����bL�df��~uą�w���Ǉ��Nm:3�$?�/���#ͽ��c�297($��!����-����1�d��^�C��¹�ǿh$]�U	��^��,��a�����X�f�iT��څ�ȏq_{���kI�Mr�qH����U�]����m�����o�g��Vq��nd�V���M=e����f:r�
K�n��_A�e���ڢ<T�E#���X�+�[�'�N���/�ʑh .�jHp�~H�K�������MdCŅ���tݼ�Hߦ��v�����s6 F��_��Mwu��Q�R�n~Y�hW���)�<�1�~����xM�f��#/r͔�Pe��6��ia��|-�ie��;;��;����l�Jq��x��r���۠%�ܣ�R��by(���β<�s^�P�[B��Y�;˨|�Йx#y\�����>��=��]����߯�ݼĮ���&����+>s��_=}�P���1�+.�6���'���(l{Z[�y&~��.�d�2��C�Ҕ�ʜ�HoI�2�22��d�#+�Y$����2iu���CJT�^��@6n�XH���EmDJO����]+���rIP�]F; n6Y0���� ���me��!�X9Y����wԫ.�|�әaa�/}ɺ+��׵_O��#�6Ȃ���G_�=���Z#�����T�K�9RY��p��m*��:ќB(ّf�M7�ԗ��A� �Ӝ��5�N�S������#�_7���	�ҡJh5�{5�d��*nd&؛����3F�9׿���������_���?��(I�D�8N�*+��;�v>�Cd��'�g�S�:WbW1���Q��>��C�fx�xB����g�ͽS�A�ӂp5�������������՟j�����;��4�AI��y6?�K#b�޲,G������]��5�\��RQw���8n�t��ߑ���R�1{b|�H��T��研�Of}{���*X�ˁH|_���׭��x�xZ�$��زԕ�eqГ^���|�f�+`v�2:�s͸O�0o?�����H�{I�Y�
^ꄅ,��A.KZ�)�����܌��`���T�k�P~�.���8kú�,�CI:����b�m��S^n���X��& ��j�H*�j >��e��sKX��g�G��i�3����1'��Jt�T��~�|�H�qm�yR�J�Fʖ!r!C|���Z�|S待=6�A̗b�0N֝�Řs���LŮ�;b�b�����)�=m�E��n�}\&Fm��DQs�,W�f}C���w���>ˏ�]k�$N���֫���썓Q��9�w�q%�/��5�d_�=X�[5�5��A����a�pؗC�� ��'������2�!�1��Ｈ�܋ۑD�8�gU4�ٶ���/�s9ܪ��G%���,�k��!�5�a��d*�NE�N~>_��v�]�&���Kt���D��h|�j �K�w�C`�|�ܻg3`;��ն��E�J8k��;���bE�kM�cF�r[>�
��?M5�L�Z��QM��)8��F���R���������G0< !�8D���Kȧ��z�{�Lyod&�t��d1]4�U������a�rP��Y?�$D:����G)U�*gɏ��5q:i�S��÷����ye��\zk�{���Yw� ��A¹4��ҵ�T�=@/!���}#1��U8A�i�樔�F*��*��b�e1C##�P�5򇄒�IQ�g�_�E���~S�p��<Ñ�Րبgл��������x|��$�~�S���Z�! ���SH�5�
�!�h��fl�n��~#͑|�3�<h7�����y�(\D�s��gd�ZJ�M����/�?�t�nw�uڧ/�+�:3HF���V\`ʢ����|���c���[����$��j�$=1�)!:a��Y	���@h�%�sS��aas���=��2����A?G\E�DeRx	���T�"�Ѵ�q����9<H��nQAZ�����?t���v]�c\]�Q���F��99�"��������s��~���!Kө){[g�6s�eh1������`���5w�V���s�#����g�L	~z��4�^f̷�J�'����~ EX3��O�|��M�#��)�����2� ����' �L�I��+z-,YjB��~���7�{ �R�@�{�뫾Jͭ��b��j�(ּ�>��[4��T�b�NKj��-��!�'���l�o��5��=R'�
=�W��+'���Q�i�1CE!�2�����|u>c}���)u�}V�jΓ���@k��gȝ��'��t�Zu	�
1%���D�����Y���$��<����⨢�̌捠�su�ԕ�e��k(��� m5OW��e��o�����
��ZX�KK[ǮD�wSt��H����2�j)���P��(�K�y�<2ەi��!����w�|���\��Ƒ���L����`���P�%Ļ�E`��"���͚������2M~�����R:���Q�X��%r�&[9��a�倆�����t�܆��|� �eZ"Y���}���/i��:��څ �j�U��f̯�:
��S|�$m� ���ܳxR��+���:���H�#���P��PG�Rh8Sր'H��ħ`�y���w=��9�Է���Q�|�D�"��5d��/2ݿY����{�F�\j��;�%�w���>���+�Isנt�.SF�|1^�8B�	�yZ>�k�h�R!j=%JF��,���Ǎ��=$�����F���~��K�a<O�&�����<Y~�x�H8�l`�\�&|�ވ	-h��`�^��W5�1ެ��AIt�=8�!��?��ϓ
��y�Z��r+7�l$q'����P�uJ�[��C��T��,���#\��� c����|�oB��򋨠�7V���qu�/F&h���`�p�贫a>�d�r�h�=61�3O)D>b����j����%�?'��.c~>EǦ3#�l��R��O�ϑ|�[%���D)�O�n��
�U���x9��f��]�1���ߞ�9�wR���g�w(�m�;D8��y�`�����g�7�h>8��1C�
w�} �Bi��a ���O�x�`������Xd�V��P��s��s���,�Wx���2Uwo��v�M���(���u붫�S�P�.PLJ���n��V��ﲰ��e�����@����:J��-�a�i.�v���������O�����jԓ2G�[宀��� ��<�F~d%�(X�t��8���3R(W�׿�{Q��k�m��+`2��f<�$Z+���$�X�?������~���mC������Q]��1�ř�5����+|�/�G��G�f��s�x�z�ųz�����R����ؼ�aK�����kP�����6����D��Ӊ,��@	����S��ų�kճ�;���HO����E��W��xt�$�2zG���:�,:�gf�eȸ���
�����v~�a4��NS�]��K_�؁�E�o��������g��i]�痢cN��kW�\<{�E����|hѥ&�B#�Zf,��>������+�>�����S�ײ�{m#�`IP,��v��f3���03�.��$5T�Нnfº�L�V��sc7/��j�O��� �N�H(��$�|��΁_gm�(�u�\F�!����Ԏ_㰳(��AH�8�8�2�5]�����9�d�ܛ���ۺ��'GD.:{Ү���XX���d$�T��I�`-��G-4�%���N�[H]����c[Pk/2�����S����в�h_N����]����-b��t� �a��S-��6���2]Y���q��T/���n��@^�!�B�}\:�-[����vt������1i���oJ@y9$�eR��B]#/�۟��x���X�VU�0���x!�.�`Wѻ�[!�م䋪�A 9H�u'�PU�{�Mc:����ޞE,V�;Q��2�Q�j�^���'���]L�F�A�,i�8t}��x�XXX�Z����0���ԯH��D����CF`5_a�JY߇�vE�#P���!}8U���eɒ^�O�lK	�j{�0�S�:d��ǗYPj��=,�ZZ��=� �z/�Ek��!���c}�A-��zU�3#H�l1���P�����c��a���H�e[��[�!�����vY��9���L�œ�z��ai�s�6�#�9lk_1������Y��n�~��I���YjWg�</�I���/��l��;m�:$	�0���%"@qY�s�"p���Sz�@r����0���ZT'\��5���8j}@d^�1u_��wg�_z�ȇ�V�Ø�z��^a��;$���P[�7��P����(R՟�W�'�s�T������>Ѿݒ��0�rg >�.H[B�^M��V>���*Kg�Gȅ=a[����������&�X���f��r�0h�B?��Uu�fS�K��Ӷƹ����O���<��Q�.e������z K=??�,��h+��"� _�F#��!`EDȌd�r�G����8}X���7 �@��g�8��0�#r�D�F�_���«r�Ȝ,F�Y����:�����t*�Ų.l���ߓx/�ښ߃D�O��T�ۇ���֖�Rń�j0�Tj�Ã/;=�	y�(�Cӥ6�H"axKm���R`��6;�KT��hk�5�]���ɛ,rپ�`��U�H3O9��4܄n^F��f@b�W�^����%��n�.�-�B|���j��?���~���Q���i� H,G��=��X5o�����kW��  (�<��w���y�J�-?�(�$�l	�����ѐ���(��8}&�ԝ��}v�HJq�K~A����l�=(I�	!Dږ��5�#`�i@���|��YVu@��h9���m�����oq�����;���旌���B^�c���u�_�ڦ1?�AIO1�M�؄���ۮ  �E��j����Ճ��^���22�p`��ǻ4_h(���&Y3��"���G�o��\���^����#m�-�޾��/���r
*��������LP�nC��g�����>)���&^+������N�M�$���P���%��`t����4���!M�!ڻ�����r'�0�C	ː�	AU��ƽm�z�/���b�C�q(7�e/~�j�5_+�o�F,a�ۧ�K(k@:�K-/,Q��������g��BJ���,�A�h���?8��s��b���/�ʜ�8��H��'?T��	�Q� �%�w�_5��>�2=dE,U�	Go(μ�%���~�aM��`��у�����]�,�O�CI(�!<�����cے!��g9^�YNs'�U��#e��]ǚ�C�B�N?����p�:=��R�j������|�'��Xv\r���b]��j��
�����}���V�A��`=8���������c�Kˁ6!" ������xV�r�]�}��,�/,��S��#��S�M@~:U��lFBq<�U�|�>q��Q!�z5T�DN0?���i4���L��%PfC\���b�j#
�`�3(5C�
*pE~�6�G��x^�|������(�y{~66��7Z`��Y��,�8�����������V�uvu�h��ч �j���IoL���v��5�Ew��I��XD��3p���s<���Z�����w{�Ċ�?5d��'���i`׈Q.4�}(غ��A��+F|���u�M��:(p�R8Mka��k��}HP���W*ލN��
S	E�E]�3�_u2� �����hw
�\�e{1��m�9#W0 �]_1�X� ?�\=��@Gg��6�)��ZtG���4���ӮD��q2?�DD�j>�;0jp�������Mwj�dr�*�H�9u�MA�8�[yʴ�&�HoZ�g�_wP@�~�>dU����g�!�XC8Ǘ��_�M�~�1�y7�j������edM]>���@Qk$-��C׬o%+N�"D�^��	�g5`�Ն,ˮ�נ!��}����!(�}��F|-��ͺ�α�m�J�w������؞zJKB^�|��Cqm����Q1@��tR��WI4�3Bt$+��
I�������@�x�e�ib+���#_yZ&��9i��I�a���e�+#0pi�ō7 L�>��n�$��d��i�����?$>Cm�	C��1�/��g>�6I����Z�͵'y�b_
����\4��!D��`�& �����9���׏�B��b���H�ۜb���Q[�v�GK���l����˨�
}i��I���*��8`�	Nr�Hفo7�J/������*9����$4 �_"�v�oQOHXL6Tq�>�h�\�����,�.CK��8l|��.���-�[�m߶�S'
3�M�1W��#&���~��ؖ�oz��+?���m�zd���-�?�bQ�0�G��!�����UE~�u�%���F�z]	$?�`�s�eG��׾�t�c�$�S��{ei[-ͱK�0�������U�;Ԯ8�AUfy���D��w��}B�S��F:{�& �H���V��A��j�啣6��N�y0�e���2����T��.<5�x�eM�6m���bۚ��˪~Q�u�Y��$c9PX��B*@�hl��Ǻ��b��~>���9�_�(rw�~�]��ҡU��I�lG7��~#���ZZZI�Ūs��P������]{��ζ�}=�*L�g����̷[|�PTT,���Ȁrk�)��LbS�9�?9Zdc&�Y��BO�,��.<���*}��?3�1/hA�m�qmQ� m5I���:�ԯb;m��Z䫤�cÒ+3�L�U��Pչ}��
Ϝv�݈W7����H� К��K�����=x�v3oq���q�1l����T�����z���H4�3��lH$3�Z�YN}'�R���!P��ыL.+ɗ���v꬛�7]��+$D2�6���� i
K(�(>����f_�<1$r&���2�N��u�>}=�͑��7ٚS�ߠ�	p3[.�P=N�\T�Q����1af�Μ�Mr5z�(i�OE Ʌ!a/��cz;��( ���U_���i��i�*�Z�y$�x��h��t�ꮀ�<�bQ¾K(�BzQ��:駖����fG�.��,t�z�T55��O���p��e�F{:;����`��T���1��94ۣǣ�;����2�g(�Vb|U�m�:���2�蠦g�e�Q��Y;"�*{a���"v��'~�S�4.�ͳ�[E��P��Y����(�\L�­}Z�@!��p��G=`n��XA��=(UN�� �e}+n�	�-��O��˓zd�)�ޕ��U�d}f�1��V�ɴ���3�~5�Ҳ56��o�Z��3 ; }[��h>���sP])��E�W���U��_�JM�P�$}m�-�߲=6 /1^�&X�ѧ�rvX���+��T�T��Ǖ&Y��e��_��A�5�7EĨ�!�=�/��]�$N�9��?x�쳝Z�￨����l� $c�aN����E�sK�����)�= ����V6M�w
]9	�F�B�����]�uL-�U�5nbw�E����o�;���s
3x�,}4�Q�s� �A5��:]���*�ث����HoW`���e�$tu��=)*���y�1���'�%�ŴW�b��\�ۮ��h�,x갛8��"'|p�ƿ��w ֥6ď�N}�I�S�n|M ���g4�,kr8� X����z?����o��L�I֌w_��@aF�u����Jr%�ɅLy������"]�C���nA��'�?~��cv��	�!��il��͑X�.�ҿՓ��-�!����b&�'���{�W2l�^�����5n�U�?��ܾ��� �ȼ_0Ke�5�~k��_������^7h
c'$II���9�o�c�hN+���Vx�%
� �>	�1�aW�
������+<q"�XN��^��p:�pk�C
M�]��"�;�W��7����v�
M޾���z[C�$����x}e�+ ���-ad�'6��VX��ɦ��Z���� ������՜'P�MZ��4�����ę>k��6S��f��IGOTuǾ��̶`�z 1�x�Ca��W���18N���p�� Je�����\�)�]��t��a�8g]��+�Rt4k�eQ��vpH��*F���S'P,����jXK�����?��n���6�=1� a�_������WB�����Dx<U�XFf&��NUfQ�9 ,2�J^l[0������ݎ������RDgM����S&7�f�'I�Q�5?�5�;v�K��x���M�<��'AN�|�������Cꨥ�Tj�9MI�_,G�Wո)x��!Ȧ,�l�iw��'��A��,Y�T���?jS����a��,$֔�j���w�/�6T�m�F�J�%jv�U�+��E�C7��y�G�h��S��OYhV�C�@����&U�V��c�<l7�0���p���������zR�˃��<�Y�E�
��,� -Ɵ�ssO�ߥ������RGo�jgHfQ�GM&�L�(�}���sI��5
;�C
\�a�y<��=K��ߨ�g6Zүa	��ÛB��U,������Y�kr�L��0r�u��sJd����s;��"W�e��B�+��K��'gfg||u�L%�9*��B[F��X��B^��S��=etXs��}=Μ��4�ni�����B���cIq�<��Udb~�Up�J���(o��߶)��n�E��\N��.s/x�yݩkz=��4��TS�B�K��A��P��N��20����7O�.��;�������M\eߖaB���K��=�8���||�4���U�O&���T�N�OzG��&���^��f�e�3
m�dH���ޢ�h����?��ۻ�?���s�A��w��H�՝~���ϑ���	�*	�:Ptqo��Y&�}(r�#��B��z��Ժeg]�I�#"���wn	�.�~Y���x̓�2!9&��C��`a�(�s���n��?���������g���8d;�W��1���Y�8!Ь�]�5���lD���G\�M�X��hm��Ǩ���9(D��V���R��$X����ӄ~n�6>O1&Z�e�,ym�8b/K�CQ�I����߱�����B|W��l����u��2q{+��UG�]V��tь�);=�����?��A�f�YC�Ǡuxrv��g������WK�?�>�á�����a1�~u�Ab���j���|5���.e��&��󔞠�DYߋ�����5��������� ��ڕ��]���� PK   �X�X�R�� $� /   images/179c08ce-6e18-4019-8002-932a24469ad1.png�z�[�a�>XJ(*�"���� A�P:��0�]"�HHwwMb��Cr��l�6`�o�}�?�w]_.v}ೋ�9�<�}��|X�k-eJ

JU��:$$��HHn�ݼA�S����p�榠�w���w���wrgc7�⋴�NO�p��������{w���	�s�YY:�8�ڦ�dHH���|�畱��s7���8Yp+��~b��x#�񋈻�jIPH�i43l�q�Ͳ�SĚ�4"^6^DRd+>�[��:�[�WJ���=I�)�C+Ocy�;?(���(�x��ZBD�$��#�e�0,Y�[曽�t?'��|ߌ�D��Y��2���I�o͕7`�6`�Ü	�����`���C(�͚ɀS�@��2�͸�H���j�~2��g��s������n���������:�#���9rHC4�NM]O�~Kˌ�S8_>��C���d�K%I�:���*E�J�<��:��1�u����o�}w1^��o�gx&d�/7 冞��S[օ��*�$�o�}���J+m��1�b���~�`�Q��&k��#W�;O����s����X�tyt�P�2D�DB�Q�ș�p)�R�!ߙv���ZJtc�.����}��4�e����2w�(*1�l�j�['?Px^�h��WD�8�v��qoJ���D��e�IC�g-��'���VثJEVX	8�����d�Mj�e��=/;��R_bK)��u�x��Q\�[W_����u��PόH��m�w�!#dT�}�N�hm�]����¨!��`i��� ��}����{h�9�a3�eHud�u�4�K-@mɩ�����]���I/r��Q��V�tb엑��>*�O>_;tT��̯�.������+mD.�H���i�l�|���a�\{���U઩<���Z��JC��
�py9D��h���=��R�h�_d��_�P*2�e;VE��iڠW]�
C��	�QF���7|h���A_�>�s���m��i�P���s%N�/Ūj�m��h۲b�-�Ώ���t$3B��v�q�z��w�H7	�By�y1�i��v�S������ߺ>֟�Җ��Bm��gx�I��$�|~L�{�[R�e�G��J�������^Jo%�J~V~Fi�����������������j�vU�+R�����v�k��/�	�0x�{<�!
M���T;��t����P�6�+J�6�Il����Y��ρ�h��O1��#/�ݦ<~�H}��^��(9���OɄ�|	��j���P0c��t���4J��ω�#';��s�޾�7&N�ط58�IB~@'O�l��<S�4�N��1����Z ����Jr�� B��DlR��a��`�}i�m¶ַ� �g�!C�d��N�&�����u�t�������[B�|ȷ��6��Lb�t�ַ[�ʀ��c		f	��ϻEfL@N���qx�~"��4�j����k�n$#i�XW�^9���!��M��S)?��RP��(����a�Ύ�*����T�4���7:�e��š�[ܶ�4����FP+���d��{�"�$S��L��3�󿲋�s����g�k������	˦Z�||�ܕ�k�M�7�����?�Tj>�}-��������@����?9k�<\C.O-�X��E��Sc�)�8G>{�x�D�\��u;7�14�N����U	b/���a�)'�q��"�[�?�}����謁Ow�7�lr��i�����G��1�������]����{?ƏL�1���	?��]q�Ͷtω�#��p����(h��:*I�f�W ��3���ښě��݈:��
�$��̿}��k�4�g+G<�������y�_��4�Zz]�y�$� ��Y��Fk�>�Q�-7봃5Ph�Mg(��(�@�G��ݩ& �I��S�Ҭ͠�U]kɒ&�X�W�����Ͳ4�֎7��O�lB�|鼒r�m�]T��M��z���jP�dx���35ǚ��郁{�+�C���L
o��ezC��&�0�z��B�"��}�zi�r9���H����s���EΧ���Nu�B{�rV���4C�,\��.��)9!�[���?.��+��?&�B����w���,MC��f�_˞����<�8 2^�З��S-Y4��[����;Vk�Jl�9�l��Tͦ�z��n5܃�����i�(���B�/�����v���[h����C
���m�1�JGӃ�-�= ��Ԣ��&(	d}��� ��_u��&v�_���F�VDox���^*��_�ER�� 1�8�O��y��+G�>��lpq��ҋ,�۶Y�2<?��>`$������s��[4��eC%e��{�0�m�r*WB^�(Zr�CFk��퐶�=}@��j�ӫk�c/���3b0|�>�7��n����z&@@���5��ڒ���*q��;���e�7%2>!�1M���:�O🸈�|ƶ"ĵ��:�Q���ojV�F�!�Q�m�Xߦ��砎��|E���0����8�Fx�<�6�^�cb"���/�ώ�-8��V_�I)?�rܒ�p��W_/V�.�8���9<�����	ƒ1�����]�:9'u����f�YD�Bo+��wwz�uv��x�_܏����_L�&���L�^ -��Z����D�[�ˈW�	��n3��5��@�n����R�9�����|_�=o�9� �~���+�0z3�=��9m�Y�����K�W�HHb���* x�݊�5��N�(�%��l�{-؏��K�A�rb���v@r�M��c�l�i���_�Ħ���O�Gr�'h܄Q<��h?�I�(� y�X��8@d9���~�/��]C6@�,��ko��A�u?��cUA맆�57�@�y� j.g$"�$� ����q�����Ib�+f ��c���C��̽�?� B^�^�2˯���`ׅsMi �2�����XyFԽL�L�s�g��潓7����)!m�
a���s��|���eNo�*(�m�{;�Ϫ%�?Q�ǭx�g�a{����	=�LHg# ��$4\�^�sc�cѺ�*sgti�*0�A^^�3���Pm���������%���?�n)Uگ������Uku/V���B܅x��@}�ԶWQ���%��ZJ��3�fe�@*�&v��%.�r��]��F�SmH�m��,<�}/���F�-�ukgV���6�Baׯ��U����*��j�]��o(�I��$Z)�����jj)�]���W��z'���]&�ɣ����<Ęj]�8�p�K�SSS"�p������4��V����.I�4�oZ'Se����%�7?�"W���.2����X}xSHƹ�Ъ!Q��;��
�L��F��Z���Z\���N?Ӹ\�J�,�)I+˴�*�4��ſoJ(s��?��V��I������<����B��7��p�A�͟ô�������#$m�
F��g"� �����v����>���������#`�E�xk��+͹�U�%����Y���\���ن����~yY66�MR?p�����V����r�t!TOj��ه�ZoC�وB?�Zo ��?m���q��������l<���DB�S�*��2��B�;!a!bS�-[��(v�Ԕv�VH���5he��k�O�-p�"� i��X���풏���/˟�i�eVؿ.�=�x=3#��ŝsK֊�O�Xu�L4oH���E&l��X����b�*�}����"�Ù٪�GzhS�E	�{+S�ƥ*�1�_̾o$J�=�I�ıE�n���jI�r)�g1'\f��ޜ���@(��
��ɤ�*w�>O�)�-B�'��C��L��ŕ�&3ZY���2�=��$�#ގ��|���y<p}_�3J:S�mEE�x~�Yn�����/]\R�s����ЍMa���&x���4�x�	dR�߰y+�կ#to<�1���L��S�j�������
�ﵖZ�iFr:I��G�����Z:��P �["�����{;q�%��A��"������)w��%�h��̎%��k�:13F&e�m��>�tBnn��qiԖ�ƍ�P��g.������UUL ��i??b�g3� �*��qfw��1�ٽ]�����
dx�E�C�O#��D���		��1J�+�a��Նq�L9���rx����bRի3t�Gژt��
�����N����6~�� g 軳sF���.�:ߗ�xN��[�dM����@�>|��;l��Z*��}�V�R86R�ȇ=r,[�J+s1���~]�d9�{��V-��㞠�+V�S�D���'��3Y���>�e�������k���,�T�p&xf�oȬMı���ætAoL)�e`0G(�����c����j���뎽��� �4�����^ws����=�d(+��Mē���+�n��M _ȿ�u"��g'�ʗS���V�l�p�k[r/�iA"���1��Ϭ��o.���Y���(�	�R��4cc� ��iPP��45�o�[�B*A2B#	�t�� �gs0�PAD���:n�j�:2)Ll��q.��/Lk�fR��;3�3�������*�zO����c���.�ߙ�e�n��{2oMH�n���^'�'��8���[�l�z�3��Z��4�-�$?��P�ޢ��Ym�s�-�n/�z3��pi[��k��@W�����������)e7���u�Lr� ����ǣ\H[)�K#�9��%���m��W��
��Ñ�m��Kb9��˸e�bJ��K�qIBJ&�r��VG%��ilf\>Re�mKX)D���oS�W��1���MF^x~}�V�k�h�x�`���E��I�T�Pl����{l��br��կ[\k'��;�h�&�ۓ��\-���ĺ����#3Y�·��kߪd�q&p�ff<���O�͏���3`wtB��lEG�"[Y�/��p[��4�}+.��	����҆���TȰDE���y�� ����O�8yl(C7�e�/��(�l��/�/�Ko��L[h�aK�]8�=��7�^%�o!bx���챲�H z	6���q��O������y�}^܌�[��L��E^ฎl�νļ=��9� ���L]��=�^���J���+�&�����f��hY�%�n=gRP��	'�vc������1��b=@F˓�;��'
�};����$�*f_��y�֍���&�~jvˡ�o���ml�&:��� �.q�g�s`�Y���K�o�掉��s���..?	":^�석{��%�>F�N)��1����	����|O&�Rqd�D}��9�V��3W6�1�;�������F����G�\����Yƍ��l]������P4f3?)��T��z�����ƪ��m������;�Hxy��W�e����<���d���g�z����Ŀ[�"fDj8Q�g�=�X�	�����`�mfh�����^�v �_1�@�Ǆ@s����&���S"�r��� �>ٶ�*nw��i��|��������-c*� F���ý�*f�1���)j�Z��u#��i�l�����I��	���)z�\��ޭ0��b�(�|��w����w}�,��,�Epl��w]u�tj� >"�޲HB*no�_ ��۟!�o_۱�43md�8��#����Xկ�4����;�v�{mcY�a#�M@ek��O��ʴ���b��)�L	I3�N��Ģ�Ed�3���))�:�؊0d)�L�mV���6�m����2��cآ�V����*�'��Ɍ�ꏈ\�#˸t��6"`�s\��D��x~���+g�<h���HԻoj|���J�0@�[�,s�j�Dtíy���B۸�m�pLV��{�[�3���/h>�&�2M��/!�>�|^#4�YqsJ�[T�TX�� tgh_[q���S�EE���N��_�P�Vn�&z��~��Z>�$?o?m�lO8:t�#}���2㏀E��T�@��F�'F�R3�eXJ�@MߟY�W joJ/lr�J>�/h0���>�g��|��#h�r���9�e�Qlrz�Ι�j v@�AN�P���=U�jc(S�}k���NJrϩ� �cG�/|��Ouԩ��I�'�E���DqLD�$�����Ü՟�C�B���=x֒�K�堟	r����s�Z�cɷ�#�aPxy�@�5+'�?h/N4�c2j�"��H��k:F��N�i���J��>_k�p��A�T�]���wW=� .-<P�L�%Wa�	И+��}6��ǂ��g��*�9��?�5β=J|���7�蜋MH4�]f�Ԫth���$*��*%��W�1��A���3~��(���Oެq�=��R�51�)�y>¼LY�q�K�U�$�K���^�*+Y\�e�*	s��|*5�6=� ��^%��6o]��؍���aOsy�boRB�F@�e����B��$��~�����0��+�H>?��8U�yA3���˓� L;�xn���r琟��s�.�3���"��1^̸rriu�A��w��l�	�A+To�c��c�;҃������]9����%_�V�^�|&��p���#l�w��k$�?ܓ�[���!m���X�rj��#0�X��|���Bˢ�ëMF�!ι�s�ܨ¿��]a�.��B�\��{��44�&�����l���|�]0��Jrؑ����$c�rz��D.�MB��

�6T	�����1Y�3_��� ���K�F�ŝ�}N�R��~�jQ^�&&�-8�|����K���N)�omo�>��-��G��X$ob��@�`����n=�}=y)�=�j"���A%���//*F���pC6_�N��yPf��X���'1�}�3S~�w׿��5�����g��T�\�[���_�+6K�|��"�b��U|�B�����?�~�
�/l;�o�|�-h�D�H>��*L/�)\F� i����x���\͈D���xzs^;3s��r�G�)Y����K�+$�/Q�!�p������}q���9-M��Kk�c��sG�i�}_i��v	]/�G̏��L~�(� �h��W��:�Ϛ��\�(�8��r���#�$���4�04�%av�cZ��jq�?�k���ͧ3�9̫i��g�Ԥ�Ot��-�߰��|L�]�!i˗�v��gēe�[I����;�����n�Ph?���w��f�bE+�y��ch�����9�!7Rv#�yW�.����P$}t$q-hN�QFu�,�p��f�U���jnFѵ�ٺ{���o�4�}[{_����%�-6��1�]0P����N�c,�߽Iv���?�_^L��@�:%����'t�w�?~	<;��_�`Ys�
x��ӓ�h�O(-I]��i{OO��K96�;+��sVX���@�Ǣ4��7gc���:�@�'������f�l�Y��w��.nLv�?�s���6A����� 4����</&h}��3�5z�h���i;����V�mQ �S���u�y����Y�;���jE����ư̿�������{��b/�w��[t�̀�xb�?h�)~t��+���N�N�a�g2�l�ڥN9�҈b�(|�MФ����la{�������eIY���Y����T�%�;7Ь>%�~?�3-ϗ�v���2�=�HH։��2g�P��p����F�r�Ys���3�̉�3�����f=��E��z<�V5q�*X{s�L������W��2����5�q��D��r='02|>� �ڈcP����V�	�]�
���T�z��ޭHQA{�'m�4���&+�c>�n��(;Xp������1�v�m�iIH"4�	�9����}R�����a���;�?�'H/u��(�R�ꬲ��d�p�>���3TM�X>4���g��U\ⶳ-dhO3H�N���(sl��<����~ ��k�:Q�E��G)��`O�b��H�XIP�H�f�:���~���Ox>�9�OQ����Y����K����o�_���r��6�� ��K�mZf���xq��:�o4��gd�i��pD~����;i���{�u0N��=Zy�[V,
�"� 2u�R$8�������N|~�Fr��G�0��ar�A���5�|�<#�2D�ͬ�LL������f.���Y)o�{�ڊ���;c���XQ."���LЪ7��߾8U�_��G����]Y�Dc��D8�׵���VY�Z��K�Y�A��X�R_�;�>j�K��VT|_�m���H9��y�J�!�L�\���7k�ݫE��ۢ�b��;?�J�0����\��ۖ"�\���N��{ypd�nx���h��3�yJ5Eg�)��VN����{X�_���3k��<?L��w(e�BD���S�]<�cZE�Jo�:��jC��Z&���x>�Z�����ǣA?r�Ի� /�6�ԁ�,m�������_�̱հ��� M	��� ��G_�M2����+�J������e����ڎKe�k��Y:��@*KT�\g/�7k���6F�;��*+�777׹o��ԩ888؃@� P������TIR�U�d]++����oz�C=��I���_�WL��Y	� R�f�n��~��wTK�������(�yH@%w}�W�/�����SWL���?����~�.`���ݱ�Z���-&,�6�'��5'�)�o���)�Z���ȑ��t4��r�"2X������"۠ʬ4�����`m{gG����0�t�D��ۆ�b���|�@��/�_���{��O���f���)��Q\�M��=h�y�'�*��K��7O��Bt3č�Д'y���JFC�Qj��H4;R��L&�ԭ��H�k��+��Rg���_6JJ�R#�0#�X&�}�r���}��ƵJH8~�AN���CCC��W��;��m�p�q��,�ƺg��o!xg@~w�H�A�c�r]DkE�wZ��³�zE#3��[����~V�#X��4R����۴�oe(�*���������ǡR��s6�R��߁lg���_rs���߾�'ƕ&J>�gv;�[/��Med���������R�L{Z��bNC����6�#��{�^�L\��z�qn����\C��F�߂9MV�"��[�L�ڊIH�dJ��+�GSEl��ٝq��7��'&
��I)o���bt���՝�$M�6��8���&=Y+�>R(bS��ȧ�U���EC9�	f�O(t/�r�|!?�f0z4C�b!���)��啭���ܱ6���D��� �2���-s%�"�b��-%-u�}��fN(B���a�J�͠�L˻dMkj���'[I���jΒ{fy���f����A���|I�×cL�
�W���bf.=�2���L��ܞ0��8�� |�=�Om���u$$��ú�n� =�۰P%��mN��� �������Llvƾ���6_ؔ�����;�cƻ�Y%��Xd���i�1��A��IB��"�d��</��_���cF��>����+�g�i��uN�;SG)��;M�����O�	�w�5ݷj�����|�	�R1+�5����C:��:����HE8�� w^��$�]Mn������H�������<]j#ݕ�yac���,�,?,���
�����h�j��P ��ŝF����*<��7��$`� ��77q�@_�I�k���� ~�f���aQ|�EGfYEnv�y���w���;c��E
p��(�U��!Ov
=[�q\��#t��&祐,_��?�0Q�[�,P�!TAٰO��\P\�L8�E�в�)�ʘi
�^��^���]���i'�dm�f���*t��2&C�~{�m/bT�HP=>f�����U�<�h7�1�P�R.U�5��>�*'ҝ�J����3큁sk���0m�W;��}�����f��_�ո-^~e�X}�1r�v�K��c�|�2�����ϜӁ6K��W~���[ِ�C���5�{�x�T�@gy��V&{:MF�Y��	5@�Fgy����5��\k���o�R�Y�6{ �:�^6w�+$���t 
��N��*8.�p#%�,Y����zB�o=\{��,�g	A\
����R����_�X�tೲ����V�e~#�f8p�.�^j��c�6I(|����͹�w( ��i�w�g7?���Qv�evY�@,��r4�S{3T����c.�JJ��S�L�f�� 0p�4l	]�����$v����lbf���&?q��vN��$C��2cw
�#k
��6x��:�UT�б7Rq���47����S�~e�����״I��0K{n2.�Q��<?5&�!�J{E��dd/�c��Y'nb��k!��~��v���-u�P���Rއ.B���W}b�E�]�8W�8��^1��#��7/�@	-!!���5^k~�!vq��7�SZ �s���"�?F5-A-_�[�^�gZhz��4�M�9f*��"�P��J��g�X�Q�;���ĥ|������*Ͱ�і�M������]�eJ�q�\G��80���ӟ��H-����RSS�%��xf�Yh}��b��N�m�U���0C9���;��U�m���ڸV�5�p5��5��������0N}�A�*;������8�������)fg�+h.�����2|W�(�|Y����<�g�P%;��R�
[�p�����������;^d/Z<�H�,6WD�ͧ�>�~�K�uZFƸȰL~;�>��j=�Vp�@,�fJ�`��c��{�e��׆t` Y��o�6x|���ܳ瘷���:��	O�\�(��W&���ې�>��q�n�,����/�u>yG��y!i$a���٠�j���!K"?0�O���?3����%Of<f�W��y!o�
T5q�K���p�X�= ����|TW$���A�������أ��|���t����Ψ�s�˰��k��uH����V�d�:�����n��0ú���l�4TS�,U�5%�5nB{i�
Gg�R�tR�`	N٧���m+3b��i�a?���ݢe� ���~��_<���ɔE���aͭ�����&�81�IU����8+�
�c�ȵ�H��h��Rn
��=�,��:{����z��?���}Lhl��m�0��-�r(T��<6*Q6o-��c���@#c[��oO��~q�*��������S��Ui
s�?���Vl)c��Ǥy���w��Y}���ċ�����ew�3��e�7����R/{���D=�۬��㬭*BO��y��9NhpKW�:�f��?5�rq x��p�m��Ż��#���E���i0�~���A��q:7�Ct���,�l�&�����d2y�5���WO�k��c����o�zE?���9�O=�(fƼޕ�#9��x��]�/�GÃ>sIE���t��\�<�ǳ��Ke����(������@
��eU7�Q�0�H&�5�)]�o�g���t�[q���@��E����Y������ѻ���1pU��(:樔GO�#���)j^����Osp��/��k�:ں�� 	r�g�l玌���A-��9���k̡(7YG���k��5��6�1�ZT��&�˛��>$��i	�~���7���2��U9HI�<Γ>y��H_+7V;,�~������z07�Q\�߱b뤖c"�lb�o)�Wg���Ò)J��+���0>�3��&>��+����K~ʗM1��ù����n6v�p�Mf,���r�4́��U�Ù~yeR�_[W�S�ŝ'4[B@څ��"}���������/,"7�].�m��,t���X�:X7G�]��^#�76�'�1M��Z�I���TyU�zn�C!���x��9���'N�H���gq����7BZ�R�[~	����"�� UC0'�O�r7���;�,�x�<���c98�/�r����O���fV�r���S��!N)?��`�'<�cX�@K[���/�2I���vB�8@��K(`#�������s��<�(\���'�EjoVE	ک�O3(�YS2\�����?�ҙ�ҳǣ�ۙ�A\
5���syƌ7(���d�,r�ʰ��E�cH@PiJ�;�Z �����Zv�cwVcw�-�#ئ#V�� T�Y�A�E�ak=�>�Оr`��Y��aZ��!��[�i;t�N��"���)� �c�r�oZ/��1�z��wC���Rp�c�^�.���ڦ?Y�%o��Zj������+Q8ʟ�}�`��P�^eE����0�����[@@ ��㉻/���ys��~tq4M3aX��s�"���U-��J�#��Ƭ�E@��^��,�r2�4������Fa2p�~ᡩ���\���qUYYy���-g0]�ۜ�r�s�Y����]�M�K��Н7�i{�sÛ놬f�㨀�-akc�j�Q�c�z�n���J���ٰ���	z֜YĄ��7wn�� (�/�P�������t-�~����u��;��.X�	�$9�E4;��c��n�[>Q>=]�f
W�ݎ�,�'�Γ���8��t�����1������;�9H�Þ��da]�sY�y)I}�6z�?B�%��������]�Wks�����1MW0��1 c8U�䣉�3�l'ƍ`��L�X�b����z�em�+2�n�-&=� =���ɠ�m�-�r��Lm{�4�D����ҏShK���O��M��f��T~�*�9��U�=����y�&��p�4?��/���e���l,������g��ڳ,�6e���VP��d�of>��g���S��o�O�T�KZw��Yx�����az���3�`,e���"���+��|z9��^��k��,� }�{� ���hP�Jύ֚%ͤF:�E�j�q������,��)��3ulz�����������F�/�^�/�p���5R�r�����Q���r����<Sסp�ʦ�)�Ԗ32�D�v���m�, z���π��J\1d��fj���<��ڨF�;�adDXk<Bw~[&vc{�w�ۄ@M���o�qpx���w���ښ����d�4�AV%�L3��I�)a�ih��OX����&�J���p��'��}�-��o��5��>Mop/�\�&��|�mՓ8M4�9�{��*V����<;�A�U�<[7�����S�ǖ��̡'�a�-b�n��M\uL�l��F9+��!���ǫe�UH���Y�aZ�7�T�Nao���.ޘ2OyO�Kw�3�R�5ͅ��.���IO}!U.9�FZ��17%�=�������,�� c������u~�����W�H�
֝��[V�lC���V߲��ɡP�V��q���e�ǝ`�L��S���g�tu;ٶ�9d�t	4��=��G�xܯ)�yم~u���<H3��?����m�0�Ur����@�����#�öK~��֤$rG��,�:y�_������ ֣&o�ң����~m�x&�K|_�*����f���s�X�X�Ywm��]��i<S���O�&��CE*o�X���x�l�/L( ^�&���1�p��8#�S,�l��qo�u�Ot��M]\��4��jeV=m��9�T�����[��~���R�rxV��{�/����y��t�L��u׻�]ކ�#���n������?�����@co}��N�O���[n�,��+<?�5�<S˅����Q�2gۥ�B��}��{ukV�����7��>��v}�Y��B�aM �y��ܮ�8��'\#q��hq6�a�E����%�Jp��C5�P�=����qq3#����TN�����u������=��	��f�]���n��ƨ��&t���.��㌷㞺kU���)�R�n�>�6��F�߫7lm�+�xϣ���7���Z�����[��C<�O��<�7y����(C��'dni���I��3�W��e<X{�M���yx��q�q��1�^N��U�U�<A: ��K�,�v�uJjj�n9�b���0�����5T��q3%r^S��j�1�i�����]zɧD#Wxx�{i�&���_&k���QL|
���i�Au7�nf\:?����7N=�2F��2Ř㜍��v�����,�����m��}ZT�%�+�K����/������w����'(���!��追��tS,A�Ҟ;�.֝�ܹ���5���"6KpSJ��Y6+{��Բ����5C N*ך��x��ڢ�F��1VIS�B|%�rZ�n��!�{;��P��m*���� /t:��26��8�͵�*��'W���=~�u��̧#�=I~�t<~�^�^�\B^{8�5��Ű���8����{���*��ۀ�����[��Rfւ��BY�z����?�}��P�G��g�7	�P�zr&c:2�����Y��V;e������!'a���ϫ�N��tb�,a�5�u����t�x�ݶ� '�-�������C�i�k6�I��4t|�m�*@�����.�r\>Lp5�0=õ�L�:�(�p\�6��A��î{YU����_�x��͔��-�ž
Y�=mp���~^�î�}s�\�cQ�ٳ�������q�J6�R�,X���{�o��&�£�V��#�Cr%㖕5��� m���T�j+d����?%k���?I���C��d66��x2���f�)֘=��L��ϦB@u�>}�"�Q���vC
�����ʚ�n�pB7V�3Z@�y������<h �@ō��ʉ�
���P�X�a .�8`�w�.�XA�����H��ǖ�4!��1��(����Q&�PB����|�`�K�;��gw��נ��-/�G9ٶ^*ޜ��N����#�<h �q��s/��ϟY��^�O�ޗ�4Uf�Ou	�8k�*�LM��,���+����X��0�h��0��ؑ�:��>Z��]���Y����!��U<��j>\��x�?Pm�S0[�M�1g�On7P�5	�w4
��Mb��I;���*���n3�Ά[����mN�N�J�������V���qZ+��}am�] �mi:@�M�Է��ThY�r�L��c���g%Ir�_����b�+X7~�PvJ�k|�#߽!��a�>m3>�<�ۆ���cn�V��O�$O*��=����6G�`�恉c\3���ɚ�S/�G}�ǯ�F
���]�	�����|v����^���\������&h�H�J�ox�U�v�l\�A^e=">�A�mH�$�<�i�5�}�wL[��B5��
�8�^ �K���w�ʤ��:���S�[�:+Bհ}k��= ��U6�i�ъ����Q3TVM}5�%�z��O�K�!�j~Er�{��mp�5q>`	Kwe�g��g���b�����,��OD3�=�Ҵ,u�D'?XLT���@?�zw`�5ͬ-�W�A��a��_J�������]Ǻ���L�~_�I��)����i��ֿ�1��/~��r
�����{ul�m�V���>�I����,5����*�O��&k������`��w��L8��e�����
���ȿ����>}M�h{�?#'اrɇ��W3�����
]��Z��Ms�E�N�c)����S���ק��*����R`��ǇQ���V��N�M�)!�����OVټ+Mm��2��BP�)���@�ؼ�B+�$(��z}��Y�vV�0��."K3����Yߩ��~([�,)pU��,�(\����1���,��ۏD&ݙ����R�C>]9;N-�rU�5�"j��;�1�kv{���O�.����8�U���^��vL�U���tS֭�d���
C�22��]�)��y��
��K�K^��&�>/8�����b��^-4�5T�1ȸ���,��U�6��Ń��㐹<�*t�b�ʡ]�eb�������<�,i��p�W{,'���,F}^0�␿>��e����;"��^/hii]�uy�+ך�m�)lmv�7���:�@c�ѥ����|��Bf'��/�3�%K3����L]���e���k�%��"�v�e�R��5]�'#�cx�z�e��S�|��쎒��O`���g��pw)-K��O=�
��n��� �(E��&���7E���Yϵ$��F�>1-���n�y�y�2��7	FN�WUpa>>�T,N.��Һrf��8I|V�)ا�\Q�F�k��G���3�������x��d�-��l���SΧ��g�Q��O������&���$�f��6�x�/K\+E������xrV%�y�q�D�O1�q˒�bD�t�81�N�+�h��!߉ى�3?6���)ei����;��*V��Ff��n|+�����鲹��51����U�R���= e>C���lA��b�܀�₆�?�OF^��Y+&300�YuG7��^'x�k�NYg�������i�$��y�&�d�`)���y	���_)E�+��H��_:k3N�m��k�ٱp�|�\Ф��ǔ��h�oM��������X� �����iW��%����~�m3ݕ''<���g�W�����:��͟����N8L�5 ��r�*M���>��4� ��t�[��܇��AE�mOM�$�S�,,@y�}���Bl��@��<N�a��%���V��/�w��>,�a�&��hk������2Zۆ����%DZ����chD���a�:��������q��9�?�\g]k���JU�?�y�9&ȥU�Pښ�*-�D ;�Bd�$d��J�v�����g�x�
ߡq�wt�{͘��%�{F�ʵ���Lo�,VE���%�����������C���J�w^e�8n0!�ϵ��i��O�n�V��n���;����y�e�HJYѽ�̀����5S�c��O$���G���[�Y���d����R�խ=�>�f�O�m�/z��4�A��!ϧ{>��͕�?ܜ�{����~l�'����{y;h�L�ˎf5��u4�%p
�69ٻ������Wo/)�
9�:F�>�Yڸ�q�z�L�c������Ҡ������*�o��}N%�O{?T"c�#c�FaW����H�V���}���h�k�-=��(`��a|�o�k�t�_gT�O��,}P vQ�p�+(=�ٸ_Le���gRtV+��*˳�vD]K~������4�-Pa8!����������/��k3���t^�2��3!UӮ��������M��gj}���;�T����v����S��x9�ي��w�OC�#�68P��o��󦐪4�G��X4�I�?/�SVcy�c�����C	��1ڼڎF�i����"�t�)�J��U=꩙����O�HcB�O6����^�=����
WCf��Yony��*
1�xC��Ť��Kү��b�yE�+�o���gM']�)�PN�J����^�����������GF��Hǎǫ�a�~]C=�D(Ҫ��,�a �����K��T�i��ҕ;�0%�p��A/�0��?�u��Ms���9g�����[�
�|rj,!|x
�`�ǍV��6\W'T����V��?&�|���]�!fb�:����0{{�Z4H'�����=,s+�6���'�A���N:�Y��<~4���b�@aQ����H�:�CU�{툃��o�$���g6ob�}���Eڸ�{��g/���"o���
a�Un�'J=ɗ�)�3���A^]ǿPx��p;ֿ]��G�|�9d�9i�j��7�M����;')����� ��)LB$�de7���v���lt���.a\�5��q������$0`�r4�~{ᤃ��l\�[r�2vU6�&i�|,�����ȯ�F�:=�m�?�����x�>��{��4�&� ��jo�s�����"͋�FNwF��l��u�=+�S1qY�+dC�$�f_SB�4��u�E��~����4��/lGǳ�c.�`:�>�q�����r���_g�gQoy��U�sI�;28}�v
���������,�F�/�\���s������);쾖?Kfk�y��ZQ���j�x"��C�/�u'�G�� RB�{4{#�[���Q�ͭ����%�ʩ�8��s��������^"�xk+H�\�v�X���N���X��b��.ƞ7n]%dk�#���k?d<���}��I3��k'��}����s�+�iWKN?�Ok�.i��I��(	��Rӱw?�Vh¢q�4����Djp���C��C�g|�@T$^;�$n��>���kM������ok��fρW+#�gbt~�Ǔ�y����y�Q0�b��	b��#�����Xo�]$�n ޖ���L��RE\X��D�(	i��u������dЙ����t��oe��=:�����}s
s/��V�Ju.˯��u4�����:������$����hiAOߓ~QS�Jx�Y��ͲM��8�k*��I#\244<��;m�=T���q��zc�v<�m�ے�M�r�������NZ��PSq��Nr�����n�>�F�(I�`c��R�)���gaZ4�Y�D��8t���в=0�$er�p��,G'[x����@�ֿ��RH�놕�M9��Lc���=�ݘd" ?��Q��`m��n�U!��|��x=��*�$�瞇ү.I�ʽ[�I���5���5���s�8��s!�V���Ե�J� ;�5��U�*�!K#1;��[s+�\�[݆�p kMN����䎏��~���~��3���H&<�=����B�*-Q��\~��xk�sr�ق����Y�0�ywY)n�9���R�����C�G�:T�9��l��5,��[Ѯ^�^}<7q�k�@j�
�U�]�.�w��4Ɖc:��-(=l<pi�~����b�'A��	�DL;�����װ�QLL���&'E���o7�e�܅b���74��(~�8c^�'����@[�yN(��,=J�/�K� �� �/5��J�7�0ˇ��;, a�����m� 3}�1�։�ܚ�Q-�ޙ
;��ϑ<�ݏ!������K"u�LXZV!  ��(|��縒Х���hC��jW���*6iJq�[�.L�w�d
�1�n���a�r��Ϻ���/�ey� ��2ǜpX��0�.�!�n�y;�|F,\A��)��>���4F�x%%�"��>�&�L=z:�w���JM1�n����m�~�����M����-ⲁ�K+���1�++<"W�	�Φ�qA�O��Lb���ZY1a7�]��@ ��ɤ�4�pɵvrR���M���WCQ���H�hz|���>� ��%n<����+��:y���7ee�^�ZS��Є�Up�,��3֗ QI�I	�1�>t�>A�������>�s��n�5�v��-����@3wQ�p�g�����+�^f�Ѣ�d)v��QC�S��-D�O��I�0ON��-���_*J^V^}5i�N�ɩ�z��s� ��:@`�:�?)o��+�Q��� ��i3^�e+_`�"��6T徯����D/:�7A�������(�{��#� 4�������_mm4��Ʃ�6�,j��D,���W���(�� �"�n��6r�P9���_*�/����f�)s����m(���aM�\�M����E�(�A��֎����L�`���SD	�航����.�h�Ƥ����e%�Fa;N�oP��0�_�&&��\�&��1��8�[�@3�nF�{#j܀G���s|lj����?�(߭:�q��ыF�ef�Ч�@i-�� ��N\ϯ#��}}����EOHT��;��0��b��ܜ�xF��bH��T3&y���՜+�1Q�ΒrT�ؠؼ�B���s���xc0���xYV�+��bO�Z҇��X���P%S�`�P�?�B����mBڞ�T������xX���y�׿t2:�_WFM�l�'w���o�D���H�/��#��qv����N}�OT}Qu�T)�,!2��]�(�I��0g�>�ݳ�g��Oy��xٹFz�B3a��{�:Γ�g�V#"W����w'��"Oo�$�5���Nf��1�Ӿ�T&'��]c��m�Ej���6��p2g��hFA��d�����l	��0W�k,3Q"t�~��Z�+SX� �~�-�#� ��<����r�F��+�\�����|���3K\܊�
�g�RE�X,�2I�$y;��]�zS���朋�.�v�i�G�9�_Ŝbf��y��Y���u���3�CܯE8�����V�TV��-gj����S�fc��T��9~��~��G"4ΥK?�8��@ �y��R�6�]���g�^~^�G��~��9���qTl�{��C�!5�̏�v�*dR,��<�H=�w����{̗�0$>� (�T�;�S�般:���Ws^w��S<��ү`���HF ߟ�>���V����l�]����\��@�â�}#����\��5�Z���5�~���'¯�&��se���J�b�ܬ��,������U���) Si�杘��Q�ms	�/xq�^�&b�;y;uz�]b����zGt���@i��\�^?W��ERt��㩂�7t����מ�鎋k䕴�V���VF�Հ�L��^�I�U� {�1�Je��ˍj��=_:��\`�yN�o�x��W�fSo*�,�����4��T��&lU�M�W��D��x} ^��,v�����~x�u^���M���fU�$�)0�����h�Q��7���jă�z�����0��* 䗗�@�Й5r���*�Q�éW�Lh���4��&S�i��ǫ�)��o�!�;�'�1z��$���=�)v"��V�J�����z�V7_@gk5�+�Ƨ�Ϭ5��71"���\G�_u$'��b��]t��8&8˒�<�Ͳ�KJ{c ����"�Y�_0�D�)�n]A���+�&�+,6�����v���+i�\���8���'~zGAdǥ_�+
��C  ������a�����8�w���@"!�|�Շ/�>�����


h�x����1��@`�����K��n��Ӧ�#�M�3<K�^s����)4k��������<<����~��MA�oO���&މ�'w��۶崂��_�%�#<j��"טr3-J�C��x�"_���(�r��n��]�T��(B�)�K�_1��[����- ]z�+�;S�<����T��x�?@~����6�%�GF}�����X��|+h�yE����.[!P�YNy�!wCh">���9��@��]E�CK��E�m�'=$t� n�ӡ�pr��������x/x�>}�?����H@�J%��ٖb�����I�uDY�������o�T1��dZQQ��}����ζ֍�&�M�����z@��ژ��
c�l�����L�!H�n��R��#殞8O�]��-�l�̘���٧C��Y�1i`h���-h��s�2��UZ}@������U�v�K��Z9��څ-j��6JN�[���o�	����*�-K_��~��Q6NR*��"��o٨!��ڪ|��K�rO_������F��;Yj���y3�?�ƸH��@�2�'N����6�Q:����^�����x�J�f0��C�r�n��l�l	
�������[�Ҋ�X>#�8���F���s	�mN�w�,�!�Ζ�}!e�1����A��&���:�y���L�m�_T����N��|3��g��h2�߻]�9�~����G�z���t��$��(�x:-��&G��L�7����Yj��
g�򞉪���[��]���SU^�Eҗ���Z�ۃ�h��&C5�2͢vk��R��_�K�TB|ַ3P7�D��!��;O<��q}9(��r3@�::mE@���^��6p���$|jc6)ca�h9���E��+�Q�F#��]��v�/��<�Y����A�������c�\��~O���j��P	��Wy�js�vǲ�^�±����wdŷ,t��Q�ם�;�/e�(7��m�6!1d9��\�+���p�d^uǕճK��wH�F��ϕMj�'�D���hhp�ڥƩE/JK�tl�CEj��#]�i2]������v�N�+��N]�6=ӛr戓�V#���pXFrϰ��}P�sg�~�'牎��<�2�»F_)�Ϸy�~'Lن��4U��D�A8��E{���q��<�_�O���lmm'y��_m��^\^�-68ؤhB�LT���A������㮴��̠���!>�����]�� k���Q�-l���ypc�I��;�ni�:����X��Ĺ]K��I��&C'��#���I�<Ж�פ˴����Yn�C#c�����,W�rΊ	w�I��3T�r>���/Ge��kKo�=T�m
���5��b�ju\G㚻`DP���y^�g<�����%6���w'j��0Oq��V���Ĵ�|��g�W�t�$�t.���_�#��0�Q��I ))ys�ґ�����F=Y��K`0�尼�E���v�}qW�fa���b��hC��3�9�÷��m[�Ѕ��VT@yj�d?�!x�nQJE���$����nװv��q��7ݷ�.a_��+l�g�7�>�B�{����y�K��ܿyy=5����6F��aۑ���\�y+�笗.K>�o;K�˪>��R�}l/#`2k��Eo&�݉<D����Jk[kc�'])�u/���q띇����7�%��N�[N3�ֲV���M\n`f��5(���+������𚲼����gN�O�Ua��A����.8P(/W�P�X����	�zq}m]���tD�fݦaL9�5�Ay��i`m;`eT����\������3 p!5!�������Y�S# y���U|��A��:^ a%�dn����}�{�� �/�A2W�
R��L�A?Y�'������No �����'� ���aB��i�;I�<R'��q��]Ҳ�EM�)ݼ���;�&�|��}��z4l�)���p:.���q���`���|�"���b�$�%L����!{��\SS��UU�yy�i�ܻ�Vv����\P�C`o��a�DEP|b��e�����w?䑼	�5��֞`3a��:N`��x�u�H�.cGw󇣂ȣ�n���L5��G��W� ș�b��9�pj�p�#�K⢩`�:��<��$ݵoCo��-�,�8'�9��T�D���G����Y��8oweV��9�W�]���䁜��P���+{1�Rg�n���[�U�V�����R�JH�����J|rrrݰkU�ݝ��R3����:����Ȟb�$K)p�1+'3��bh������0�eK�Euyl�x�%鰬 �����[�>�u��_b�v@?<�1f��dH�.̢RK����b�h���	ͤm��Vg���f��1�h����'h	�J5,����"Oĺ�8ҡ���1xSڃ���F���j��W�
2����L�\�'��Q��������ϕ��y"�#���g���l%�۽��W�ڴF�48~V�^;�Eհ�Q^K�G�4��(*/�+�,����Bgm�J,Z����+/�.v�%u�sM�n/�먺��X?�
:yȩ�;9p��@�	U����\˅u
s��1��CܭO<)�ү�����l���`��I"��J���&�G��zG��{���0�q�R������	s
�t�E,��u2rř��~��'.�^���3eaf=��0*��V��]��{��Q�%�#B,��V,����Z�v�gG�a�x�m>_������i�޴6F�rpw�����]���/�x�xpL�&ùF���Ař���oK���A�2M��[՗Lh���A���3�4$�\H%��1"�k</�L]��HZ+t�����y�[<���@�zYD\���8���� f+Q7o�:�<h��X�n�6f�#�V2R�sנ%?o�9�gּ���b!�
 V۠Ôk�VࢻFz��nY͏��_"O�p��f����< ċ�@��O��E�|�����U��1c�Oa�?'/mh�.`s_�\��Ee,�w�g����z����w|�fB���i���~��ax����R>��2&MQ��ƕ���+�ֻ�Rrrg7H�F���׎�y��E���lA��e�֜��2����Zq�#Da�(39j��[|;�S��l��P�(��w�Ǚ��R?]hՙԼ4r3�Kd�^�+KD�t�������r{�!��8����,���Hnj�ғ��h����� 3��Lŉ�w��H�3��~�`k��K��v߳��[���,{DZ/�$'ȴ��N7��}^�#++�H��E�~��#�K^�3���$�k�ʐ_�!��]�;<��L��W������;�&Х���Q"~&(Á�V%2���P�(�ϼ=�	s��n�>`�}�+����d~�M�䉌�.^�&N�T�a��l/�4U`-z�Êz�i��ZGy?�[���v��B.e�V�k��Gs����B9MpMF�l���	��{΍F+���Z���j���E��5��i����7��v������v�)���#a0�U�D飞�q5�
�K�T���$�`�U%5���}���j;�����i��T���6T��-�p��/A|������ǩ��-���=�jk�j򹏖[�ү:
b8�˓�
p��"�5q��|�^L���ȒLx����5��Cl��͊Q͑W�@CR�o�4#�4��_���
@r��* j��]���I@�o��C S}s�>zP�nYګ51Y<}(�_g��W[���I����'�����m+(C�㳟Nv�>��c�t�?e�7�(����{E`��&$88X���G��������eg�����O���[�w�,�B?1l�i�G���k�Je���h��w�`>	���Q�G�\�c�~#��9A�C���nf�@�0�\� ��g ɬC��J�#�ט,��8�@�Ӷ���q�i.eΫ�YVZ�������l��zɷDkԊY'&}!a�c�MCk�x�ƈf�"�x����-��n�yDp�ގ6�Pe����Qk��l�� �y�&��� bi�´$߶������?�`�7�\/((h�a3?Yi���Uy���)2�$P�}E:��=�eR/X#���N�4yo`}҂�\�{�@�;��@�tݩ�b�6�^�0���)⁇
{���29�&�ߧ:�F#(�Zp�vF�;5�h:*�Z��Cdmדm����W����r�G�85��ſ�G�%g�]�njڕ/q�l��,���E���� 4��1�8�:�ܖ���@
T3�,�qGR��ppp�^�z5؈��fy�y�.ԜY�1��{y�<��גr�d�S��3�X\j��hs�I��I�%`�ώu�0��}"Z`��aǀ�+}�ž:�����CǭtҮ���z����G`9j=�}��4��%!xZ�����Z�e�@v�+�s��G�i��JX₇f�LbEz����U�<ә^ON����7,�X�g��b7n� cD<Qd+ RW�%`[�M��1�kt�[�h���U��\mYƊ�yK��ˊ�bRy`�U��ܨ��%_�Lj�/E�����5Gr��ǈq1_v ��Y'k��Ϣ��K���ٕ�P�ﯭ���k
�R֧_Ϻ�Go�U�HIt�������N4f~�5Ln1��C�d�.C���:�GC�֧��w��#a�Y3�E��oM��(��Tʦ,���Leg�*]j(=�H� �N��^�o2�� JH�}[�ކ�lO�H8!����Lk{�®ɑߖ���U8U2tg�X���Ga�6���L��}�Y@��?N���ד�K�s!�vܰva˽t�9����ZcccWМ�Z�+��RӾE��, �NL|ÞT�����F ��ys֟<�S������K���o���L�- ���d������FKr����;8����{� ���m:��tz��{<!����=�]��L�e?�&�'��ʦ�OuW�ڍ$���:�E�쬰1O���B�����9z��Ծ�����ᝡ�� T��Axt��z;CØb�����_�\����6#�k��Y�������n�9<I����D��	���W;P���7&t�<����u��ta����-����Js��9Mk��GtIF�7$��~���h�B���Ǆz���-�M�e��~L����G�9E���,�b$��oN�~�@�)�ad� ɸ�.���[����T65��87� ��9[?@�TvL�>��nq38������h_,�����yKG����y��q"�a�Z��JW���G-�$�".B<�x���"��(�q�j�㗭��O��<��RL�;�;�.��lR4�ɥL�D6��5ioj��^V7(ћ����D�zO�3=����ui�-�7"L��}���s<ĳ���V��-,�����d���JJ ��}S����%cN���[��#�E��d��xd:��l��L�hs���oZ�a� Sߕ_���_N��_��n�!�Q#�D_���i�8�)��zޢ�r8�p7����4��o"P4����^��Ru�&뿹9R�ٴ�O�r4���-		�f�����k3,����l�!Z���(�)����w�w�?$��ɉ0������Q��b
)��?P)ּU�KJ�Cۗ4�0N�&����>=o��?�`��l�w��d�?�u��s����S�X��E�c�+R�%R/�R�7Z�R:��˫�'�����K�pk���Y��tU��C
i�
{! ���+ާ�ermpK�����E�����
GY9(HU�����2����+��t<�.��sɞ/ԟ�.g�����������9���"Nz�	�S�M��
�[��jA,�b��Ud-KR�V�q�y�̎)�n��`�U$x~�p^�\�=�?	���_ iFD(���2���{���#1}�k�~����m���s2V���c;U:us�P���B'Ɇ�@0���Ds�G7r�$h�8��%x���p�fW�E�R/�Rꜞ���+���i� �c��j*���h�I��a��ᚿ��I(1�3�%^m5��4%w�wt%��/�(�j��X�(x�ۤZ�?iM�/X;8�e�����J�I�I�**�3�ړ�|����S���z���g�l�N�fnO�InPQU�GZ�l�#YX� �4�!u�C@� �� � p����),FĄ��
2�暺���g������j�"}⋳c\2���s�뼻��Q��9ћ�7�7���0�J�Hơ���4�>��q��#n�9�*��+��B��!�'����[\F��q�m� �o}7(�J,[aC�_�ՙh��S���l˦ꪅ�,�	��$��,&g��j����[�:O���^t�.}���M�M��հ8�%b�7/ۯ����^�u,r� ���X�8|r�	�pߑD�7��p�Y�+F-ᅏ'y�ϭ)@���5��xNB�ۮ�R�˂D��E|���}�F�!?�jG n:ռt2���CkV����KM�N���x�,Q�y ,f `��:�v+$����.��uz�^ۀ��b���*�
����E��!}��/���b�觺@�h�͈�7	X�d0��w	A����}vT�IE�UR�"ؓ�	�#)M7�h��>s�Ya<���]�w0wi�fp�.�fׂ��?�ym���o׌��=e���t��'U���Յ��n���2�D��������M�eO�X.'�m��'�H�nqG�t�0�����վ<��I�f;#i6)k����s?�	H������|����WdA��1)n�h�v��X�N1�|������TTqޞЅp$��������T�B?i.q�""�?*�s���!� ���`lM�M�}�7:w2��h�ˤ�&����s����C�;���I�@��c��A�_ʖ6U)��rE�5�l��!ݎGB���P�����R���?l�AS	���M5E
�V�fң9�A�G� ~f������o�il�	��ʬ`�sf�w+ �w�F�F�w~�B���E��4��~(���<�,�_$���Q�#@.s�9�p��TUU�o��M�V��&��D��i�9��hLf�x��r���N�>��K9���_��߿HĹwGA�]=��F��R��?K�{��Wy!%3�����Sf�C*��vwzu0�S��KG��Xh)5O^j]	7%�q��j���C��A�X�H���x�߮u�o3K�z.�=h'�����B��POe �80�S(PE��d\�E����
2U��3s��w[�E����hN"�f?Ju�jn�XTvv&�gސ���P�Zn��S���g���I���=g��;�������eNo�?�6Nx������6g��/��4�K���pU����A��~G�"�9�#��e�1�Q}�����$>���o&��M�>��O��K���n�gw̷'�1��-Z���@�r	˩�:w�g��nt`�hv�^�Q�\2� M�!zfV�\�J)YK��*���FH����_W��c�5y���Ǻ�O�k��o��0����}�|la��4r��NtLG?m	IT2��ܻ̽7s��kt8]�1��P@YlC����h,I�ƻ���z�3��>z)Xo�n&:u�;"9�����������iGN���D��G�J���
C�͜pe��i�a9��D2`��+8�k���e�ECV�W=�TѓXՁ!�����?ֽi[ZZ&y,�?�gKz��9�U�)�3��?���3����b���֭��{�lzr o��À�ȵ��Er��B�*oء<�0���~����b�Ԓsq6鲛�We0����f�"J.�	.έZ�*�[V㠛�8,�t����n�V�ρ���`\��E��>��ֳ�FJ�}ܨ����}R	���݂ՏZ$1&Wx&�D3�G�ٚ�O�}/�u�o~�3�％�,��.D��: �e9�g���&X��s�&��WyϬ��t��4L�q��޿�ߵ"G���v�<W���.u}/�������������oT#{��M�z5P:�n|'	"9����?���8F�8�����tv"�ZM3��\������a������%	u�R�6)-��2�[^X�a�f������A�:s,��S�[��lG����k���Dq;��,xRSyf�Q�����C�n��p���?��H�):��<9� &�I�J�1��@���Y©F�"��H��}��Π��Q���B��]q�Ӑȕ�XJ%�Ӽ�T���ت��=-��EȔxd8>x��|뗦ο�qބ/Lu�pr_w��utG̻��пO�q7m��%k�فxTr~~���}������P���q&־[R�g�>m��ێ���_��-tZ��WԢ�LP�ԗ����h6_�����^j�k'S����s�"��<k/�/l�M��*��l�.0Uj>�0ѳ^���:���
i�AÄ���(�nY��]�'x{P zȻ�|t�ΰ�#�5b-f>DF�e���ʑb�eaq�y+���u{6��W�U�N�S�{x���eJ������ĨKJF-�:���r�N
�I�U;(����Vm����"H�U�̲J�ߍ��U��z��H�*�½����h�.��#Ű�^�����V�|�N۔�/�R_��yEY�h=���P��;nG���N�����E���Kf�_\\_�&����~"f��-#i���=�}||`�Hx�����,xlL��n*��b�}h?i��ť��J9w~N�y~2-x����m=��������K&r�a�m�3\��E����!�fFlt��T$���!�c����l�$s"����T,.2v��T�+,��Bt�l����Uخ�*�yA�S����6h�!݆c6:��N����T�8~qR���s�X /�ֿ^'#�8F1�b�]�B%���sጉ5p��Ǜ-�������W2x����l�	�Bf�&w���M+����r����f�'Ϳ��Y�<���Z�/������y�=\mއ��:3��C-,�k{��0�dy�&ؽ�W�l��M��dXu�?s�|UY+�~�F�pA~CX^d�d��?�i|�q2ƒ�K�ڰ�0��pMScC?{I)�a�ӵ�T� ��m�x��O��gϨ����y4�+-ⒻL]�t�#�f��7�k��w^��Z|
�Z�e�ծ=j�c�a>Ԏ9�錡� n�����:Nen.�4ĞP�%p~�e�Ap��rq�nY���C}�m���;o�Aź��tǙA�Dv.�����D�\�^R������z!�`2�M�tL��q�,���:����䧏?a�Nnd��V�w��
���/ �;��J�z��I���(�鉏&����{�)bB�5�����2�֑�6p�oS�4�H@�y�
�B��L���yOu�����
pjո�![Z��7�\�T�c��h1�ؔ�e:&LYj��dp� c�i��G�6�qMn�-�V��!��;�@LĠ���t��gC �Q���Џ�dl5�����N�E�Y[6�fX��3|��,�W/�[�y�W�����0{�æ�?f��T���������A���� �E�+�r\�j�U)���Лɔ�w�
��S<]�M�جM��t�{
s5_��b�VW �݉,ǳ���*�@ "���\�� ���	��FF5k�q{�p)th���>���&���p%l2V'�Z�9/��>���p���Gڣo��W2��3�2|����us�j�"m<;��⭄��.ڟ�`0Ե�uF��E>O���YK0�M�u��a�-,���c�^^+^	�C��w}z���q���gk�`�X�|��]�K{&|]�F�$%0�S��t�+�����[��rZ^)�������ۥ���'+m7w���1�>�εV_��S���>��z��;�7v_�g�����V�m&Hg)d_�3��wi�==�1����������;[�"��k?)�j���Ύ�ׄ7ՙ(Ů�y��/�RBa1��]��6f���XJɨ���S��h59D�Jʨq䃌*R�VzH ��-��Ր��iJ�tr�s��:˲��r���(D~�>�e�I���Jq�]��l�_�����6_ z{㜃T��K"��{��5�W=�7�nP$T�sB"���U�l�%^��(�2�hTv����c�%7��[�����lEbh�B���XV�K@����[''ޙ
�9��%�����5)�r#�Q!avɗ[�/Õ��;�p�W�&��O>���8�l|%�wk�.��[�V��}8�ɉ��h�?ο�n̝p!��Y�9��8�­�^�F��#�`��ϪDI�����v��P�#��J����G8�_�-A�K����q�@X�D�����f��,��<��H^��gwj5��\&�uC�y�8�Ȟ�yB���\�ׁ�`Y�+���,S�v�{�:�FZYE��e��Ï�\DH�<:����d|��7'�?�����ʂ`]ht��3�̽M�ӝ�Jd{�1i���X������;���^3���q�Iݼ��-VoJ���ʺYڕ�	XG#��0jB��{J�`@/�f�.����4t��M:�R�ŃqT���i�EI���r�ܾ���6`j�D+@º�b9븶�x�4�0�i
p�5�bv���Q#6r�Uh�Bx���O:lp0�m�-XS~Ȟ���ʹ�/�s0g�&��~H�a���Gq�zh3<��X��N��^�̯]���k����H�O#,{�\b�dہ|�S�@������j����~�����W�_�\��9r���v�=����������94�i72��/]���i;����t��r��w��M��R� �E|`�V(���8�x	Ε�f!d��VQ�f����a6�d�)7%�\j[���TH{Z����7}`��k�k��p���]�Y�w�6��������0����=*���o
lC�T���'��"\Kw��O��}�S{+_Q�L���˲>����� 1Wm0���h�I�9]��K�zv�
3��3
�Tx����\�5w]V�:}�Q����[�߹���="j��v��)�8ߖ�W\���X
p>p��h�0�ZG����x]��-)1.++������:��F[[[ ���=��y���Vy׵����O�v?�@R=�Pu�;*���5S��`��B�B�/V��O��QuM��ݰaʎ�۫��Y5Ĉ^(0�hm�<&6Q쟎_�z��G�yb�.�-H]?��wZZd���ű߹��@�=�zu�T��HCҕ!o��80�����4�Ѫy�*dDk)���_�\��f��GՎ R��R�}�kY����`�s�=�3K�(;�;�IEs�x��Ip�l�޲M�����2�̯q�X��'*��22�Hy��*����� '�[P�3F���4�a�.�������G���Vђ 2�6�L�4I_�1�g������w�x����]/G��1�_M�lD����A�!X.S�4i�$���o�lÓ(���~
ϩ�n�!�T��n&�C;�3&��8�q�7c��J'J��f�C���*���'�(�r(��֙h�����l�T��Y��a�,�m�jm�������=�K���-{L���3�r�^�ʀ��+��M1n��>fc�?�F�m�?�v�zHҦ�:G�H��G5��w%�JFOV���&��e{�$:�NbU����w?i��h�������0Zd����q;6� ��IE��բ�SC~4��X����Ug�@�.]�&r���):��@h��|\���r�FQ� ��ۀA:;��
	
o����m&i�G��5��Y;K8��W c6����'
:{�jd*�+�.�H���6'�h�,�p����z�|���R�@�7tc��P6o�qGA���U�A$��!}�J~�
��Z_��ob�Z�C�߮Rc�<Ē9s)AWs���Gr��ީ7��ZO��'���,��þ���̓[�J�sH��z����=7���^���V�k,|,�7xv �����!���D���T�
�?�VI ��m�V{_��yu*PT'���lI�B��>�	��v�/7c�vK�"���P;W�6֠������cY+++[���K�K.�,�f��"�-�Y���1Y��6��P��,N��<X]U�^�&(V�C��O��e�u��Vz��ă6���&f�Ku���_�m1��.�2�CEt[r����T�A�H\�Dڿ9�����?0�+k�cP����_D��� �H�" �!�!"]ҹ"���"-% ��� ��H	,]K�ұ������=�[�qv�3󝙏�sw-mW�=��|jG�O���V���¿��ZN�ۦ�=�=��[�۬��!K���	�������t<A�o���XX�;"wKn 1�7�	]�k�=2%w?�P	z[�6/�-[�A�e�l������'x(�	W�S1�~���~Ǒ��_���	��-Dh#�I=�,P��ڝ���M ���K��#��b�����sB΅)P��5�����E�1 �%���<n!��2�,�q�c9��W	zV$k+=D�ݨ���E���-6��'״�y_-7��ꏐ��fu}qu:����1=`c�U[��8�Rַ���֩�ǒ��s��.���u�-��X��D�}�7�kq{��4�^/& �R:}�
���U8�?�*�dE>�������!WϞ��� uTT��X��nA!�s��);���\=Ǥ*~�T�����;�I~`I�?>�]/_�!@��~?(vzl��`t��0�� ����d�f��er����w�36�-��A�����'�����G��91��D��!a��DX�S�xZ�vu{V�VZ4�n�|�{�1�K�[�7#�#!�
-R��P�j��ɾW%@A�c�J�W�п���@ѻ<�%�%���G�R�O~��o�+�نw���?\�)&]�x���Er�8��TF�)�2j���kk��0	Ǔ@ Ժ 5BJ�[�ѿ�����toUh������u�?y�lQ�b�!��es��q��]bo.p�xA��;f�Qj�Nɥ���i�z�)��R��1,�"d��؉3/�_���#�����!߸q[z�6Um0�m<�Z�2�?f_D[�߈�+���_�d>U�6��	��� Z��Y{¨n����9.	�����o��t�~�C�q���i�W�ITǻ&��8�uDA��e�?�,|�?�4j/��3v]����t�,K���D�ReX��a�����Oнkm�SnsK)y���J�T,$�Fٶ4�ԝ��g��5�܈�'��oؗ��Թ��H�
)�,}��S� 𥆮iD��2)������?anm&`� )�8���4�����ᘜITG�Ɯ�q�O,��B�����"ވ���e��S�[*�R[��GٰN�OgO�F�X�G�iFP�۪�z�c>�V��o��D���&LV����
-n���L���ֱa�lKa�2
{��%�����NMX}q�?��f 1��O��f�hV �ɧu�%�'餹2ǃ5���MıCؽk	=2hX8�G�j7�1��k�(|iF=Z�7ĥ�w�������Ės^E~���!��h��X�� ��q�ښ^�^��� oSv�r8���r�i�F�jKH!�t}�]gt������13䵃��n�񃛋�xz ����p�@ą����k$t�����v6������/�g�j�W�����+ou���@!�GK𛼺2��Q�>[�i�%�)�,jN7x�:���������!�>��໮�Eѕ7X8�T�%�\w�1o�ϸ�=����e|_'J:�j��+M��6?c��#��8�֭g���;�aC5�m]�� y_����C�%����ɞLt�Wz�tB��s�ns�|g�W�;f�2~�jS��o�3�F�3�-p���>����a����ك�T��.�N�) _��w΅��Dޕi�����m�*}?i8/+cY�ZʡX�qt�%�؉�/~����� ��������)r�ga���A̳�y-b�������&r��u�+�`_y���w�h�hp�[咽<L~�w4BK+s$��4�"Y]�ݱ�Գ�����a��/��Xpvљ�:+ٖ��Ðǌ�°�V�[��"�f�"ӛ [�ٲ�����>߲���?þ�X�?u�F�/��i�^���ȠԮ1����T6_$Lu����)�[���x/,w�&��tU�kr�[B�NR��i)�h����zW34^�s�[{�ġ�T�y���k��?� ��e�����jA������z�����o�b�Lt�6��C������j��S��:�g�V!�@�5/Ft��ܝje6/��!Q\�=��a'���h�#6]����"^7ƛ''1n��5�V�0��y��u�r�N,�Hv��mP�H�Rt4�.���&�`9ۛ_�*Û"�پ��c~��0ؑ)��|�2�DD�U���B@D[����E�y�M��R�-	�=��ÄǓ��6�TV��r
xT�7���2h�x������;!�<r_�e�7�CL�|��'��H虈K4V̏�E��wW�]M��eS���n������r��؋�so�f������5�H$�æ�#YMsK�CS���Ck�`J'�y�_荊��o#��T��z`]�lj!��Թf��1�W��9Y��&��l��,�
��$���((��q����y��
"��u��zH�[ޠW,#t��0!�D���c:\�P-��-UԬg�����ej)�o�Ι~�ER���s����oʢ�������%�6kf�ڣC
���1#r񻭈ms�����)[�[Ǫp���CK�n�[@�k����x�h��T�p��S�Vя+�B}\~�ѕq�<�v�3���Hk��������p���<d�d��[�~$�V(-��Ȟ
�l���{��%8?����Σ��W�pd��K��:��\��:�Hom�߯��1Y}�.S�҉�?�?%-;fg�8Hf^wf���Q&4iٮ�s)ϴ���Vyo��r%��Ā�ILǬ�{٫܊@��������W�&��|��Z�R������טQ���+�0�4�����[7;vg7�3>�1�� h���j�m=��1�5�R��h��}Q�&�a� � ��D$�j�w��� ͨt��L��W@�Xؾ|�����1���W�� '9�����tc;ZHX�kz��X~��',M	裳�H| Ј��M\;����lV���N��,E&քw.1��r�ҫi8�Cr�95q4V�����V��Zn�3g�k�iV�FL��q������˽:��>����4*M��o�����E-3���hR鹖��5&�fD�0CG~d��֣��"_��[�&�E�w֒�Y��SN"��|�!��;)���y��D�b蒡U^�	 n�R�5��Pc�@��:^��c�ZQ웣n��Yէ�+��J��+ɓǎ�Z1SK������1���\>���5o�7��?-<�\�'�pmU���᭦*z��ΙE4[�c伩��E�����ak[��O�m�/'��tXǪ蹭zY+�}Pȋ�q$oe#����^Ѩx)w}Ѡ�ӂb�e��H "��i�ɋi��T��KO�Z�'��q����G�5VY6<��K֌�a��ͳ��iՒ�C�^�ȱ��w�c	��9p���S~�~���l,�He�wf#����b��'���+eR�j�S ��L7`;��ųU1��z�*�O��'J�a_D���K�	I`v�0wDG����H������pSw:�!mʦN�#�o"UÎ�EV��;����KOJHטu�^2����0/��t�>k}U6���(,��/T�l����W�Iq��~X�ϗZ>�N:>1�h��1M��g����&.�jA"I�T����(����W��y�.�e�Y�-�Mx9�iDt��%H7+#* .Ir3q4 �� �̲0|}�#��A�L��y�m�MG�Y���Ij���p���>!�F�V��r�[�(;M��]� �	4@�[c��⦧��)l4Ĳ@CR.X���qRׁ
 �4I��RFu#��fL7��|gwML�v6�h\���f���W��&�6�x2ޭT.N��\(���Az���,>"�����K��~���E�����/�T��������l{�I�	�@��//Ɵ�ހ�c֝������X����1������Xä�L](c���Hu�1�0 ��Q���6�����cx/�C;|�k��yv=�)
���iS�]�~����+�墥��9�J�&x��a�h/$*U�I�>�D7�����P}�x�|8�W��a$���<Q�ٌ��[P�?�G���xC�a&�޾�ɛy��� E��5�=}G[�Ւ�"�u�^�=}!y�?Yq{��)�̅�~t��1��4���Jr5�;?�f��a?t��ܐhd�w5�����!���Y0n+OЖ`k���NCմ�3s4$�A|BL/Z?�xYj�;�Ր�W]hc*q*ݳ� ��C(�����m��0ʵ�-w��/������SE)�\/o�2�$�q�S�ֵ���O�����F��^+l�Y��*�6 '���#1[#?����5����U
W�ߜ)K��)#��^_�Dа�kJwO��
ҭ��-z�7V*�����3�
֠�H��#o���L���n�@��l�����Z��A>_s��>��9��!�a9�c�ޯ����A�I �]CG�%�!.�5���	BoB;�R�c�g-瓪���獪�nD�H�Ǒ�� ��X�6��,���*O:���ps嵙����5�~jN���z��;�O#:��B�=�|�g{��P�.��%���{4o��T��za?r��$H��jCs֊�G�=���Ā�'�V>��E8�P�q+8y�:��@�뵞#�X�^�~��1�m��4)���J��q�� ��M����S�^�,�döe#P�8g�dO~�	�F��G۔5��\I|6�e�� �f��hzL��2t�wja�׹ҳ��n��[PL�$@�d�����W����e��ng��|��7w��Ҿ�y+�����h�=��AN4����C�;;;�:֢i�gg��4p<B�M/1>j�Ư*�9�p�6y�Q$��-�\Qʬ�bl������浌��2oIk�CU��$费��6y�^�H��P���=Nm/�cS���<i~�ν����,��2�'��%lm����j��E�ל���m��+�9��'���v�D�<wN��W�M�U2y���O� ��?[��*%��ӭ�����^`���;��x�/3ц
�3�eEy�o�500�ɓy��!�r5��/p��NV���4�z	U�xߚ���w4p&8ۡ/��d�*�v�C������>�l�ݚQ�^��y�N����Tr|;??_�P���?�s]�P������R��l$������kX���>al��_K�W]��`�/����h.7���S�8��\�F��!�}0��2�i>oC��1���Fs��w��u)��*��&)>o�П�׃]x�����?
��v�x���!,�AUq��m�ZQ~��L��g��\'h�b�e�/	k:�G����[�'�ƈK�����)�7�{�w��&6�3�4��M�?A�'#"y��'$lt���
-�fꚌ�.�ӊ��� �S���9�^4� o��[���؁��0��#�ڒ��{�!n�R�$��1�)�)l���!7-�69IqZ��:�VVR/��������)
J+~9G����9[e�4OI��s����l�Ih�tP���RF桎�ϔ\�g���^`����d�Cȃ��bmnޮ��Gn��qk2��D�Rh!�fZU���-|2�o@�q��t/I�Z]�8��
v��ŭ7P�h�����K�2�W��8S*��7��+*��rS�k�̻�5�'S���f1:�"���d�5z�}�ӫN����$�W{��ƼK�J�s̮�o���b�eBmK9�~HR�t<�׸/�NŎ=20��f�FqAD����X����=�<�T�]���/Y������{�q[����&&$����4����LƄ-��$�kD99X�^N�?^���R�OlR%�u���3�J���7��s3+'\J�6�f�n��.$�Ev�Ŀi]3�l+5���Yd�.�򧴷�(˼�C�Q����� ��z�B���8]�Q��0�Q�������6D�I/XC��X�v�_Xg�m�nJ�5Y���+�K��܆FЖ|aE�w֑R�@��*�m�KFx��t�E�:EQn�x�V�=E&�|�B����M��p���o�_���/�Y\��+&�O%21=����bY}�nk#O2���"���<ޯؾ�0?_�4W>��2��0p_�}��0������ā�U,��o����1�r)�a��s	�8���D�c���F�n_��ژ���
�✪i�%Ne��u���K�0Q���ʤ�\_#�'q�u$�c'�֤��&ӥ~&����v��0�*�����n��H9���g�:�g��pv�[e�O^�Ps���޹��OH��k��v'����߼(A����~Z��z�ş���6�����ʳ!�0wn�b	Km�ڑ�k�G������.|Q��qG���׎u�?��\�	�-aa(UF,yP3_��-ď��>3NhI�f�<��|_Q/������Ў�S^�W�ƆX��!9�=������K�C��h
�c�Tʸ�/+
ό���;Q����Ճ�MQ@���ۍac�s�ؐw̘�"σ(�#�d���\�Z��쒺y�?L��kG�_Zd�&�N6�pt��R����W奋.�扷��<�
:,k��(�����\{���N��ެ�|wݰt
�YȯSh�Å�~t�6�aybA�.2��G��<M�.WC\	[��v��dN�K%�#�p8j���yc5�<�÷��e�����!�3��*����ӕYK��Ye�rX�^�懻$��'d\���._���x�f�P|.+4� ��j7�̍ʮ�������n���q�Bv~TA+.f��?&��B��h����������
c�>)(˕�I-l���8&�a��'ς��6�g�J�*x�<�(�������4�~�3�o��^�D��d������<��G��1i����p,�������I֏S����	G���k7���K�����t�wA�v�����ʇ��G��Їųj�&��i���	���v��@OB��3+�[��'��9VG�Oc%�j���A8�8����~�F|?�<���
?��$�(���<�"��:����3�(ݖ�S\�!�T����݈�P&V��^�Mw7�8>��"����io�n�H��k�]�����Sܚ">kf�pdGKv-�'���n��-��]�w�M�21��M=~�HF`�S���!�Iz�!׫�{F������0��0���'[���aG�7�y���ӳ��k˕�K�OŃe<Y����[x���Q�1�kY�f��N�zn��4��=X�0�S�F�)��g������I��uD����hݥ���Y��b��=WI�B��oJ�ZL�:B�1�(l�C�O�3�������JRDw�F�7o�|@��B�2� '���1Zb"򽲿)�A:���9-��ەK��=h������+˒9��P`��o�����8��]?O�p��H��o�����F;GԆ���2Y����ݣLtNoE�Xa�N^SBF�?��G�U#��3��X����߹�b���w饒s��e�˒x�!�yv9z�7Fm5����Њ��Y��4���Z��ȷ�0�_���*2	tU����(�ڹ
[�^IrB	�v�����La���.���O2�j��5Dկ�d7�n�z���(�L@O�O�_Z"�f�㒸���_�QMIS����)�V�͵���o" �����Z	�Q�V�b���[r%Ha�|n��{��;.�U�9׮�i�A���J�4"��/��G���p���vhBXʃEzr->�P�Ah�y�^�)��Ũ�Wu�P���bE�ҕ=����U���X��80qߺ]�W�e�5����-�5�ţ�hDX2]���$�=�o���E���(�>�,|��W�A;��:+;a�V@���8:ʧ�<�Q��A����F{K❗u^!�H� y���������b���q�1ek&�Q܃���:�MmP�(��HpXGB4؛�ζ�����+�XXLO�'�_���
��{��*�\���I�G��$��\Q�K<5�0t�,�:�/@�ar�C�}��q���37","��T�8����x$����T{;���X��3���E���~�6����n4�b;��r�×�6����ζ��"-�3$K=3��$;�`�:��d�L��U��b� 4����!��rl�O@6#k�/��tz��ǌ��^����b��������Mw>�J����&f�CT1�"�u�s ;�8�tPo�.����!�W�a#1Cd�[^nn����SX���'�\^��~��N�T��?O�������T@m�x �53R���<��K!���fkä����{>�Ψaˮ�h�>���J������΅{¬W���tiS����{撶���d#��E��7��V_��E����ް�X�|b���|����f�lj"��U����]]�U�IF^1h`t�F1���ZM�e!�Ipԟ�k��6B硎�!�@��̧:&�crJ��i8��1��L ���^o�]���r>;�^����%��N�2�b��D��*Sf��m2�_I�؏�����N�ŗ`(*�GI��/X���ׅ�7K�*&�w�]:��he��!<����)��\�d�/iLq�~�I�o�>jc���wx��agyZ,�b�x���{A�p(��xu�d``0_**�[��Y�D��������d����.���_���S�+�@��	x�=q0#�"}+mݘx )��J�BQ�H$�����Bk�D�`�����D����VBgA�mv'x�r��3Br~@����~��f*0jw?q��桢�S�:zx�@h�s<����j��&���� '��c:x6(�ABT�4��)��0�,�Uh�~�V������_��em�KJS��\&A�վ������?�V}2Ƭ�7i����6+]��W��*)�D�JϺwa��׵'�}bh��W�����a�sZ�Qgռ}��mo�Z�|��l�s�3�K"?�@"G��!H�d'�/.c�g-��/�)�[f��#d�EE	`�ܻ�x+r��������<d��Q�;1Nq�_�7P6Lx���\�0�|�+�GO��O�W�`d��Y���@#� LS]�,v�����b�t��9�IZ��|��� �v�J��	����b���ox?@�v��:u[?�men4Pa��wٺ�A�~(h�6ۙ�����N���
�`V��r%2���Lf1]��)y?Gx��}�DPn@�=�5�֣���gh�r�dBO�+��@	��=Dnd���GAJ�gK̆B����3�{rm'y�zz��a��/;�vfv5|,���Yy���m�)R\S���Ǘ(�@�>�GѴ�d./�K���/�$S=�؀����a"b�?D�$��+R��A\�7n�ϱ~��^�q��?W
�Jt�Kd�&T�a't\����X�f���Y��s��odH�+��l��@&�r���x�	�:�E&�#�����f[�:$�4Cw�ܚ�����:�[�J:hM��O%��?H<~ם`���VBk�OX,�Q(Zwd��0����|B,��D_�K�u2��._̶l�<9MMB��{oS���'��7�&�H��܎w�>Y�r����L�__�����/�>C�!��a�?>iY}�F�3�>�w�i�o�-��I1�RC ��,gI���� |��(:x��?��	��=be���y����,AY7:�sغ�x�	�H��ژ��w%w���o���r������v��ں�<*�d�/����s[��|�4^g��`+��Q������S���.���l]yW96	�b�Ǖ����!��}���<�^����|����h~��8����}
pbb��&�ևԑ�9K~���j8�-Ol^g����B��Tq��H��uzn���Q��2A�,qF��`2?�	_�bn]N�c
����N�)�JP��2B&��eE�~N_�¸���g�T� ��d]\[l8-jTe��:d��i���PXGX���|��h��|��G=O��xf������[-�I�/	�4��;z9OW�˽��P/�=��t4	K���'ȲH1ݦ�`H�����h7�����_��VO����_fI,I���]��MK�.����Q"+A$�k+���I�~+�>�#�J+�@R��SyL��jj}�nv4@�c;"�\Ph����'�XeO�e�?<t�w��ߙ�K�MW^
M�ѯ|WZ��|FK#�g��kd��;gҵ�+DYik1[<��&�U<�X�J �2�K�3s""!���X��:�g�ځ��PS`�ؖ�硧F>�>h���5���/��_m�<&�Z��q_��6�`���J�䯡�Oh'��or-�'��y�:P��7#�g�$�'��z ;��'���=Y�*����ܴ�yP{��a�Y����vi^�:$k�x�u&�^\ u��U�d�&O�GvEy20�|Ur��Q�?lЗ���o���G�z�-qS�GL͚+(�$?u�f��܌I4vK/�a6󩈔��{���,N��.]m�l�W��b��$/*5�����؁U��K>4y����΋����[�����f�-9��6>���V6�f��_(��J��,�
�zwh7H̾nhz}���QZ��%��2�[��*\ĿQ�n�@"!c��ⓑ!U��ee �>Z��t���I��7)����V��׽S;��صQ��p�v+ʁ[�3���9�{>��y����M���=[+���V�'Jl?
*��M%̆P����H
K���((�~����<����8��d]�i�4�X�Q��\�A���C'�m
{�(�'W|��j�M������pG�	v<��u>KM	�P��',��oɐD����1�A��	��HT�>Mm9���x�����	陋��1����7���Z�j�8��Ua��?�����h\ 7M8»�����ڱ�X�2@0�=|�u�#:}N��#�n6�Po�:\:.��
\�qX$����L�����݁�q!#ugR��q���9���b��G MȀ�D���n���ੑ���t��z���з�K�y$��T��[��dR^��4��	�{G+�5VT�ku��k�T�ReĆ�!��Բ��ʓ?7���OB{���Ax������wt��a�$������ ��*�ܟ(�ٯW�\�C�!W�����`�ۮ㮻�����2q�1���NQW9k*'�&u�����\CŎ��Z щ��-ߪv9+�����a~��˲�uÞ��+�w�+��S��<�/?�b��g�TJ�H�[xK&�o1����)���x'.��I�\��k�kl� ���h�Ê�Q��V�E��ւ�BdH�h?�M�D-2�nqNƗ�C.��i���� ��:1�g?d�l�M&:������3����^�c�|Pa�mH@9��h_�e���=hO�С=��ى������%����1Ĺy�׌=rT�'p�μcWݵ7Fa�SMZ��םD�|���">�=�0������c	�R�-�T��Kn����S�t)�p�;�f@ Z]=p!�v/�a�)�[`B�{�d�0�w�[��[1R�o��'�'�d<R�+��@�~��iOe:S��a���(���*%1�FJ(ߤ���~����	k%Q5�-C40x��cT�Tx/q�pw�X:��fE���z�?�Օۺ�x�S�a��{�=aT���P�L_B�ˆ�E�an��pP��&1�lW3��&�n���������ߘҟ�%׉�_I���}��FN�z.��j�C@�����������A��:�z�㈃cV%�7��e�F^����^	�ZR�*|к�e�g�WÜ�1��Z�Å��+���& "��y�v�X�(^��:ڝ�*�v�����ʣhʮ�nt!Ao�F@�F��O��S�+Y+��ػi�1��_����V0:̒����'Ԭ��$�'M��`<�_Rd�S�ym��mL�iR�Ud�R%/^~�5�<Wܼx��i,m���C�h^�~��9�&Y��?��!�]� ''�'�XK,&�	�=��$`���^�F�t���=ޭ�wl�L�D�]�t�9��osu|�f'�#�Z�}	�i����l��#��ٙ���Ϣ�B�f����m;q*Y���aM9�*���S5�2�_�W�-3�?���.>����B�E�C�,~�|D�md�ڔmhR!���������")����]jM��L��%@��(
ſ�����d���TӋ
�����UO�8�	2ݘ��;�2^�-eY�J�WJ�U���6G˓�T��S�+`�Gx�J�D��SX�ZدF��
(���}Ʊ'x����9hG����a�v]�؟�I{b�cN:�e�KW΍�r��YlP��V����-���R��x�V���g�m��g�˺. �LC����'�1P��4j��Ax���$��������SӉ�ϕ��;ʾ�%m��:	o�)����B��������u�n�CӝrA�������LH�~ʴ��4}yM�p]��Á�"�tS��1��6@�V���ۯF��W9yh�ʯ�Gz�v_a��3+4�zu#f����q�g�o&�;����:�l�Xz��x�����~{n���C�G���A�|�.��ڭ�/5����R��)��$"]"�fŸ?�y��庮l�);~�g��b�.Q�St=_���&�O�B~��SD*ae�E-��z��G��L"�ymC�Z)��a��Jm�Vy��\b�ѯ?�1�M{�{ϑ�E|�HK�{�"���\�����KH�����]u[�jרC c
�.1C�WX,�K��t�gB�}}��Wo�G�i|�
ݓ�X"�F���hvV��A�(�9 �L�#�\]���G���#OQ��W�}��A�{ �/�8h��p����`���Y��j��h�����c�j�m���p��SA��X�����a�q����l�ʲ��?��Ћv�ҙi>ȬJ�|`Gg�����:`=?�+<=`ѓ{���4KV��3�W:���dL�k��,jR��3i�LQ���Ӹۃ�`_&+�D�w���~�ڿbYW/�4���T��´R�e����- �<�o'��Eo�~\6�j~��K�:����YxBᗜ𩬥�;�l�ҕn�ƚg�-O��d�F���T�ŹXt���\�C�L/��^ltAj����
-gE���J�u�v�����[oL�p��8��Z���;eP�:W�͚����}�0������$I����3>���8��4�y�{P<+?�p|"l;½	D���� E�s|D�u�?��W�lU��x�ט=�K 06d�6�$���E	��O�(]$�V��w����D��板%�j��B����طv��z���痣a����\���p�$�{S�a
�^�f '�j�qX�>-4$6%��K���g��
ؿ����.5����
Y�<p�� f��>j��K)��N�����Zu�鮊L:)�}2\e:����"�Hx�
�Oz�1�K��n�	ZP�g� ����f�v̺�?����L.�}��`�&����©�*����i��$����߰Z*�)e���НZ<��r7���h� v=��g���_�˓�����$
��:nҩ��H�NK��C�9?Q�,��f:��c�,�� ��OBQ�5\GVh}�ܳ��e¤���n�f�F��J��
�@CA#�:j�"g.���m��X�p�#Љ�3� ��F5 ������������%�oG�E�^��&�!!���-���I c����7[���~V��&�Uړ*�JQh�T?�8L���}�kJVK�O�n��gM��%�u��$5f���i�a�9���t���l��wG̣����%�f��5�$�(�����g��f��N�~l�E�.����� ~cfy�52V�y��'1v/���_\�~-����Έ'�#)�)YR�����7��o�j���s�q�(�J� ����$-k>�8��Fak��mR�?p:{A$�A
t/"��a�5U��s�;-ʡ]��S�A��H��zy:w�ې7���&�a~���V}1�|W��Owl%����؟Mvb���b�3�X���A��\���ǔ^��%�<����(?�!�k�r���4��v�뀰b�Qm��ok3}ۺ�s��D4�^?��
\�u�D�^�a��Ѡ��'Q�G>ܤQ$,s���5�����=�=�1��}=o�%3N��oCy�M--쬀B
�G}��0�%�\ω�Yom�ٽ��m#��8�����������%v�ի0���iQ>Rg��J��vQ�X�����+J��UȖ��Z�oUf ɥ�$2�o-�U7�6�4� GZ�q��ʐ�[y�"It���I����
�Z�ͼ�<~�R�=�B���*��y�ɝݷ�w��K��3��,�`5�����0����(�u��J��Zjp�k�!���<W��_���1#Q=����t���˛�'y�l�n�a���7��b�͊f��̈́ٗ���]�/;�����%� ���$�N��V�'y�R<"�������f�'.���8�����ê�FW0Q-�Q�6���G|R�F��u�z�7���!�1�M)���F%}�z�W<bS��W~�G��y{�K
��)��#}�j�s�|�j�""����S*]=y���\%��f�!��B�сiVO�j�>[(� �4?��t�j�����A��� nPR,��HF����~I�O��uF���2��^-��l���^�s�ŧ6��	 �7��o+5�s�x����<7d�D,̶�^ׇ�� �ϔn�JnlN��e�7��a��^V-�M� c��r0�L�p�i��:[�$�Ч5��""x�0�Nc���m喫��*A�Z���'���������~�� �P����)�;䓄��{�R��i=���n�k�7C��`@'����8��X���;z�̻Tn2ei�Si�+�4�y�o"����+ڇ?d�|�b�v~�$��-��Fݯ �����N�;��h���,=	%�G���s��1�{�M��s}��ΧZAV��m��;x���l$a�D	w�h�B���50��o�Bo���ҙZ��� [��~�y��h������S)�<�^��9�C�SE#��OP��(�}���b�q\��a������j�{�]�=SI��ajM�W�}M�@�uƾ������_�5��t���p��(���ϩ=I�����o�fo����\��Xչ�<!ݐ�&8M�v䨐K�d[�!�Q��W.��O��OT�w��wv �St�V<@�Ӓw�n�E�x�S�� �P0#�9�q�GX�Y��B焷c�4T�����6��)ah�j�l{�}�ջy�Qo�T�k�'�h&�A��bI�f�;G~m��4l���et_��� i������2��,��������p�9I:Ŵ�O�f�����4%�I,�9��6�Z0Mu��"Lu�w�.'�Oi�a���W��XT�2t��,�*A.߂ǐ&���	a�B�/�݋���*p����.#�6��ʛ]$_������tm��+�K����ª���t&K�-ʃyr_}�nDB���_�G��s�+<e�	k/�5��֣a�������k[f�j@��
��:Qƌj���{�ݹ��H2�����~JD�b@S�c���~�uwԤ!׿vVv��ڎ�М�@�	}k,�����3+���Jj�1�9��&|@������A����W��.q��3�<)"� ���"vHo�t�LSA]Z�HS�zF�2�'�a=�՟Ĝ�҃�)�چÏHw5C3�ܝ����q�xA�=xm(�D_E�pmw�TЅ�極`ˑ���H�[��ϙ�Dvs��&t�C�w�&��-y-b�o+l���+�Y��҈^rT#�ĺ������w����<=))��M���IS��PA?��Un�����S���z��o��*���mlC��|,��_Ȥ�]p��C����Ȅ��bi=</�1�c���]w,уS������O�ʻ{�s��'kUu�|�;>�;�Lo� ����_I5�U
R��v����7��n��W��K�`^���%2Ϳtf��7��@���<ۃ�%&�%U;օ]sMc^�I�}�+��kc{�\h�9	M*T����x�J�N�E_�c�?�]�3�S#hr�0!܍A�/E��KtT�����D�������P��{X����5��@�b/Qs-�Y�g���`�m|��g+�*�Fa�l,��\r���;埊�8*��5��9S�*!���L1�~�D�x�['��n3uV2�l�K�lf;�D��N��;�W�u��X��[t�~T�y������D�e��E�x��W�a�X��ݒQ2�՜'-A�w�
T��c�{��#vم����'�Ť8�1��*o.OA3��<2�`���C��]�t"�=����4�"�Et�+�=��T<ŦA ��>a��"BF8V��pfq���P��`�c�#������Xa�C�RF�*M�p}�D�P:U��+��p����)���v� ����6�w��d�-ſ����j,ތ��[�7W&��fKx��𮞛�FH\\ԝ	d,Z��P\��k�jSA)�L:�vB�F�݅d�
o+�U�W�������[xE�}a�H* ��#"�%=�4�%�HJ7��ݎ���20t��w@�����޵�>��������]tZQIؐ@4��{W� 6�J�9��}�_L�����%�� ����:*��������A���=8'�F~�����R���O��r���Ɖ��8U���^'T ����~"��4��{s
|�'/9 >�<;oV�bFio��Q�<�G�?绩
ֈ����KtʥI�#aC�)����w��|י�u�>�f�n��<�0�����4�1�CF�c�O~�'�o64���#y'���F�2��M�/6��`[�78Z���˭X��{�_�-5qgz��83F?F{ >:e��&�Hϔٷ�.�&�uD�W8�������<�.[���s�#�scG��K��2�����^c�8cu�	6�Z2�&
��
��`*��� �Qf0� ��a�[>^�)e�N�v���YZ=�:w����H![�dU�NtH�$h��g��+���l�s3��+�'�����:�l��N�����7(��J���O�(Z@W�)!�lb`V��Ʋ����� j&�jD�����\��7�2k�͑�ݗ"9��Aρ�[�ߪ������07���\��T�lN���^~�����'�Z^���Sx�0�ۃ��NL|�':�f��t ]j^���ʸ	��W��d�;T?\�ud�L��_0���R*����ΉG$'F�";H��p���9
N���M���(�ʖ���}�N�Qђ$Y����U@O[z�z��]!��a@��Bĳ|<w�!�y�|=i�[|C��⣭��:	s��X؉��WC��<jY�A�6"�4�uMw��$�d��Oqyi��
�Z�(��0�Źݺ.��]�T�e: R���}_ �2�J�6��r�cD4�o��(�t~$x��	y�F2%i���Y,Z�V���K����f�|��9�	d�L������9A�<��(�� �ψ��S�i��.���VL>l5i���]���
ȋV����Y����U�3ޠ�|!�9��f:u`���i��wh�釐�?���H��AZqq���Fl�	&��8VR3AQ����{3�¼�v���S���~yjYGa�q�Q�m�saۈu�8�ĉ[��z2�nT��:^���q ���*?��^�)�PÕ��ViKm��؟yү�k�~s�v�r�#�\b-P�|�$���� � 
"��I�����a^�
9�nx�p���~�O�M�[F٣���7A��AҽZǉw�\̃������"�Hb��A��faԊ@�\dӾe/F�q?1�pF�㥞�\����5�K���=Y����!�x1�E�Rn���
�pHekzy���C3l���8�5OQh.��X� g�+�C"�W|n۔7��+�y���|�8�9&�$2#��/����=m��Kst< ��v{�;�33�fP:�E�<�OwW�����z����m[��ц��>h���e�}���Qt#�-��T-�
��k�=v��"}��F6w�~_�@�_�0b�?�z/!������7Ǫ�`ǝFV4�\�����;?��Kue_z=F{�2U�C�! jD��OX�oH�۰,�"S���]͐�(Vs���Ȏ�o]$ǿ1��ʮv45CLJ��V�^��^XS�֟}��v��yyBzV�������I�E�
[,?�0��"+���&`X���2��CPU�_`���d�M�!s� �;���c�H��6��˞y��.�&�C{D��69���;c���p{�ո���C�A<�T�-��;/���i$���N����˫���b���`k?�}m����}��83ԣ�[)��S�FV:�w��*+'ɗ��&lyl�#�� %3?p��	��4�9�pѰd�D�»�(]�3�f���_/I7ӈ�J�q<�z<��Aq���oC�9Njӌ��۲�o�Ө]��-m�A�F�r�r�=�Cy�.������c��h?1�'b��׬���O��WF�/ńC�ܗ��#��0R}]l���>ϥ�j�򵟟` П��prpg�� Ņ��>��Ҹ7{��w?儵� ��w���:*�;3�հ���ɒy�M���U��+�*D^<6_�y �u�i}#E[�[mKOA��i�Y����Q�U�geV�k.�h���H-���>�4�u�����&���"G�u~���ƅK������]F�>��h�������D�w1�\�+�#�g������]t�-�����x//G�pi�ң��`�f�/%����r8nI���m�ʥ�/�QvP�:rM���֓��%��]	&�]���4q"z�������<� ͓���y���K���P)�M�\>-�U�C�?3b	8&2��F~���
M�2��ZI:*5����'S�1�]��@�y�xቖ=�n݊�~���$6��]���v�.���!�[�?�׆�j7I�U��m�4Q�\9�c��t�*Os[���Aw�'��խ���={=�Y��n;���t�%^�^����E�J/��ŏ�H�K�`���#pO���c�`G>b�l�KA��+�y�/��~§eNv{iB�h�i��b�L}��3@;'u�vBXGq'j��5O�T�Xhn����,���;�GW���4t�|cU�.��e��������;���������9K`P��~.z���܇S1pp������"��8�.>�mJ�lIQ��J+d�;��X�����MF�~���<lt�h�ap���oP'�
�++�y��5�W<zR9�1�uj�,aenE�@�W��i���UMv<�3+8H�Pn�z�T׵QT[h�<�����ˇ���o�K���Z3�/eI����4�=�r�Z�"0����_&ɼ��b��PJ2����=��-9��[��ͭˈ�u=6S������co��ɌT=p����e��0:�5�4�䊡~�e������8��*�J4�����-�͞˯w���g>�~��婀���{�,M'x��B𠪘��|���T�/�e�<�y���'�Y+�Ś�����KMh�`p|��o�G��~J����z�����Za��f=J��x��v6.\��~���]Җ�4�����'q�B��-H���H������%��/l.�o��y�T��7�_�p�5ݙ�u�y[�r�|��A9���r5�ӥ��Y˟�|v}D|9P�O�.}P��X@O��K�T��s����h�O�l�u��Vy��I��������nvYY���DW�Nw��y(���"�WxH�bԣ&��>�S.�0���JG���꽡�r�yI؍��-����CLڪ�׻��e��;�%�ӹ��f]yu_k��� �S�?�S�}��|l��Q8"R[]�`��$��Ua����=C b�\�)?������ګ!_i؞����n��v�ab�-M���s�:����Gp�_�)?�(�	��#lo=)�c.�ؓ
��C�-���k��!=�/ɲ�Dݰ�Zi�de��������h�7�U�$Fs+LK�p�׮%Y�>�<�i�`�W�O'ߖة�f�r��w	�?��}�n��r��uD�N��3񋛇Q5&��l%c^]�~���qĿ3�G�E�-�14U�̋��Kĥ</8��;�\��H�wGL���d����!���=�����B�kﻨ����ca3��Q��G��n@mI���F�iO|��cY���Uv��~?�޷o�=�Rh���ˊƭa�`vR.��|�ÿr�z�1kV�Fc]�v�/��Z��]LQ�m�Υ�ߴތ5e,�m6D������sG��Hy�|�z7�F� i��e>����v��	0�F�ްj�q��t�l�%򦟮��W�<���K(4�Z?�*7����>ר�<��$]�����?q��[	���O�����Ĭm�R��մsC�ݖs`�\w.����O<��3W��TV=1�x�h���[��r3�7;����=h#;�|��Z�B@Z,���[;��T��ƙa=&B���+󢌔�w���[�&���2?v�g�u��)Pf��;�\��HH�A��I����wn}�ͥ�<�w���_~����ר=�DL��5����} k�-���%��6
�����<��7^�aIp!�ŗN�M�Û��׻�C|�9�;ą6sY�^���DG��n�f>�}���&'DC+��e�s�q�>��6r����a�f��+����m
x��B�U]C�]]iŝ�Q���v��y���>�ۻ���ޢ�ö�Q�>�udP5jͤx�,��',IaT,�	O���WzQ:��䞑:���ø7@��#X�d �@�!}"Y�T������}�)��V��u��1��w▝���Q���_}aH�G ���9�\|�!���X����r��F^�i�c-��w�!�q"p#�n0'����{��0��i��W&9g7ǒ�K��Hn�.#8�7\9"��Ȃ���S�0/�.u�o�(�_��<`�r=Y���je�"���w^��@���]V�0��4kHDR�����ݸ���{�<�ѱc׬�A��X(�@�:���xF�7`|;�D�P��2���̧�7��%��C�3��QM1͉q�|���Rv�k\-|��n DVK� 3����S��q�����#]��UAL��0���c9����?xD<�d��b_�Qo�E���|��7/�[�����ڼ6�P����L&�~��'e��-5ֽ��lc�!�y���OiL�}ص�s|"���:tK�]A��x�n��XZ����0��t�d_0z��^E��W�{MB�
)�^���F��o�
���]Ҽu;3<S��e�&�,�n�
���e9��[k{4&#�l�-v@E���a`�I�r=#H�k����e�H��`|� $ѤK��B1I=4����J�T��
<�u>�T��Z8�6��N�_ ���
�҄���Jꌕ�iQ���a�Q���<��J"��2v�>��G��T�ޏ%j5���q/���H?��f�CE��]�[2�zzL��M��\ZN��LHhOP�E�s��c�dT���{��D:eJq�$#���W�D�$��*;ޯ��Z���(��(2ɪ��Q�<	M�{I�jǈ��s��+E��{C�j����ݥ<2�-+��
�l�2�4��W����0�M*Zӓ�П�UK��6���0<�Z;���ΘV�I�ˣ��c{ȩ�T�|I�|.�/��~�#��k�k�+�r��h����$��2��-l�,bd��I.�^0�#���ɖ�J��L����fU=Β/����B�Yl��Ps�g����fj�=H�`�N�:�ᇝ���Od1h_���ɞ8R h��_���9���b��i�I�8HW����|0R'�-]:�!M��5d�(�iI��m*��Kz#�����o��H�
�U���e�����W���r��8�@�Ŷ��E����	�Q��ە�$���/ɺ+�w,���y��t&�I�=6%`}�_@"����y�-�V����\�|�	8��1�)�v��(��I^�>]<I���+�=O�h��ֲ���DH���ۊv�ws��ö.����Ӣ��l�6��y!��7��^��D0�gZ_wE�_-��RN.S�P�EW��oe��������°���M�L`�z{k&���U3W�(�m/�D>*P<�8�V'֘�����/����yC�6������]�e�yXs�_M�^���k.&Jb�2S/IX5�tt���-*�
ܲ
C�D�l�C&��~�+.%�oJ8N�[�
���g��h���_�Z*-��џ ���.��G&�V��-��[,L
���U	x��C��{�S�+,�7���Y�M!}�m���y�~�N�����:�����y��:e*�� j��5b��{��-"k�Gz��C��4���A�w��«�CBR�W���Nj,׀V�-�}bS���8TmD+D�'��(z�����
�N�.�IE`��W��Ɋ�9 ��ؑ��I��W�f�,O~�m��825è@>¡s��-��ֱ:*Q�2�`Ӵ @�����q}�'���!䇈Ta�7���E�~�?�yn���q�Vh��g�\�;��^��DN�d��c߼j��kA�Z^L�G�L0������]p���1�,���Xh�Ρ�v�����mԓ������Ԏ��{C�1mJz�nF�:DEe@�(�q����IǨ���p�۽�e�~�Z�U��׎=���6�!���d1B:.k N�[��+�^H�Z�Q����a�Yu6�\OҔ�}'���Tܯ��Yϗ� �^�ԨX�>s�}��)s�b:�v�݌pf��\���<t��MvM�������%���$uCX�9��k?���<�&YY	���xu�7k|u]ɤ�֗.e��i�� ����^����42d�[SЭ��;<�o&��郺��˨ފ�cd�e���'G��b�X�c���$�r�ku�s���e��y��u��~��~�ֈ�`@��.���pa"0����w�q���1��ix$�:�[����Z���f�o�����OEt��7�D��H!�(�k|a\87�������~�8+�n�n�E�E��*^^�z@���������d�r�"ć�T�I�X�>���=�l�1��G�k9c��^�Yd,4\��ښX;ʧ^�E'����闒�2=q'v-V:jF��;�Y���|䨼Gs2�M�B��r(|q{SZ�J4����auYZ�TP9�+��?��5�u�����|{�����Bq����+˰%�����퍜3�V����|Cim�^���k�s��镛n�b�<Dza�T3�")��Tq�]��
����[�+5��ӭrC�˩��/�|B�#��
��$�+�	I���ߖU@;z�#VN�=�9OJV����)�2�M���j�_�Q:z��d@g���bX�2k脵�W�]W��ep�ا��0���]��Ӻx�P�g��M|x�wLV̓�{�+j0�����vJ�փͿ��ٍGh��Y.6p���.�i���,�GC㕽��:آ�P	<0M�}�a��X�#.V�"��8BkDK�?6� 6�V]�l���T�&��/��h���=�s�����TXIݬ`��[1쳆�T���a஝���V��G�>
�zt�`�g\G��o��7�ʊ�ah}WpK�j|����yS���'=���ɱ�[,H�NW%YF�eke�K	���-!5���	�繖N�h�1��3���*)I��'ަ��W6�����vi��H���W�f~�O�����dv�����lEuj�b̀�.�UqPur�_
ͼ:�^4G��Eu쿶���<�"=H�Ɔ�Ol���~�Ã����v�D;�ja��7�&[o+Uc���Z��xdA���Q��n9?�i�t�\jF~A�[��^Rѯ+n�f��2�e7�|:�Yo2��%{<_��TalP�O$&�N�� ����"i�W [�φ�\�i��.ݕy3�&�P��.K��Zr�� <X�4���P�6��u���#wߙ�6����D��i��;{����_n�'�������%�J���[�y�\���(��?��>�@��b���E�kKa����V[���s���
��cp|��F����OQ듶g���,����96\��	��p6�;om�]@��K�Qq8� �{�)Z��r�5�S������kw >�P�֞���z��Qd�<^KQ���}�<1A܉����Z'y�I[�?ΓU�>�?R�շk��4�ޫE�$ӭN����ME[ C�#5`6�'��� CW�${��[��i=��x@E3��z;wn�%C�HJY�#�������{ �C�M5q��RԀ6B�`3�0	��"|��Q�_lYȊ��E4�]y'��K�H��k�����,����%n/�p��'��{kx|f��/�x�E)��F�cc��4�qȚ9��5��'����r��O*��]6,<<�6��?#���+a)((�,�ov�d�h\���3�N�I�!5�xA^ ��z���T��ϔ�bX���PHc�ue�u�gơ��=��>�а�m��Lb���7��7]�
{���L�����T(KO�t�s�^��N��?*���zR�,�]�������e�����w�N�N��n��-�Zq
�V%}��4_2z����7�B�-��2B1���m����A��N�y���W�μۇ�G[��㝆1�g�Nhph���g�l �㪮.EE37hntFxU���K���#��N�_!wm��WM�>�ƀ�CD/'}Y
���_���&
��|<���hQP�((Ko�!0��x�P���8�D�,���\|sR����L�a�m?�z6k�v(�H�!��=9�2�BJ��z�%�(�)'eG��nj��YA�F�u;����S�f�>Δ�7OQY98b7��Ob����<���1�y�_��?�u���?�%kV�L&���l��^�mM��Q �2Vh[�P�rn��,�T9-�B;i�W��	���Ѓ��[�	D�uԘ���Z�_��5%���"�� #���..bMH��)N6*i��5b��d�����긝-'\S�8��3�˼�BqȘoQܶ���
��?Ca)�ћɎi�wj���M~׏5+�M�꡷5ܞ6�|w3H�}��!�c7��aqR7��>�ٖ�_��7����C�_�+�4V[k1^����C�j&[�Y���#���ѸC�z�.L��<�����Y��h�a�a�����t�JI�su��u�������z~�H �@�ch�ݲ" �|�vI$ٍ���MzG�y����7W�aNb�+�j'1�^��S�Ĝ�r����9��o��VCs.���F2��+).3����g׵�9썌��^�@j�/���K�p�I2%����:�����|���8��,��AU�?m5�ȗ����@+*�)4��PMnk�E�c��5�ߛ��5bѤ���  j�Zc�۷4�#��ff�&Nnq��x�G�dN
c��@ �6�2���?�nf�N^��2�/�(���{�l�3OSsO�x|-����=gd����̐qss緼h�)@�.���5�	�kv����Wx���m���K�zMfVHF��$ŉ�]�_�n_�D�ʵ�=M�FE��r��;C`��ͥ�B��U�[�ʧ�����@i�O�gMY=��ݴ�/�ÁJ�q�I�}X���-��:�=׾}D2���h �D�A�N����m_~vxFWJ}ʓ~����b���!F0}Y��X$?�b�3UQ��?TP������]Bh���p���񓺤g\�c;��lH�-B6S[(�P�;��x<V ������Ps���p��e��뼗i�`��_mI�C�ZC絰�5x�[`W�M�볞��|�������j�<SOga	���Y�E�k��9�s'�"�=�|�#��V�yv��.Z<���A	3f�~�k���=��¡�xH��H�'I�e���;[2��;�m���$HcoG�խ�+��\�����T_9�ayl�X���? �H}>A󹵂��l%1W��(��Oj�,G=I�ZjÀ���]]��A�u��QݼLo��(��M�.y�^%a�?I�ۘKC�ܢ;gD\=X(Ш��Ο���b��{��'�o�Rҡ��-A������f#�;n^���<�~��Fm;*��&������ц!�{f�8��WL�C��3a�O����׸�T��)�վ�Z�%�N�M���i���D�9(�l��f��9v��������X�Ce3_��or�7�+�ʟC[��s���Ở�c�������f��T�	Qg�8-9ݡ��&:vf�k�&�Ɛ���`�E���V�le�e��k�bRgGѲ��B����Ј�ac�nx�^^�Vg�����`�_8��O�#�r�����;�1#��'�v���o�|�G+�&��F�Y�.,%,��������㤆�(\���)�o��$j^��W�7��I��4#Y�tBν��0�XKt�l���Խr<"]~w��^�3�u��<)Y��n�{��F��>����4�[��i��>
T`��8�>T��E���\T|od��I�����&|���Zφ,���;t&�"�uC�m+�ϭ9r���Oԍ���t��)me}�v_-O%���槩��\��R.6�B�j�F���"���rM��;�^� �
��[����jR�	r�zۈ���s�G�\L"�D#�;\�M�d[�n��.�D=	)��f�,�b�" �=�vFQ�IB�Ƞ
�ÿ$��c�~7O6!�&����褵Iڴ������!��p��O�~pív-Y/3��ea�N]��STn��-!A���h^{��h?�Q�R�d& �`Y�	�jk��������Wr��KU^%���n��b66m���5�4��t9.����g�C8�6���d�Nˤ0�R�g�N��b�
��C�(�\(�ޭ8���HG������B��}Y�6��H�ނ|�2<����)�m߁�ܾH��oF�t:]���E��7�]���
�\�rw�*P�$�4��[r9}X��7=���Ы�-��y����a��9�dt���D
 >�3�{����0�7_�@J��TN�-�6,��4�G֞]�	}g��p����Id~��q��&`O0�"Ae�!�|�#A�\p�hB��\~���H-��|*�Vf'Om�N��e��e�>�i?�9��ݳ6V<]�P�7�@�}��FQ��M�g��/�'Q�/r�}�����1 ��S����8�P�u�Ȕg�N�0e�5�? o���ҡA�o����,��<�!���'T�������8G+���V���=A�S1`�٨��ԩ�ʱd�\F��"#/���!�_ڰ8�Zz��3�s}�>|�y�F�f�r���c��gz��V�
~���OE  ����aRjK��7(H�ᔲ��s�H��q{C!,����I�������Z�x�¿�*h��r;@l譋�7�'G�D�{�2�fַ�ć���j���`fe�٨y�q�Ə(훖�t\U��vTR��P��?��s��1��r��U�HnN�
,�����{�uͰ������k�>�z�@e8�|2j��7M�����a4i_j?1^���HҠ\ҚB����[�#��0e ��55	����/���$^8�<��ҕA�t[�����_�[�MGF��v}6�B^Y��xq;�Q(�(lt�wb��#�
�J1�j�α@!,�)5�|�Px��'��\f�W��AE�P̑j�o����$7�D����V:v���h9iO��fA+D��p��f�r}"����,�0�����~=Q
yS�ST�M�V��/yf��"1>m���ѳ\G��H����F����1��/�N��{:������n�$�v��Rם~Y�i&��g��+�����(9��aq�4�?{����$��v*�����g���N���K/o���� �Zj]�8�(?@l���:��a�D�4]&>��sE��Ms�HZ;U�C'A�ژ&���(��J��t�M�CM���"�J�fI�����;�.����fS8^���H�<l{��<(V3�� �i�����-'>�E��P�kf��O*Z�@Mc�<s���L"E�+�K�h�[E�-���vCC*�hqi'�3��]Ɇ�8�p'~�U
�����ˋN�1���m�5E���7�/�%:V|��;8���J`�	ҕ��:��.w^T\T���:*Q�}���-�,����J)k@��H�IJ�x���D{K@�����"�\��{�`�����3B��?i�u"�^�:�+6q2�\�]��3g��%�K�i,�Q��ˎ	���GCi�����u��I'��v��Vhߤ鍅n��@f����F��m뷗B�Q"{�+�*���%���T>�L�ʘ#��~�u��u���B�G��}jG��Osp���nݶ.�aU@ZI�3ܝ2�c���}��&���U�G0�V!�����ħ��7�J�S�����]�"��r<�M�YI�p�:�E-n%V�ͯ�{���r<��g�M|��ԏ̓?���ǌ�2�������G��U`���Z�Z�l{�#�_~uF�{�����j~������N��;�"�����-u��!Of�Wy��3���V���=o!__�3�o��ف�?�+k�]��a822$<�J���6��c�e�K_����&1��_�3��,����1�	��C����Z��*;-�ËaJ�������@z��`G�H�@6�]�7ep8<v"ƈq�YD���X.�KW��$��9?1I�TCQ�e:v����惜���0�]��m�X�p��n m�dH�+��a6�/���>l{fQGC����$,��Z�K����bR��*��@�w'nF)$O�Ъc2�O���xS4ζ'tk���)_;{�÷�C�A����v�ga9�Qt�+�D��qw�
ы�awn�[�S����b2S=�gů�V�7q��o�6�]�,�O�BL�|%nZJYU����-i������/���g�Qԓ��y�::�ꮺj���>;���;g�V�p��G����`��2Zҫ���E�Ya���ƙ������؂%.=܂� dp=�A� i�^�E'� ߝ�Γ��i�Oߝ7t���A?���5��ѪǗ�OHnL���:���1�In`Qps��D/Ğ1߆����6�?��X慎�ݑ]�������.�����HU=���e-���}\ۀ�抗kX"��ԕ�0ֶ����$z5B�+�|o����-Y&aźԳ�� ���z�z2��uW��QHL��/_Z)]��@Nn��E�=up?ؽ��/����k�5Ř7�N�#7�L�f���`����x�:	�v��\]T���￷ P��ne}x�F������� ���>��;��2�_�9�Խ�S�����q��[�l�j�aҬ�:]�a�C���$���2��g�t�B&�5
�)魑-\���q z�X�fȿ��j���cwď�\W#�p��R���I!����|�8�˟�"�x���ˍ��>������S�T�MC�~��
���
.�E���](:�T������׳*�q΁k��N�&�p\�����%���<&�l�)5/-�V~�l��5��i|��\���zF+�C��d���ޮ��x���^��@��H|��X��#|@�d<�����u_~h�ʹ�_s8u��X�o�yu�[R���������֦u�M��v�`��f7�O![ݫ��m�����bk#��'h�C�����J����n92�l��N��#�4�[����_A�����ϙsʟ�8`��J\NuU�f']�&-}Ɂ��b:�����������zN���+�� f (�x�f��D�ןIX6@�mbܲ�� �X��hs�#���i� �(O��9�\�|,�W���
��db_Þz����.�u�G�Gu�����Xf��$f0`�2�^�dw�߁+zެ�� �����;^lܼi�/L����v����=*���P��-�>'�/�fy�3p�e��~hGQx�ǈ�����a*����Id�+J����GjN.Md6c��|SE#˜�	��>i|��V,����!0�������C�j�,���W�3��5y��4A�CA
��h�j\Bc�xB[+֑�\�s�t�Nz�BZ� ���c�V��]�ʿ%Y���V�!���(��8	j�^I��!���!f)���敘��H���%ob\��E�%��^_ڇ:���V��ˊ��C�X���w�v���(aG���N��-��A�+� �W������ϸ���r�MVZ]��G.�M�st�h8tx����%��&��Y(�0w�~����#74',G�����PT e�q�d�kt>�Z����;LKy$#�g���ؙ��yRL�p��zW)��":S��5�X�ل��Ӂo��~��ڠ�^��� �n�X����� R��Q}�� �&����	�k��ݕ��N�(�Iq�d'�C:���M�M�^o��b�L��S�B~��﮲�W	=5�܈07�������DFH����~1�kf�.bx����%r�L��������i$����l���`��������q�S�f�QȖάcB#�|,�.�auh��GmYf�'sƀ��̘޲��VϿu�+��������~	i�jm�,�]�
Ԗ�
��'�߁����٨S���t�j��|��]
֙$H�"�e�A"�.�g���*BGh"w�_�,��p���Q���o���R���A��"ۆ㶋�l`��gP������N܀��0�ҩƇCkE���X��e��?�^�0��s����8�8�T���O��jm���M��pW�����pf�t��r�.�k�%z�"2�C�?����d8J+(1�TQs�w�}�k�+t:�de� ��T\y9��bC����\f�Y�u8c�}t���y�p��IIL�+��^i�^��Q'��H�D{3�����+ɾ�i*z�;��ޜfMVCKO;�q�����_��S��%$
��
q�5T��q���3#H�0�z C�{'���0'b�AZ%��7��9���yVWP�تKhG��IL�`������v(]���qN�T�q����WuD�Gz�k���t�9q�/~B�����4��)E~���j����$��>_�:v�F[jSNj���%'s��}E8�1��0��p1�J(��Z��m���%�����Y��::�0x˭�n�0
�a��� i6F\e�G�U�0��;<��7?iꜬ�|�����Ȍ.��9.*_;g�#�ߓ�����ff����i�j��qcǊ�-(y����'��Q�3~I�S�5u7j�Se�a/����z��XO<Y�$gh#�X���h_4�^��܌�-2}D�jZ��tS��;�j@��&��2���&�7�V�x�Ҟ���DM�Z[��lh��|ۉ�� &ΔP �_p�v}Px��)?S�7z��Y��z	���P��aÊ���.֧-��X�ߑg0XS�~O��}ف����D���������E��Y��v�1��p�vql5��6�5�	Vp�##!!c��G�3�{��kIF:Ϣ�r�Fbd*�ur�{Q9�h�&�?��-g�{�{�ԁ\���'Ea�q"�	b�Eἱ�=�!2�>�B�X��;�B���ⅰ-��' ߝxg�|�����f��Â7��~��`�x���0E��W��4�?���6�8���Mq��ǯH���h�A����l׊�����V�Ƃa�W��k��P�b�M��5Ԗ�F\�鸁���N�(���vx\�V�?�&A�b��R�1k��e���oR�e&�3�m��,ؔ%���Vs̞�65z4�ۄ�ܮ}��<�j�ѯ�@�|���;��5�gϲd���f�6��3QU��9�ʰU��ģx21D����	T�xa��҇�)LhV~Ve��Q.��g�f��<�߹Q dӘ�K}���QiX��xH[=Yj�����?����到��-k�9ŖܪU�]ܚ�=�ϵr��5�j��|��2T1����Lʅ]��t���"U�U#���~�5E�;"��~�jܴ`^Ə����m�њ�-d�mUx�j����si��ف�5To�,��`���%`��Q�u�,���O���lV��1��|R%�t��T�W�/�V�I$��OJcڋLsv�x��D�#X����xK��	��&9Ari��5�[g�Z�ܪC�����+yYՄ����H8����M��p`7FGֶ�1��樨
��υ�YʾH��O2�Q�fY1��Y4�I�x2v��D2�vY�| �Y��5�k2�F��*(�" ��x;��j����>�ۃ���2k8�Ze�Ӱ��,�
����e3n��Q���[O��2��T���G8�������\�L�"������O����ս�^/I�y=�[˄�.��x,���B��C�41����iK/	����&�)^r�u��췥PN���:$p�y����$fGV�̛i����
Y�>\��ۺ|+�Y"����D�뿩�v�UVsȨ��#�ݬ87�Z\�����H�=4t������8l�����ֶ�0�cY~sB<�3����ı_d-���x�)ٯ�A�d�3���F�h�&�ɬ�*���z�F�����@�gl)�C����ܱT�֚��ϙ�c�G�4��V���O�d�+�~ &���/1Ü.������ʷ��x!0��3�L�E<�$�*�&5�=36���t�*d�+'�ٽw}=�8>v!����+Ƃ���g'Zg��1=��v�O��n!���C�� �-����,���o�ц�Չ�>�ptuO��yL
H����OMˋT��9�kd�� O.l�=dkHG{ jUզxt+i� r���Q��ҭ{m�{��������R��Ǿ\iLջb��^6��s�#��p|$p-O%��`��3�tɏ��C8�u�`���ل�uؐ�@s��Z���2z��9o�I6��!�:��X10@�P�'!���ÂN,�\cE�A�w!�k��A}���u)�i�b8[Q��X~���˲�u�	�y�^����g�d��Vws�U}��(����t��+:K�n��*�kXN>712v���:��l6k��u��Y~NK�B����v���T=-vf�p?�����������r�Zz�J�<���\V\�M#�m����Q��F:��V�_˃�=�>1gF��#%L�X^��s�n�@��~����4cs��R�H����h�C(_I�C��'C��m��ez.�XV�4����J�g�k�je��_�ׄ޾m!*"ҥ���t����HJJHF�D�.)���"ݝݱ�	l0���y~���kw\q����t��]N���oI�5fՑ�Y�ӹ^������_�����83<S2"�0�z��_ϣu�h��Ok��K�V��!Y/��gf �8���D"%O�5��k��%&cv�-�y�'E�)aF��b�8hZ�`/��+f��W:h,��#�8-i�����yF$,�C7F������/��;<�[l}]!��)��[5�$�y.�2�]u��{���^�h^�X��v"�+��ǧ�M�V�8�M?�h�b���'O�W,�,��ݷu������x��,!�_

	�~�i�qE[p�x��_N��=݉�I�S�����b�f��h��%�8 ]�z�L�/"^��*u8ZF����(x��囗wh��(��A��n�ܐ- ��I�Ӫ�n��M�?S/�?��c�y�s��Z:b�:�2��Z��3ّ�[��,6ﰖR�m��S�{5X|+��EF=��y_w*�}e�v���[Gc��XX�E�B��L�C���\ԡl����%��z�l���㤘�{����ZO��£ud:G�����'(لpΈW�N�e
 ��_��h�C�.��a���e��I�g��t��kW��g����o�@o�]�o{�M��R�_�x�=+T��'��&�ѼiFF���
_�b�e'���D专p����$�7�������e��.f3-�_$�l��6A>�hצ�����&z=�&|��Yw���9To߼;b�C��#��QM�H'Y�O_��J�<�����[��0
�G�|�������Ț0D/ô�d�~�/�5G�^3�z
R��1�
H����7N#od�Gy�y>U�@�|��"�i�5��yY�䇆qO��~�eQ8�;��r�	s�sR�y+��뽮r׶V����&�:m���I=l�'�-p�nUu,%��f�b	%�uI�/>)O>����{�j�9���a�����c�'�1�9o��H�t��Y��2�>qE+U9���z�r-����@M�O�q�ˎPB[�����l� ��Y#���iGk}�[=b���U��C~ARU�CZ=���&K�h���[����xE���r��$����1u�e �oك�(�j���'�����D6�c���J�l��1����irC8_�N �U-�4�;�f�	˒��p��m�c ����'boŘ�i�f�0O�B5تJ���Hb�aE�;�	z2�?O�5LC�6�:��ɣ�ɔ5]�>`��H�b��r@����O�m�ܳ��W�fW!z.�mx�����u
�C���Otx�����=��v�����l�Y^Ș�Bi��DR�/w�Fi)�$Do�����>tV�y'����590ç(��録����肜�Y/�卂���Y�];�V����O�G��V;�Hd����C)�4;�l	I%Z��Q�qUc�HLa���?�_�e�=Ah���)堋��HK���Ep]�K�5H�Pd<5�;�k�I�J	;;qT�V>�j!��;��}��!��o�c�.����w'C�Am;�h����c�$.����|��1�kxr�C�l~��w]�ֱDkV:��)��x��Z�����慪��m}�z4]������9�5�j�{���dmHOȄ�|$*����ތ�]9͸���"����d2�+ck�I/
xK��A�w�$t}l����f����������n���Cq�7n:	��g�O��=R;�؝�ʹ:Y��1v�|W�T����yx�Z^����xqs�d��-������]j�7#�������S�!��^z%N��j�ٔm���ڥ�H	����?"��G��j#jp跥��2�L�QM�r��Yy>Z����va��Eb�s��9�4��G2d���u��鏭�ą�n����\^�;;�F�}6�t+���E5Z?jTJ�x�`�K)�H:'�(O�.��7y14���Ι�*u�ԣ�W�JX+��L���k7�޿�JA�D�����@�d6��h�`�Wj��b8:Yݶ&/��4�$����gdWy��>��%pV�����\��BF�d	�d�j�r*ҁ��=9BM�s"y�+�L�Ҵ���p':�T�O��8Ɵٸ�)H{�=��=��E���Y��͓��Q��w쬼������4�"[�p �O�VoB���#V<9���rPf�����y�سT�|1?)׬���?��������[uCc|tc�t��K�ŢX����lX�Ω��P":�"���yHL����֍Dje?���0������$�Ug6ٰR�aR�|,�֯t,��ӧE�ku�-���������QN�7��3�����&b�o���x�����h�d� w �2Ր l"�/�H֏�׬܁�F����B���i4S��n���i���������\[�R�y:�H�)������B8�Btwf���>6�K&�譠�jF;l.�������֕�n{��fz+�3��*�����#�۩�\>
 P'��h�Ͻ�s�d<P��(����>6��y��<?��n���翰n/�˓
��ͣY�0��+�)I;ͽ��t�M�����*�J ����ũ!U&K{����
�E�/��K7��*e��e[GGqy�x�Yff�N����͇<z��XU�`�4 ���.�To��v�כ6��]��ZxJ�FK�Ve2��!�>KM���.��2@N2��J[�=�ސ54��r���!����1�
���dɝp���j�=�UH]ޙv''�<�e� �R�O֧��D���-m���v�|��Yg��qVTm�����롌-9�}�n�@����I�ò�7kVH��:����صr_�e|����~!�ו�-+wǄn�]-��3v��E���'_�Ew8����gA�'� ��~�h%�QdK�j7��e�dN�XV4�ޤ��O>8~qE��6I;1�m���5sz��k �.S��r��h���'6dZ�x52LO�Ȫ�K�[�X���3�'�����[}��B�;���x�>���ى,uhfQ?��u~ߏ�&q#���*��j#�;���<�l���7N+9����J�|뫄�bvt^j�Wd�H?
�h��
FF�c��n�<%۰��w#��F;׼s�q�Z���E�UL)Ѳ��ک��L��e+6����C�$�-M(���y��<%�7�����M�qK{V�DVY܈+jH��l�x�䅈���\��L�4�ܻ/x��^_o°o�?�;0�o��c<)�k�3ɑ	�^E�qme��$�k`�Ih:(�J#�V�l�M��7���L�ҩʻl�|fXd�;�Y�&��%�H�p2�a�M����=�|��6Uuϋ�P�����ҋ�s�+S��oE��@<v��\"Sb{q��OܿO�n�ݏ�r?��<�l,;��5'
�2�����6�*���䋌�2���CI���}.)f�9���x���M�`f�4���������2��P�5��������Z�x���"�^�08p�/r/d�E��Ґs1����bff�!I���=�ў��\+�S�g�T�*��˕6ʀG���^klE��.EܧL�(�R~NE�0#�ɕ�Q��A��k�w��V	�<�(j��[-���I7�ɲ��Nu��r����a˨�/b�q��l�/���)�!D<�[��=�Abk��ǜ}���I&iI�v�?�)�;'���s�Q�]6Mh��Tv��'�q�)�}*�T%~���EC,`t�f������&[�B�/�<a�;�;("6���n���!�?�oX<��
��أ��:���ph��c�3o<��_l��^	<�|�������^�5`ڣ�
cj�?��B��=���sG�0vz�q�����.fa�)�y�F��Ot� *��mU�ג�L3ʈW���n(�1y�S�;����7v2�f8�����B�Lbi��ؗ='��Zv+��U��Bz��}��H���o�P�Ҳ����=4͸?o�['�F�L@�J��2�mvh�j�fљ�����:����4q����]}��;&��� n� �k'w��iA7'��U	��`�θ՟���κØ�3�7��J+7�7�>sܸJk7�@-�v	��5k�2S�R6�{Z��{�_t��-�4lk�r��3�|��#r��(�V���E׻k�3�NO���z��I.�?U���嶦Z���zx��ޔ����~��bi}l!_t�Rg���t�c���uZD�Jt_j�dȮ��8�X��Q�m�k~��{e�3��w���:�2�]��Ӡ�쐌QL���Q��$J�v�P���\Nث�욒mP�S�ڏ�s"jN��Hb�LS�x�l;ZF.�I�y��4?3��A������g�9���~�}�w�E������?E����3��@�n9)�V������W��5P��0k�=M��Ԗ�J���}(��brЊ�t�g�A��<�)��;�A`���ؐ��"#¢��p!2�C%{�Ù��ڀ?zL�����2eP5s�y}g=��z�)�c�O�����?aR�"��	�/4�_��z��3�`k�0�;�@-Q��V���|5� ��xN�gG�H��ϙ��3��	�Kh�D�lZ�8G�Cp��`��t�\d<��trh��h���rr�[9C�$c�r�tJ`�6���hU�`�lU$����<���3�Μ_�z���p��Kt8H'�v�<8��6�[�I����֩�H��'K�PK#(�-��]��;bM�E��eg��hVF�G��S��g�MüQ2bIƐKR3j�]�¤O1^4�~���X�"4d:�W��9�r�/�d]�"���/���7�^�t�K�IOt�i!$�L��|.��C4����9�6��5�����]�?{�,r�D�!)��%��΀uǺ��D֬T?Ǚ�#ssc�'f�����M9iܢ1����]%�B�R�)~~�g��W +<��z6͖�JNԨ�ݙ��8�#���ӗ����`(�[��zqlEYk�	Gg��w��ky�wnn�V��?�����hf�pM��,�:��_ժ�4z,�$a�$��euqFH���~�RƯfĒ�������!/�$�LRy�)�p����-��7�k�Cm+?���ޚ����=�2��S�a�ޟcD(���m��z&�!k0�J�=;~l_V������ �|����U^�C�lȆ����@d��\f�Gi�iȋ�"���W��[ӎ9���M)����P݀c޳����>�{+�(V�iɨܰ��iF	��#�����@�d��}�ߒ�3���#s�Oɏ�� Ad8 ?sk����1���2#�-q۩�!����M�C��+��ă~�����%B���5Oh�j���Ƽω����<�z]m�U���e��,�L��8|�+h�9��/cB�/��M�%�Bw�W�=mY!'L,�c:��V�1�Y��i}�EF�5����wm[��ӻljT��!m��ӷf�e�Ǧ^cTLj�x�%�4A�>2�N�ܣN5����7�L$~���D��F��	J���7'�Rlށ�*pӺ}���}�(���`1�n�ɷ���/�	�یr&D~�S��
��[t�� ���6[b$�j�l��珞R��x��%3�k.�,�do�&���L|��g�>�6����z;6���4�~2q�#��>8����c�/�3 ��8�o(��Ȩ��!eu��J�o�w��]���ރ�}�߽�>�m*V�������MD,��%�3:7LX�� B��`�������Eѭ�c�y�ؕ[ѿ��V����C�����<�[��bxNdhOE8�8�׮V��Lg �AG宺�%��§�/C�,�e���M?c�hR�'>w���G��lwC%��;��<|�z4}P�<����*�]t��C�i��>����4O�V��ʤ��E�-��E�|����>ol�:C5��O�e�8j��J��HzlCS���ƿ��cA�/ �a:1#__+} �}&�X�S�D���	@�4�O�̽OL"�3]նb|DP� ��+�
�[�=]d��c>�?,��}<J1]~n���и�'d`�s����ō*J� �ou8]��1������b��m�U�_�8�x�u^OS�*uw��t���'}w�N���kڹ��|tx!����x7"EiF�bX�&��Y�������x߄,Cu#�:R7pHh��hv�� �r0�G����fx)�Y�}D�y�ǎ6rLҵo���Q3�ó���_���9sʨ-����7lV�"��?6S�}�i��	�Jӣ�m�$�:���������j���!�2%z��U��Òxu�˵x���Z}��߃���E�W!9��_�J>p�d<����<��֩^�Hj�j�@��@�@Y5%`��HG@��o$c�ِA���'��k[���;���$��!�h��'�s���a����$�p"<�D�@���X��-!ib8RX���������0��bE�BZVYH�D�mG���$�R7vѢ5;������x� �};f����}�W�Z�]��0G<]$̢C�������ރ������{�H��yP�-3����!D��w�1%S$>a���t�T��`)�� �U��˺Q�5�̯&a8�:��2�6���q���'���
]�i��o���V*��Ђ���E�.�[�@ٍ��-�o
�2�����]?p�(q����ߗ����5d��S����Si#o|�	Y}���y$��Z$q׃)�{�rkQ����۲�>s�%�?Q%�ė�
��@O�'E�kW�[v�@C
b`��]�Ƕ���w�:';k����IT��I� m�Ug'�hچ����5��3ߪ�|D�U�[A�������[���\�ڂn�綨�����k�0�A�}d�"C�}y����B�fvS��
�4~�lm�&$X�>aS�x�j��GKèoN�h�6M�\})B~ ���ƒ6Y�J�j�_`��1"F�7�	��Hn`	6F8�_Ԝ8��B}�ӧ�^�a���,��&�%�>��)L:�¤f7d'W��Ɍ��}!��o��	c����6K���M|d���S>B-���P0G�����2v�ҭ=�4jSi1�d���W,q�&�dV����q��S�Nvp�I6n��@Cr@�������<Y���"��c4�#FlG�^�A7}�)Y��1z~��ڹR�X�t�Ǣ�λc����ԝ=��W�Y�8�*e�e>~푌 z�R1	��׻)G�P2�ƨ�������N�#��!_�O�x�r�	D��]��Պ��N�%�[k0tAUo���� ��6`�{,���5����`�_�W��}CZ�prݴr��ݭ��q:]�
�� �u�"��S�;o�-X�����_��'B[:��\$9G��
���u�F�x%���Z�}8�-�]00�T�J7v��.FB;�A"=�������zc�����OŦ(��o!�z6.�0"���=py
�J�d���Кjj)�)l2Do����/��FC�HNa���vf*>�Sxe8 �U?��ס���/�#���%�'\П��e��u>Y���W~��I���,����'$��~���qu��O���RWw8c�sZj�^�Ԍw!#e���	�ת���u��՟��?s"�W�jciЭ���YP���[�-fO�й��|�61u���-vт<�B5'z}���t\�@�o�@��U�%��//�[so��+�����$��i���X㚠�C�U�x�U���#��c5цg��7e�ň��&�`U5�<�3��>�p�]("Q����c��Q�E����G�7���Y����Ao�@2�<al]�(���䒖�^1_��'eW��`{i7������|�i(if�MAl��<��˂SZ����(���}�K����bG\pJcG��E������6md�K�����&��uC�yR�B��UJ�#E���M|Z?y��� n��vM!i��3�"�!�}�#��[{��{���
��ە�� O��+����r���+JH	��GT�(Z��ؗ>�U�H���-J�3B29F��ȢyP(���l��L�.5(D�<��/�lT�_�D��įzs�_%!�VƝ����s����{�W�3�TmS�Vz��co���kɦG�խH:���	?'b��|}#��r�y�&�4��^7;p�,��m)8#t��l���kkl��r�ؘ? (�ǋ]��b~prrH������уw�k�Mk��ڻ\p���h��2������O��waG5�HJ�伪)�I<�p�p8���O@	��2��w�l���-�g� n��]��̄g!��&�7>L��fpM}D�4�6�.t�,��K0��-�+�ʼb^/?#>�ʛ)ؿʭ�<��gYx�g"ޫH���F�Z}e�� 6d�ƈӚ8VB��f���ҟ��F���-�h�VM_k9̿DH
��HM��O�i�:����3{$*��޶E�E�'`��9�����Q5h����5T6�AZ~��Z��Y�X8NJ��ѳ����ٮ��ʹ����B��g�o[�Q�#�GY�Q�a��(��u��O�L\�>r�����ٕ�8��"S���������L�_{�c��<�����A�=eb�^}�F'���D~>iM�N�CÉ;�-?$���Ђ,l��+�O|T�bdM ��ԕ������Z^F�(��鷥�$1t%�Ǯ�15�ěo��yoe�	!�j�f�	H�i�%�ڬ�+��yB����wOV���#�o?p씱�+�|ҒH-��G����a���5�w��[>������G�z"S��|߇�`ZYg4d��W�����i2�.��&O��oI�ZU�N����X�h6.Y����$��[�Wn����lKl�aΠi���.���S{�\�Ja_����$��	�ܕ��@��s�
[��o<���l@E���!�դvH��nɸ�>��[?����Kk8{�����lid�9�|a���{���t��c׾Ԧ;��,S�7�48�L� :,�#ټ��71�7��zG����}I~���?�]��ԋ �"t�W��� ������&��ETM�^~�D���c�o��B��3gp������SAh+8��'���wg���7�����B���Sm.�@���Ӣ�c���a��8#m/�-��\�aޫ���\Poy�jۗ2�D�L6��P���N��WW��y�WD���:&OQ�'�C͒%�r����s����۔�i���˯�tp��Ҿ&��>����R�}���p1��h�6���l8f�F�z�q�B�|[ܕ�mG-!����]w�K��G҇����}6���d���ګ=�]_���jN�;��@(�i�2�ۘ&�g<EH���w��2�ËKٕ��S~��Jw�ٕ�!�fE�����G�[H�oe�M'����d\N��q�S�ĵ6u�r-��=mo�V\�yџ�T�N����	;p��#}Hzī�V1��)^�&�� �uwl��0�5��1��VEF�w�l�7������&C�3;3�"$�]��^�&ď�ѮzF>�x#2_$9� �q�\5xWy�@,T|����y/���)����)�Uo�S���,����n?�B�Lu�n�����p�^{�ݰ�PEa�b�"Ta�<��8ʣN�v� ��PԮ�%~QEK;'�ٛ�N(�5�E�������H%>t��c���
�-"*�\%;lONҮ�T�d�΁ O���HM%�IMZ�>�&D��w;Xn�M7�Lт1�v�*��Z���G�K_�N��w1ۋ7�C���2�$Ք�g�0�ͯ����O?��b�kK��-�EO�VJ���̖[ٟ:�F��������#(n���,�� 9|��E]�O�Y4»�89ޙ��Ĵ$b�P� up�E�^��r/ ��|ڶ�%Hp�?�(a-3�֋�3x(Y�Ox��vX�Jg�gN-�R�I$uYצ���t����M-��(k5�����oǖ��6̃��#�?� 6�Ix=�`pI�zUZ~�����~\�6D�l�3��)c�J�Νi\"�t�L^a�M��2Z袰?3���ѩ�<ґ�ƽ$y�0��/9S�M��z�+��J�)o|`�Q��m��I������٘����T��<_��;�u!��g�ɠW�t�[N.��x)�qnn�\�=ZD�_`��}��f��V���s��Wt����yf��(1�-�wu�⫽d���##d�ᠠb4ͲI,-�UmJ̩�>a�lsy!��I��ֻ4��S̭�FD����V��%���4�,�ر��(�j�j����0��R�Z�A����]p���s�#�!՜�:�:�d�[��{͖�g�V&7�P2q��a�L��}���ax�Ǵ#hA@h+D :QL[�"Q���D�Hh��!ar����BOO ��R�B�Mu\I9��N2<���?t~�9��˫��v(��J�gp)0��ٔ{,��~H��o寋.o��^�o@"�����p6��v|�.+I�n�w�jn ت�_��󻰷�u_T
oX#�U�-�R�Q�-VX�)�V�g��xYGxN}�o�����$�?���y� (�f<�0�0�~g7l�Q�2�D{���8<@�P�:]/�a&g}�I+/7��Jy�us7ǣΧL�j��~޼��A��dzҩ�OK�F�HYٽ|�9��Fr!1���m#�W���C�i�5ByY��L3}���}���+c��ǲ��l��
{���/�X�WS���&<��2�Ԏ�|C(���SP#��s1�J���_p��O�׶�l]��g������%G<xE��΂�m�'5k�/,�����NSx��B�͞)�=���5� #sƪɓD���\�
{��l�ոBӂ}(�M�St/�7$V���	����hK�͡�Ac��hM��3���:C�%�@���%O���O.Z@]�/��=�}LZ�Q�n�ٯˑ���V�t���[���9�g�̀5���.)���Q���6�ޫ��`�P����!�9i/+N�~�HX�ٍ��>�¨9��[z �R�]���4O)� I�a�,��o &B���H���ϓ��{��g*�����W䑁b���8/���� bӛ3~
�i�,	`|�s$�2�<��`r.�'u�8��Xw��|	#��lOG�fV��/�Ѡ�� L~I��%ԾOy�!�
S���*i65u�c�l���}��J�LmO.��������)����$g5Kd��$7������""��������i�#�7��?���e|�ʌ�V��@�,��uEU�$�qHo�;��������z�`f7�����@���-�M�a@%�ތ}	��j�CC��7Ov�h��l�l�r���n����LS��(Ω��I9Mѥ02��r}J�[�϶��"�ʍ�d.�D�Ɉ��;�b�������^���]WU=C�EL/��g�w�]yi�:,w�������ژ�`<�����>BN��TL���ʏ�9�%!#q�:�z�py+���4��|�u�/�]�$"\�����.��4S�߾k� Θ�^��p+�r������X�t�5*Ư�r�gDx{P���:l7��%���[���2��6{�Z�3.g.�%VQ{�>��[���s\ж�0A�E��{�vj��i����s��\����/�?���d�o���ߎ3	S�-%���j;%,݇�Ps�O�6Q�l/���>��[�D�ڮ��������;��z���˵�����:Nč�h_�Ќ���#t��$�^��4�s�y��w��]��@9���8�ȜW�[�0U�˝GH��f�|b�}��=V��� �t
�G2]�F�%�#ĈV�yd��E�Q��T�a�E:��J�|���f����N.y��8�J���Q6<?�U�C�>�,"��^KX�m��f4��_��*�N�s��˹J*z�6�D1>d�AzƆ�$��oB}CcNtv)�?(�W��3(�_i�NZ�'��Y�� m��ۉ>��e_b�dh�MLܜ(��n'9y�'qǈ� )@�΄��J�.��`a�q���f	��Z �$}�nxC�yБ<O�.i�N�O��fT*y>:��[�x�.��3x������i�������M�Y�=S;)�	��Sǥ��H]�߸�PR+�êll��������[,��jwrSI���^����B��,���rE������K~`_�=�>g4t0��i��M�~'.T6 ))P��]�Ĵ>���\"��ЉX��.ic'\s�32���>i�� �If?����T���_����0���^����� *�~��[N>�<�Ih���p��I��i�f�6ŋ��;J�$*�O���k�@>%���O��<�q��p��-i����+�CQ����ᙈ�!�����<��-G�F��]���=��{׸�2~�-�vs��;���A'|amLmD�
(����"P�}���dx=h���Ȩ�ԯ�xq%���ή�о�N&]�rC����JM;���-��B�	J>2�!">�˛)�M]��iD;2�krt��޵�.No���a_欄nk������6�Ȃߚ-�^��W �a3���*xR��0���ڬ�����@���&�d�&Ո�p|�׊zc�1�VB�0�S���Y8��k�[��=��'���W ��\�!�'�՗I�,ZW�87���;��8�/%�f�>���N7�)"���|[�����FvJ��̩�s��t�\M"a� F��-�+t�~�:����ǨY|�Ⱦ����p����^��Bh���b�ӕwT��d��}Wo�n���aJ4Yds��u��pv�o�;6�c|�o=�|W_�{k��^��X�C_��8�5��ߝs�w~3Dߣ�I�K%U����k�������d�H单Oc�l&b����_Gn���W~�ƪJǧ��p��φ�v��'P��R㊧�E���q}Z�O��oj)��Ie/tO���X:3
�]��D�MZ�b��i���>E�v�4y5YX���<��}{Y�� ~��
�ӯ�N����[��#xݨ�O��f	͓�7]�	Z�0��>�� �Jr�^�\��٘�c1Q'j��=	�����=&����Ϣl�.��'n���q�s�bf(�,��ud�����/>e�%ŗq���s����{�wϠ��Q�z<�6��1�>KW�q׌D(�X?�ht'sGHz_jK��5v �JQN��P彰�,�OҰ�TQ���$����z�tr���jR�B��TY���&]�A�Tj�g� � +&.�.E���<��?�8��3SΑ�l#	\V�g���-��-���!nO�f��	�W��n%����vĽ�}�G@;�V�}v�d�]�Iֺ��6�G��Y�눕��;ܾ�	��6�XV�����ԭtY��ݷ�ӷ�o[�U_�pFK,�w�7���,.��c��-�rK��;����f�Y�K��B���	̓8��{Gg�@�. v״�?�����������t�W��R� �������C��#�XZ4@ԥH"���>��䤹��:QP8�����}\���5f盒7�BF����;��і��V΂s�#�í��tf�ι�ocu������,�zkH������l�$z�q�~C�/�a��̝�i!�Q����Y+[��7��<V�P����!��؇�m���X-��I�)���I�"ƺ$9�F4,���xhX@��q�l�~�;��K��N�� �bP�
ѳ�up�%Ҳ��Z�͗�X���!�P=� �O��Ƞ��>�U۸���ѡ��l>ϑIX�e��bج$��#�<���c��$��n�M)� 8��5��0Ψ�*E*�N�DQ��.>��tzO�G?!?���	�V�;xk`}:��S`u�p���β�*�R���O��i��
�ycTs|Q04�V�yT���	���3h-A �(��.<�+�f��Y���b57N��h�G��kNX�hxJ�\E"jHZaP���k/#)��*$��#�>����D������qq�t$�S�8�}4h?�\�< 2ڂ�se�(�����U{u����LsLn�@�<YJ|`�B=�Yq2z��y�h�`R�C"�/���|���q�
�[3�1�˧�����E� 	�l3���{,*p�DP��u��h�Aws��49+,�D�_o�~M��=�PX֫�	��4;݉�ޥZN5zڞ93�̯*�fВTI�|��I{!R���$�m�R(�~�I]~�(;�-$���'UK7�$��V�0�xe'���ծ��h��H��_*~9$����6Staz�h3���8|�?�Z\"�~t:�#�%�L�~pGZ jؼ�Ι"9��w����R��P8�W#i4��c8&���@�a����u3C�/��D��2Lm̜�΃�,�Jk�#܋�z�&�ȼ6��H҅U���vV�SQD���O��ψM�]U2`�H���p�?ɾ�v�s:C��'1v�.(�q�42��
X��t~U/}�3�9�sB���VƉ�߾a��xE�|��L�g|�)V�����>��R�E�����7F�ZA�8� �V�w�{��MG~��J��F�5������2VG7#�Ѓ�q��I�Kۗ7�+�Df1��Y)Қ��Ph�$��	Ԫ�kB����2��� ep|'l����n��l�B��Oo��h�6qM��[���yI�pv�v{�gk��Gl�K@�Qy3��O�4��9pG�|�c5����Pu���iP��_��ٓ�,��թ��U:�R�������$G3{�b�k.��x{~�P:7\:n���?Ž�(�d�m
��綟�Mi.+�E��?�gb�G���/��*KI话òZ���#���,��%ބM�Smڊ�3�^�9
���v��R飹����=2��Ŗvs'�(��I��gF������g~d��%�a*p�Ӑ�^�;�bh��%��L��$�4骄�+�|����[�*9�v�>�y��dJg�)��堑�t/�(14��a7M\� zԲ%j��8��4p�0���ͼu^=>�i�4��c���[~�)m�q���KF/־��U[�g���c��b�B�@p��$� �وw��:�V�1 �b/��oM��h>���vp����NS��И�#"Pm�S��^�	
�",�g��2x�p�A%<��s�/e�O��yW�Hw�/��w�?OoA���u���|��=��[ �o��.~	�����x%[O�c���*B�ښ$�MW�ı�5��X7��1����Hl��ݤm{����
;�kf1��s2��&�#�������-N�+s�����37�����O�5m
q��ڨ=SL�*I�I�jp�k(�K�1vA~�$�3�]��������Lb{��eF�����)�y�����G�� n�w��j)Et���= �r�ƛ���/na~p�L5���.����8���~�5��75�?�y�4�x4�������u���T��n��y�7v�̴^�B�Ғ�BDJ-��~m�cL/�˕U.�y����mب.Y*�r�/.<�����G�fM;��p;��
���ƥMX���Hbo��4K�͍�j�q(��)�Ia���E�*��6
�%��\����IC%���6;i��W������w���r2�|��->�n(pα]��+|$�KB�*.��HcߵJ[��ޡ��jw���*���'gk�K?�8��#h��ߪ?��9c��P�$��bL��fw@H�b�{�gi&���<�k��YD���Ž$Q�g�d2���$P1��,IIgW���ܴ.�5��;aq��ݶ����	9��@O*L��ΏD���L�t	LJ���n�ȯ!��%xCQ���Ѭ�.]�β�#+^h����d}M]�� ?R�ĆQ�t0�~��b�a3u�r�U�e	Z������e�]zX��n����b=i9�^�ްe��L�E�I���tяʬ�!&ю<�
&Eqo���?�| c�(�îA�o��7�^>���b)�i ��<�X�I8_~�[�.�J���|��ʠɜ6<��|>�Y���7V�+��َ|T�iV�=z�S�F�����j�T�崛��b+7��~z�F}ىwº$O ,�By��3sj�#V�no/��2��j@�o��fM�S�
�gy^����[�TD�/v�!=���
$أ[�\�H��~uhm>0�N���sj7W��0aH1�	a� 7=4-�;������r^>�����ghx6��Y��k��`A���<R��J=�A}��r�ѳ���!�%�ˏ9�9^�:
���	Na,�Z���J߃^��h_vU���#
}��u�.� b��m�>���4/ v\�d���@ +�%��4B���CK�e>?�����zV֤arQ�����}8����X��،�*��_��)���m���,b� �ȟ�9b^��'cu��E>(�?�ӓ���P1��4�,��yG�շB���y,Hj`��)'�֪��l���Z�e����<��	�ޤ[��a-ӊ&ߵ�w.�$�b�j�Us��Z����@�o��R�����ҵJ>vx��/H9������_̇�5��4i]���u	 =r3���O!Гv�zs���H��~a�r�H�ָ����_hU�bF�Q��f9��,i��,Vi1s��g/B�|��_�6�q�wk�'9�xy�g�\��q�bMq2NuO�ɩ�q��Q���`eT,l@�R���u3-��6<ٓ �\��T\�#����m�RU�RiըZU�v[�vmJ�-Fm"�^EQ�.�{o�7�C{�H�������~�{��=�9�s����}�[y/�����M�%���'���t��'�k-��	��Ա=a7��k�kT}�ۛ~��8�Ƭ�����2v���z�k��eMf��To�f�[m3>,k�c��x��&}��-�0q1ٍVk����Iqo"�CÆ��κET���F��;?���:5(a���������~[6h/��!�Tx���#"Jbt� 3TG|�����0|/�0�SRw<i�<�5�L�uTC��_� �L�̔A����y^%\㝙��ݻ[������Q��������յ�;dSs#�k�J%��q�:\���)·J
���W�AE��|��g�w�4M?�Nm�L�찥��T�9��\���Br��w��/@9���uQq�xV q�Ǽ3ܗK�� ���$�et5�vM#����]�
��oT �4�@6ng���l4c��*z(���W���/+�k��gؓ�]~!��1���'z��8��I�\)xEo��6�w@Q����ގ�}/���)!���8��dP
��H}��~�l�����N#�jT����P���hU��0����V��B���{���aB6t�;���#�D���u�]e@���]�(f[pq�^���4=����&@X\mj����u���S%�*{��{o�Bָ`Gna�ȴw%�ؑ�P��G�6'�mZ5~U!����h�6BdǢKzP��տ�XK 8�{�~�5�����OP�r�������wYq��	�N��k�����zJ�9H7
 qaWZ{|vXs�#tď�F�h��B���֓��A=�����P���]������Y�V����K�M3	��)��Ry�)���J.:���2~Xb!�wk
kE��~�c��_.%QƊ��I1@m�TG-��j�nR`����o3KA�K=}?�z�E�|�Pua��!|%o6Q�U��tUi�G��a�:��I�Gɣ��yU�'?�e�*(��+�f���]��܆'����͓�z�y7��
�,�%z��Isr�Kq�s��(Բ��f�N�����ҷ������I�5g�Q�{]��Y����e��ғp�V�P������ѧjlxe��&����:����"ę��ffODF*|Y�X��`��d"�z|�}�=Ƈ���c lv��՝��G���z9�/|�����4r�w���f�
�L���f6�lLA�X�ڤ1��3R�aٻ�d�ڍ��.�{������C��n�&5ayY/o��� !B�{22��g3D�"���s�Xc�}�$>�@��� ��s{t�������A���&��c"aD�Ҵ�(�HʌM�C����]V���4��w�����Fu����}�؆k��l;>��T�,�S�e�bպ}"08���K��38�{S SB�/_��֬�����E�W�h�#�� �������Y����˴�֊�:�o�w|�5O+��*��~��JU�=<��#��*����)=޹: 8��ý}�4.�q�s왮�?��!��jy�G�"*U��-3�9�Cz��3d��
Z65v��"d򳰫T�͟��	�<���=l#N>�Kz��,�>'1�'���I��aU���g�%"�o�#Q:�#�"5��#�=嘼�9z��qNd��Di������_D�]UCw TS(X]N=E�>.Z}����+��֗��p���a �Z�5��q�t�b��CM1����q&�=�^9�dD�쟂m�|1C�Ǯ�J�a��e-ǫ-�̞������'|9��s�ΰ2�F2������P���mS1;�N��ȕ<���!VU��c�������[~��I����_q��Q[�8�@:#h�:G����������|��C����^C2��iV��<qW�MP��I�붸»M�L�9�ބ��f���]���>�(��e�S�6�d���z��-��c��B�"-�n�3z)�֗Sg���;�d�[�/>'~8{4&@�[��>�[�ҽ�q�pt��I'�N�'�pV��-͚�VT&4F_8*ݱ�à�'KODh��s�70~����j���/Iј6�����g%�&���0�fi��7A<���jZ����<���W��ȭ2�L8S������A�%b�g�'qTH�]V�i&h϶S���/|T(m�����>���ϵ�C4*N٤����u[�y_G�[���l��߻P}�ԅ)Bꌱ�U)z2 ���*V/�f6�����_�&h"�+<�!�Tԏ�j9�3zf���el֜���E�[��ǪՋ��2��t��ج��+W)4��$����<��z�ؚk��rX� �bOO�+'��鏻�O9B�P_rB���Q�-��[L��K�K�����k��4`M���2��嘢aMo�q h��c�l�D������lO�طQ��	z^�xR�ݚ|C��(X!a[��������(
M�(.��.a�Ǆ��Z��5��_!siq��@�x?&��;ɉ�p���L�R�{-�q���|oA��KǤ��Z4\��=Jq���~�G-:�f���G���@얱���q� {��K,^�s��?m��ө��r���X��4�J`�-+^�PT��;������M��O�}�}���!�Ƒb�;���K)���p5�y���3�7���p5��f�K�dKM��k�Z��H�^�rL�շi�v��Z.�bq�w��&GGz[���&O4m�WURyB?�UYi�R�(��m��������x+l�Y��5$ ����ûX.7�������Gtew���&�-#�=�<��#�H�cL���S?����(J�)��j�z翆s��Z��5��)ɧ�n͟��&�Sr�cy�*UW���*�L��p�����e�5��"8�{��I�ޝ9��<�N{��e���S'�}���|�W���^�0�*)ʨZ�̉%ؾ�U�c�{$�xU�BX�z�1��޾t��=+��E=��"���?t�L�8|���=�~�3��i�����L|<sO)��_4��,z�cQ7%?�W�#ł@m�v*(�� J�u�_B��n�E��a;�w�H�:�&	[T�T���z6<J}�8������BSG��<Oi��E�:b��T�z��{�r�@ˡE%\W1{d�9�@���(A>6_�ӆS�������Pg(yi�Oʡ�2S�v�DT^`�%j�ۢ�h�Qg�U�W=_�>��۞�z��6|c4�HZbY|�t88K���.�nEⱗ꺲b�Tͧ������(,�3��Ju��푲�vկ���i����w���	g�d'�����`#2�����m�u�K� �������p9�q<4���Ra��) ����O|�2�ձp����J���ns�*���<�7f=y��e�܈�h���g\4�H�e�--�6`�����ᨴ���ٞ?�Z�V�V\L���QTM_D�M�0����@����H��kigIh�A���!vP����ME��fYb��'`�˟"��ֵЖ���:��rً�ߴ6�V�>40�����]RZ�p�a��;�jZD��t���ӲO۶����vjޤ?���L�-$�H��Iĸd�NJ������Owf��C���f
^�'v��_�+���b�^��p<b����1�{Ty��������'�΢$Q�����E=Z;��]�g�v���/?@�#��w��J�.`U���� ��o~��j՝�kx��*í�fw	�>��x���y��ꤥ��)'V��hy�sHe{/�rb����/�R�4_�K��ՅZ�]0}eH��ep�9JBזϫ�=t�P�r����b�B��v����1�7ǏQ>��J�,S�C0�K?�4b���s��K('�"Q�X抌p�jO�8�#�/a�ގ���&d��Q;���R{K��(�$;q&���$�57�Z�'N}ܳ"0�ּ����E�i���܀�ͼKҶT��|�P?9d�'��ER�EDm��N�;c��O}�No�m')���ި�{��魥�l�YiA������36����wN1��0��P��iv�A�\lf�Ǟ�[�J���ؔ/G�.����'���Ӊ�S�2S��uG���?�6�u�Fmy�	����a�� Gd��q)�ձE
c�"�_/���m\߇��������o?'�܄y� ���s�pi�z��,�u���&�	G�<��k�=�ۤf��])c>���u��/q�/��f�
��<����@��/��q� o1r	gD|�d��X����dm��~Q��&Yu��DZ�t{���ֻ2�8P��V�XW$���\�w��cG@���n�^ր��tC��ܕ���E�^#'�w�Ty�n�g;�h�9�0�2S��8Ʈ�Dv҉r}�\�D��-�6s�_Dv<￷��C*~#�� ��4��x�<ظ�[w�J���Y�� �V�9����I�b�X3�K;s�K]Pp})~K?^w"�����~cA�S���t�0+�,X�sd��-8Gm�v�/� ��-	\���%�g�̤+�6Ʒ+ w7���D(v�1t?���1a�[��Q"F����"��-2c&�̻V�߿�>3�a}-ЛBm���ۭ���"��!g�]�E��f��d�eYMo��H��E����E����9�YU����P1�Xׯ�s2����K�
���{h�J)k���t��>�P��X��G�<'83;<��u��y/��<�$|��	��K����MV.���q���j��k~�>��C�]#T��~֎%hkR����$��s�p_&K��PW 5��"a���i���F��b?^����?0�,e����Dq�J��he���ʾH�
.��])EE�mA�S|e��e�T&V�[G��)�~���@Sו.S�ٲ��>b�Al4�7��+���e��L�n��NO�ڭ�G��Sa�$sL=xfi�C��o������0~��i��9:0�ծ�t?�9:�z�z�����=��HF�0�9{��y���x������w��iH�3o�C��w��K(���[��|ۄL��M��w a����ЂR�j�F��^��k����Iť�L���e�&�Vf�uI܁-��_ƞ��N���qKĊ�#^�_fM>����y�c�©ڧ�?	�Q�HFn��x� jF���wA,~����l�Y+ݴ��%4�B���TY�w�RH��_�I�ʚ]q�4bP�A�P�QL�z�w�! ��V����3י�����߉����uWhN�c��\PZ��^�;g���\Qd��Β��
���-H�eYJD���vwQ��t����Q�.6���O��q�[�mC��r}�r���kd,�f��\Ѽ�Wひ��f�|��6��8~^����R_7�!���ґ-=���p>��uA�����Q�7�T���;Ӭh��#aQ�r k:�E�r���\!����F�-�ܞ5���:��I���m+̈N�*��'���>/?�L!)��r�Iˡ5�a��8�=4<gP�tʮMܝ��+q#��7�T�d �(M�z:�4�����H�*c4f����t��
�Nݟ�#I8ˡ"s9ۀPyE`�Le�d{=���ʁ5ړ:�w��\���>.�0fq�Z8�BFm����#����92j�d�����IL�B ݁�����߻�� L��U��#��l�Ǿ �1��]��̧��)���'.��{�O�]?p��;�}<u7I�+w��8m��.U����}�{TG���ϻ��J�*�9�,�t�qy�ZxN,%���9�҄¤���>G�����%=g3\��pyT�@��B�lyZ���'U����D��w)7Z����������VRė�{@��k�����f��O8�
 exM���RSR�i�۸�1!���^�)���?I�w��o�JM��*��/�]�/����(��RѦ����Jz<��`u��X ��&O�h`6GT���.�d��ޱ�3��Ui�K����V��Ӈy b���ŤV*�FH�Y�q�sP�j�co�ؼ��l���?��\z�&KiP��M�j�b�)vyO9�Ͼ�̑��ɖ3?���
_����ңBO����ߺRm*� �>HQk�-���tEg)_�M��8��!k�=��2�@�l$J�z�vھ�P�=t\AD<	c=zb�?��~Dtbd�)�3�L�O�9y>}���-g*��ï8ӂj@d�H�A�ص }_��x�FoU�����ͅӫhp�Ur�g���N�2���%tTS�LitAj�<v<"e]ms��M�������TFH�#Y��;R�����>xP@�Y��c�;��0N�zdm�ڶR���s-��כ��y�8��%�,�ڕ���r�u/��T�wJ%U�_�B��+0�p�!9|���繀䟴��bvg ͑<�5'�"��?Ns���y!���:�]%�ty�$\�����>��; �Ψ�3�u��s�O&�#&����-�`��os�R���ߒfukS�#n��5E�X��-�^i�/�T͢�����=�E�Y��t]���Ol�Or@��=���k~1E(�/��ׯ�F#7^f'��B�^��� �_${bt�8�i���5�����U��xtJ�1[����A�DNG���f,s+����z���|�MtN��d�E%�E�ʙ���
lcX[�Sir��\�@��΄v]���J��Z�.Uf�]���(�\�X�vL��QrY������{�<�@w��tʔķ���O2��"�Z��&�7Ѭ�l1��F��S�ib�8�	���,��ȧ�)m�d:�)��ֿю���mr�ԪJ�5D�����hA���;�p���(�*J�?O
[�>��)pAˑ5-!dУ�ԛ�E2�|'�f��PD^cqNC���YX`�g�����<K^� Ak�iOߧ�v��*9Ĥ1Nl��lmb΋3%�C��1kzV�F�ӎ�^��ؙ��@�3�����}�6�4ԋD��c�Dce�Y�Q�@�G��R�{�/�t	�5�5[d���߼�^)�q �TX�kŀ�w;�[���7ʯs�,⃶�e�N�v#�pe��	��P�� 3�@{MQ���N��ƌNuo����fP�9�"/꣑���~f�Nr뽉\K�Z�{%���f�b
=2>�V�|b)��q�;��9����?��"Z<�D����[�h�~��J���ݍD��Au��]�2AÃZ�B�o�7��������c���n{9�l3��937�j��.[�N�_�U��v�?Y.˖>�Q����+��|k�����V��bO����>Qқ;�I|�S�@cS��tq������AS<v]N-�E��+�5��q�<���nq�sDk�4Jg�ц��f^�Y�����`��#|K�K�Yj���\�?5�M����q��+;Y~{�۔��$h���� >����E�9�eK�QI�Y7�.���H�ܓ���}�@��Il��e���hH���2�98-vƴߟ�mc��,��}˥r�O�4���o>��I�э2A�鈅ң�
< �G����k�_�q,������ې�[��7ۯ��u]�~���.A�s_GKW�:�W&їƄ��OZܺ.�Wv�X�~���uߍ�H�����/�Ե$��yI�{���@�����|�5��h�"K��K�E�5���z�����i;�Ӕ���#�q�{G��Y����HR�1�-�
3Q1�kB͏��Ț�2���Ws	��G�o�"R���k��1|��j�P!&��:�l�b�)�����^���［��-�gQ�dx�h���ې�����fb�c6:�.ܵ���,�T��.�y�2��!��A���GC�m����R�l��a��<TS�G
�Ym��[��A������["I�~�i׊!E�|�Ğy���U�.��K�۱�p�I�Z��ol�:�4�+7�r$|E6�����o�*�y�!��'����6������o>�I%[_���rׅ��7�q1|v20g����)���ŷ����D��>b�T[�1ϑ�����m�˸_J��b��9k�n	�&0����g�����J�Y�#����ڃ��;�\�Ol��^�a�*� w-3fi�^�4@�5����:�?�"}����+��h�[�Ը��)�(8�VH�cI�8�εѹ߯M��R��)q�v@,yn��|�@��5�h?g2��8?�}��T��2�tU���n�C��Д�!N�4����y�冥k1@�F�;5�٤ZzfG��wJ��o�Ҵ��
���z�gw�U
��Ql�/�5��[jՎ��(L������ޙ����7����ˠ�v��wA�	����fZI�]]O�M� ��v�ڣ[��"���� ���yJ�����NV�X?��?0<F�@�ko�z[z��|p������=Լ�Ϥ'�N�o���7Bc�:��?N1[�{e��k�t���/�Q9�q���Yg����2̰�$��l��pt����ُ��j��+k��e�z�ϗ'����¤GYj|�x~!fl�#��_�j7=�����O|�.'.|}"jZg	�X�O��%�F*YM��@�"���z:e�<x��!�����OZ�<|�����J\���'�jnnP���(��� ������3�sƹ
p�R6UI̹���+?�\�6�B0�v4���d�䪇���͜��%��z�^����4��`��@���ܩ���1���F�\Ub��D�&�Γ��׏�'�O;��f�'�cn��[�����I9����߉L��P9̩�]W"|��1|�Rt��׷��r���[����k�]�����9��wT��_�Hn�w�XW0(l:^�k"#ׯ^��:������G�b�YZWY�j_Y���$��բl���QV+�T �q��;$/_������;n�
�#�_�Q�dW�.��z�Ɛ�Y�H����<��$��-Ƙ�"�K�Q���B���d��/y��04���ؒ��ez��0������xG<��4�F���hՅ'�[uAb��Y�]n����=�]��s����'ډ�0@�'�		;o��<�v��}ql�ߟL�?�8��yOsE/����wVW�/�Ƣ���
�re����y>Y'S��Gz���x��|�$5z��+Ћa,��-sqھ<^���T�aQ�NlNR��?��p�M�����i���4�JU%C��x2�����}��C�׾`�����D3�3l{� "��Ѻ�Ȣ�U��q�o�Gy�F��'.��'�+
)�D�A���ɧ�׬��b��t�jD�v�	U�*�,��ïyM�B,8��F������ ~���	=бO#�2O1�)�����/�:�6���kà{9ZB�~I1j�<�ȕS����̻[w�U�:!ɬ9����Q9_R;�)rR(`-���0�o�R҅\��P�փc�QQ[ʤ��m�E���w��b~�.`�a�d�Tj[qZ�ڧΒ�>�w&j����L��M�d#K��X̍�M\�{�V½oYSL���5�|j��.JW��ݠ�A�F�^f`�?�1Պ�M�]��X-]t�#���9V3ȋB�@'u�i�]�j����'#S��`�Y��ɩq>t���hn����;��g�W��6>P�ͫ�\�� Da�L��d�

LE��MM'��px��:�ŎP�R�VB�}|f�qk�U#U�K"�O�W�{n��I�>�}�Wmay�/� 
�ଝY�(��y�L�.�R�'���_#�.}�Ѓ¢�]�x�����0d^y�4��������\�����AM�/�ԛ���}�m��X�Y���i�T+���EL����Ҝ|��9g%�n����xh��ݓ�t��}�{��%��67����k��嵋z6x���\���˱��r�{Ue�7�L����*��xZ�>dͻ�ޖ3��P.q��Uԗ�X.�F'%g�8��|VB�ؑ,x���b�k��.��}����3�^�d��Q�b� �.� �EOW��zZ[�����JG�8j&6�5�L�C�iU��k�j�Bo#p�m~K�����!�/�ʑ��a����;�MK�`g�Gi�qX�$���oV�����}�_�>�1�3m~���Q�Q���p�7/�����L�Y�.�.E�B��W	g�W^���o8��2������$�.ȭY�˜W�^Jޠ���K#Sr�$ݵ�vuvd�F��hߕޔ>кnt��p��q����= HKZƟ�v��I���>�f��Ag�-��R:�Fų��&_B?Y��@�O�}'22F��kB�b����<SmT���K��bi��5l����/�W-��ɒ,r�p�'��934%�S��#-�<�Pbg��vLo~�l}���K�M|���Y5�Wg����[ 'ªoD����^�k�!��`Ա�uY��!�S�a�E A����/��ބ�\���C���ѕ�ZU�륻��uU�Ni.��e���گ[mu��gߑk��r�	��Do�dF�5���/Δ}$�T�T*��!}&�q���?;a����)~�k�8���aX�v'��C���6:	1|�˺��~��8�vV9%��I��.��L&�h<��^sĆ9��],�D鿠ڣ��z�xf��� ��;,3s��`V�D��G4/6��n��>cD�s��?u��:I5AR=��_�Kz-Q����B�>H6/,�~ȴ��Bn�/7R�k�K��N_�Y.���φ�"�<eeN���	܀9�:�n��
F�̫�������q���n���i����}�lc����j.�M(x����tP�;}e�e��e�=a@� �q]v�u������.a�i�"��_96�HQ�!�c0�=������˾0��$pMa��[���������?ƄW�~Y�w�=�uߧz1�-q�k����e}����R�Z��-�n�EH����t<i�y���5s�lӑ0H�� �+ ��}��WBDj�'f�˩���0���W�0��f��¸H����%1�_,�'�|?�B4�x3pK��!E��kn�s#��?"����z ��6�l�mX�E�����z�E��>F�����ho,޾���K~���Cs��bff��+��abwZ�����v�����(4ʼ�59t�����Mّ���j������Ldh~wV�P>�|��zJ�F��X�`LX4�������c� �}��8�������0'��+�Ed����I��Qb_��]�D^j>
���f������d����w��M��)b�)2<j�_m>0��h��bZ�^�'�(�lۺ`� (�5�K���d�7IQ�(�ʖַp�Y��)T��e���_�^�3�j�Хuҕ����ݞ֜Y-�Y�qk��k&����LK���o񠘫^U�����Xi4�f<U�ɢJ��=�]Ў���wȪ:C�ߝfy�BY��/T(1L��Gw�#�s��V�Ì���N�kId����_�������s֓���9[x��U�S�?��P�G���0ٕ ����C�$$o��@Yz><U�qa(�gq�	a�J�yg���/X�ś�F���	N1
���D�P��N1���>⡐��[Ϟ6?|��q-��A��c$������sԸy�)�6Xt��s�O�P��kAf����p�� Ѕ1�=����ܱE��MD����O�T�>�M7Js]�Zf�t:����*s�"�s+�]$��+ᛃ�׾�
K4}�����
?������e=�7����\�\fhP��E^k�~��ɋ����U���:��!��T7��ioO+M+�L��K�*s��^�bF\���I�y��TF_l.��V1f�����e97�O�	�m�[��q^01�V�ڴ/�ɴ5_��M����r�3��iU��F���V��Y�`B�S~�z,���p�&�[��و_�70�I���' �gvi���w�O�5�=�>���u;�Z�䷻ц�U�WY��ؗO*����M�>}��e�9�����x�+���
a�d*��G��ƌW��L���O�F��X�
�R������]�>j�Ew�������.�*i	a%��bq��;�0TᩋS(놀)=���iSx�J��v)�4�K���f�<p6-w,u�Eq{V���5D�O�r�k�x��%Z����Ù��ž=��v<o���M��©C��{�#{�b���`/�⍰/��Y� �YIo`(*�K���`��;)~$ϥ,�2��vذf��L[s�ǹ��Q��ڀ�\������>��3����p����?���B�H�F��)�M��7 �rwD}'n} 6�����o��fx!┕�E�n��mj_�*�W<Z�\-����D|�¡��e�j���\�.��>�Ȇ���%���ev�LL<W���b�1|�}�zux�,���c!ۤ����(MͲ�Db�W�OZ?@y�����y����35�նx6A���l��SO3�V�+��!2�a��_C�U@d,'Qy}�l^z~�	�ݫ�`�ѳ *5��eL"[=�����5I��C<I-�ħc�Y��z��SY<��[��!�;��[�?�K�ў���k����ص(ܠ&^��a�D�}�.�)xs&Ct칅ʄl���"֙�'�Ѿ�FJعdAz�Z���V�����<G�Ή2!���0�ｲ����&/Bƾ�\�b�/����6�dC�����_���lk7���>�m�ak�G{tJ��Fwn_s�bܼ.�`b�S�;���q~2���G.2a9>�&�x#����&ƣ�Sȁl4��z2�_麏j	⯎WCI�9�._��I��r =L��En�f�p,;��H	h�����>�zBP���K0PK'��P�Ưt�����^&��h
�S3����S[�Rj/�]��8��F؏7�p�r�����4�IV�Gޅ^������v�r�^��|g~���������NS�G{#��О��)�h���y�v�C��ê:��}��[h�5���G��y�=`�x�J�pv�ژp�N�s�`>S.�l���\�n�nS���Z�Utza2&�7W�}^<g�|����XL��*�-�}9��ȀhX`��y,}d��;����/��]3g�������'S�y�g������>�<u!|�������<����
���qБ�@e$�/n�B.w��~А��u^^^�w}j�[b!����$E�޶�sO�f墩o;n�]��l9��K�J�k)7��B)��� ]�EUӦ����5���>(,�EO8x(,Y�,z]5�x����e{�0�|j��>�'�T��(9缨�R�����~��/��f��Ҽ�Mg-Me�S�l��k�;p#@m�����ZR�R8!�n������>���}x�>�R�1�c+�^�Q�=3q�{���C�H��kR��g�� tK@�L���f����:V+�4��U������D�m��r	k�3��W	���ʎm��-�B���ʴ��|x�|�-�e��7ϑ�.�#.~j7xmo���k�Iw���Е⚇ ����yyƹ��ڭ*O�}Y/J��l��gI�.���/�"���q��i"�Үsg���q�N���V!�f6Ưm&��؉^$�օ7�MRf��$$�@���m���M�O-��Q���r�y��)]F�ׅe���,���
mF�#�7������T_7����I�Vq���Y�fUQ���$3z�!��[]EJ����0&�a�`4�El�*פF�iϚp��1�|V.��,�Z�~��⛴C������P�7��G�������ϣ�u�Ā�F+%)�Z[N~���>DOG`�OƜr�0j��ߓ��'�LNg�����K�g�={�73���� )��[���5>'1��="�> a������_^����D�a��I�BXQ�	U]�P%�Nm祤���$0�Q� �t�%�a�Bz��N4�����ܿ�tK�T^� ��q��Y{��>���g���l�[B؄pvK��7�����o~��E�Y��K�>�6ƣ�|@������O8�H��2��ѽ�:�&�W` ~��O@R�WP��W�o
/�-��`������������vƍ��4��cӻ�'���:�;�0W�g��~��ܾ�U����&���b��+�e�n����[�_���]�2B��W���uX-�uz(���!��I�Zlf����u_'�4�e�ٚ�6�b�%�������t׊c�
��1#� �P$�5�j
��L�e�U��7c�QiUOAj�w��3��x�\-/�f|{M,ǧy�*)�_"�܌��P�e���O�%��.ɶ.���<�T�4B���c#�Aމ����R�&B�p�n����W�_.v�_L��k���R�t�����<��8����(�u���捖��<׎�\y�9)������ʷ� B�Q3�����|�_��8>t�A </.�u���|&�5����*G7&��-��h��Za��J�\@v&��m��6�"F��weNH���Ρ~��4��e_�&���w�������}~�3��=#���ކ'o�z;�R�b'�~p�d�~�&���L�F�[��E�g��M;>��4ɴ�Tng�O��ܛC��n�i�[u١ ە��Px͆�H��k���6���^0��~�O3ӏ��|"Q/�t�� ���,V��%�y�,6�z2p^5���I���5�#O�4���������%g#$Ez�3[������f��m�7�nPj���=���jb��w��Tr�I�ݽ�P����,��ۨ,���C�E|���H��D��kF��[�EB�|�v"�Q�+�6*�-z|�?��O)��2��Yg��Cv�~?>&��Q>)�Խ��N�rӶ�7d>�j��H�f�y�T���ix�ZQ��>Uw������UW&(ǜ��(4��x��nqo�܀Oh�
�@0����Ne���?05)�pҞI^��;y�|t��<�N��Om�.���Dd�9�]���
�}�5�繱?�7&��bBP!AF�Q뻵�ܘ�B>�A"�m�)v�ͨ�-��:X�Z��=���H�QhVo�Ĳ�W/$9�LQA+���	��JeI�N��׏<1�8���l�˞H���#a+�s�i�EI_�/�a_wxl�^4zxz�!ܐx^@�ߥ�U����T*�%�:�{S%8U����	)s���e�������~�� 9������F����Є����jw�FP�)�,�O4�<q�z��.��#��������o����Q�=�P�7;PI��<��uqK˨���Ø&񜉄��с��� ͦb?\)k[o�U�1�y�OI�i6f�|����1����@�mLD�y@������f!ԭ9w	�,�}�B��j����=[���/:97
c��(\������ī�i����3#���୯�?�����]5ᡆ�WV�kP[$pdy"����N����v==Cր�]�٭QMpiL����ha���-�,ZzUE6����0K{N~�F�S\�"n����S���t�%�����A��,[L@Ԗ�ov�-�p"2�S��H�>7y��������QJ.�O��8�ꋇ��6�(�&���;���j��RP��zO2DFB_�w���8ɳa�X�Y�n*唤�c��.����S=�7����^�T��Do�k�����"�S�Ś>#h���Zק>���8�A4]EvWx���Hr0�>A��bᄫ���N���uo���a<��{�?�_(�L��T�;*]��I��/���J�M�JO6x��e���11<���"q�'�}4����ͻ�;�M���$q�8�6������Z��R�L��#�hኩ�GyZ%����w��3���_�w����Ǩ��_K��y+ �Ә���~��z��7�U��5 ���G�M���U�D_��~�Gak{Ä	&�Z:<��	A�R���'�?�I�7ij�(�|��)�D�6˸Dw,�ʹ�I��6߃܍�f�M�Ԯ_���}C���8],Z5r�^'�̒����$��	�e�-b1���������H1���υAc�l�BW	5��v��z��*�2�F/���ư��H[�����9t'�/�8���u��.1��Y\FH�;��Ct��g�l�D�ϴE��;y�<k#ˠU�������};ɰ)Pܷ+#3��8��zvQ��oT�$q3�{��Ω�C��g�(8�0f陌d-Xfj� H͸5�W˭���v\�}����a��O� l��6m@��O��/�"�6�_K��w���ơ�v�{[̕R��d�X��ݏ�$��VT�jS�Ϧ�Xɨ�+Kg��������,�>���lc��]�~�Dnf^�9g�@(e1t���-�{���#Y�����3��3vƧ�.���9�'��Z�:�M�H%��(�vJu���ʯ�,��_��]bU
��׍������uk�$z��c� ���S����g�4�;c��Gow(�	�j�@峺ؓ&�2Y���U���m��;����Zkc��Ԅ6F��Ww%����]:ݼEo�mJ���h�=�/�֨�ʻ�~w�㰞�ڣ����Bw ��C��Ǧ���y��	�z`��V��w���(u-�Boy���E�i�̓��s{�;�Ñw��Y����mh(uQ�������e�P޲��ğb�C�i[�]���K�2ӄ I���Q� ^� ,_���QU^����S��B�^���3��^M�ˎ��Ro���2�������d�����ZmU��բ5�Z���ڵkV�Z	� FUQ�R����N"�S�V+Hb�"����_�����r���{�s��s�+Dq�<�]��&=���ˤͻ+&O�u�fߎ��t��<~Z�l2J�<��Ws���_j/$!��G���ޏ�$;�z2�C)�>%�C��O6�Ylwwl�����E���z�N�1V�[E̞�iYi�]`�IИh��f�������/)��%�=뺨r��(�=��ؾm�_ڨc>@etz�y*<B�&A$�=�h;�P{G)�d]�����3\}Z�P�}4��)U �^��+G/{���c�[�6-���c����k�����霼���\FZE(�⏍�Y�QZ[�. �H�k<�W�͸�]IS�!"W�R��uq�����9:�P$�e~��|9)Ǐ4��\C�"6�vI�u��|���p=[���p	(CN����"�v�Q�T�T)�����|�#����F> ʙB
\���tfI����ޟ;�T~�z�)�������lݏeA �/�ڵ�Il��p�RP�[��N~n�U��=u|c�+��M���*��`+���%3�U��`���!��3и����'�%����<m�X��L��YZ�\ ���ʇ��5���9A�9���#���`�Ѹ=��E���@v�KЈO�H(i[j���=�8�3w�h��R�����t�H2����gh���GN�d�y>݀cD\��߬�������M~�Ï��	�e3�	MQ#� �I�2�<�(��1 �n�rUsW��^�4�/�rh�2�v�$"^I��,�Q���މ��؎]�I5���O��D��w�����9�$d�̎Ӱ�DX`>���u��XŖ�˲�
�]~�d� {�t�N������n�����v?�`���N{㟿2]��[�u����n�C�E8�NA�p��јO��kևujq�����w�H�b4ؾ2Ρ:8�n�p�۬2����A��ߪ����,���~���;�f]�{{��؅Q��ѠK_>۰����U^`����6z4����/�<��r�Ń���ScSk�G�Mv�ɣp���KW�~�_ȿHzx��,
�JH�A�@����5�S��$\�rUW�J��X����[%�e���p������".@��}0mh�q��'�WNo�el�r6�Ut)�l�|7�Q�Qy>U��:U�P;�����Y�_U)�$v��*���+��� �@�� b}"�Z�T6�?z�;0w�LS [��?U�f���X	�y������q%�"�_�����jQ��W	m�kk�P'�:��=��eg[������5��%���]~˽��QF0��[���gE+�?�΅9B��C��3|�J�-�J{r�=1�b/ǜF��K2'zl��g�[�����zU�������x��NX	���O�;Q����/��F�U����{|��j�X8�kq�P3��bq���RY�h��i�Y��;H�;�)�f��j�ɒ</��=�Ĳ%�j|��$<p�p�� �o?��T�~'�Þ2^��l��@�@f_����Lץx���l
Ʋ���7��+���1=��]<��TX��q��ĵ�7�߷/uc*�[27�8��{�;���S�B\
d_�_�\�<��=mXk�1=7FV��즒O���L�2��[y.p��=ގN�ܕͿP 7�M���
�Vlie�D�2�W,�V�m� ��TrBŦ��N���S�'ܲ/@�z{B����-��П�+�H;�c�eG�����bf�%T�����t~zwӰѢ���Nf��wㄗ��v����|V�x��[�a@CXIOT��~�K;���;��ˤ��4.r	�+:Z![}I�����']�&�}7�k}�I�3�K���B9����]����+v�
^�K���,�M�jR��/���
��/��4b�����D��Ѵ��~���?�K�$Ī����A�V=��cb�ۧ���\l!pd����L��48��~X�"�>��a%���n�+�c*x�r�>������*���߅>�c�8�6k93ih��V�e{r�^�W�Ґ�*m��[�?Mr�����i�K���K}</��1z�}��}뼬���];�u$����W K�ru3�������b�cs݊�)7kP��*�e� ����!d��0��M�����+�wD�B��E����R�:�a��n�a���<��)Fլ����!Ƕ�R�zL���ɀN�@w���d-��1Á�uM6\o�,Lվ ß;=�����I~��˻n���K>3��G%�z&w��߼���Op�nO>�8}%��+j��W���t�ZSo����+����"�#�o������_�Oʼ�T�����sv/�
��0�M:���v59;d�R` ,]����}�A0��V6t?g�H��.?
b�^!�z�t'�n�����xt1*�@�l���Բ�����Ti���ۣF�7��%����2ʿu�β#��.zgO|qw*�3	���pX��w�ع�|.��|�{�ԗ|�����]A�L!�
�7%j{(rTh>1t��[�)�t��C� �����g��U�1+hw~�:m�� isb�]��z����������9Vwn_i˯<����4��I�%D���`�&�������S�UgoR ����>�_#>vr/6���\x1�yh4�_��5հ�]��0.�#�����_׉�H���mۗ���6�	̇���&{@��Q�O$]��z�Uh�|�Kt����[֭�j�UO:�-���C�e�d����'��6n���Y9�������+T!�o���h�����)ִ�y��/ar�hT�tFf��'M����.n"Zu����������j�����1%��0n(�KE����[��ш:/���Z�5�Z��B����J	r;�~����V1wZ�?��!����!��3s��z�l^��YA���K|P��:O��j=��Տ,YF�ypr�(6�b;�z��Hw�5�.�|�'hR�Z0$!�ʣ�{�~����~M�N��2WY��ڸN�d�T�Y�GN�Z6���Nu�����ˎ�ɲ��W�T�p#���9=�ڤkH	�p���nu�WRr�QS���w��b��5��@=`�_�DFF��?s��=�4:���F�8�A!�e�߹���o*�
���\�h,�&��q��"&$��Ȩ&�jW����"�r�f"����ME����o�VT7M�6X.�ny5?��/��M��)E)��
���0��?V��}M�>�ۼ6b�v;�8I̙%���[�U�s4Ռ��7Ҕ��F��|�n�UF�]E ��]���鍥1��ӄ���(O�����鲵�����y�G�P�%�r���2�Sӧ��ɝ{ʾc�>(���� l&`�̥3&˗��#t����nH+���ef�"̣�؇%�c�ء�=Q����}i^���~��n�b�ڿ�>ק&�C��biP��ָc����a�ޞ�;&���Xp�I���^t�n��S
Jb(l<OE�^�_m�_&e��5p����Q��\��L���c��gָ��i7u'-�$��Ն�"/�W�6d��!Z�D"��Շ��?��4��f�>��,�f^ �H��T��������٨���w�M��e��x�I�<W��n�h���#�tMm�9�}�5�K3k��6����2c���q�*e/8���h��^�(�|C[V�)W<�����f%QK|�Q2(�^��d.k�ػ�MIf�:�Nn�;T1�O\*�����B���v��,Q[�@�}e�Ax�>�=�t��cV�x��R�D������=�W�������`=� �!�܍8�'�@l�D2�J:���Վ+���G�؞G���R�-�g�R�8�o'��V�Rt��Ͻ��Q�H�UޕCU�P �^�v�$-�;�:��&;��=|�D^�8� -F�����n9�W�(POd��udy��N���l�w�`���/p����̸P�\�8��a������2�W�8������{6�~��(� ��\�L_~ҡd�5|@*�	�*b����ԯޫv�۰�ꮗ������0N�p:HͤWI8�� ڥp�Y�Yn#��i0l�
�l��{�WN�l���.��/sl�{_V'}��3#�+%�NT� ���R���Ŕ�$��%h�V��&��@�4_|��~w3A�K�`0~:�;1�wd��d�9n�1Ujy����W�T����*�_���t���	���%ձ0�9����_��u�݇��ۧV�PW��&7���'���}���7�R�n��N�)���Qd��s�;��?��w0�ܳ9�k�*�QEX�����.X\�'�H��[��č�'�K>l["�z
�����L�E3�=�+:�"��
�N5�Jӣ�̤jS�X��z�fvjE��_t����9�m!�^�\����d���A !CmygO?���v��	����b_RY@�&@��mng5��^�ۺ� 	��=�#F^�̚!J"lo�yp�Қ^�� �n�9:/���췦#0��}�_C(l49�7z4�7k���SGG 7�Df�I)���A����M�����"�;S��S�O���Q֖л�l:�����PL
�}|��DUs?�����uy�OeD/��kOf�ˬ�r-����F�6ۘ1]&�z���e<��{Օ&������ܪ�[�+5K�}>�c*@�I\�Ito���<K����^��_p-.�~�"m�t���Ö�a�s5u��j�6R#�u� �5��:ӳFWA^��~slZ�{'%��x�D4�����4o�׏�7�ґ,�Yd�̥� �|?˪omؑ�x�+u>�%}`4�����6*�E=�~�F����r���r{>�O�ɸ��p�/S�M
ݰ��"�V�&���e�h�XH��$�CJp�3��@�	�ec����_���`�'�a��9�'��~ߩ �(���.w�W��+�\�
�a����N��mU�xד��U�`|�2���&�u	�G?,���Wԅ'4lz���4.��V!�������UA
נ���U�f�BzL�4����������=E��޳]R2�!T�mk(,�Y�y� ��4_�������u@D!�4�"~,T�x���@�a�R�<I �����kZQB=��LG�T@�dڼ��M����y�
�UNT~�@r��˥�W�z��嗣`HrK_~�!�<�UpZm�]���0�(�5_��dD0j��f��qeO�Wq�S�-cZ�������2S=J[H5I�wg�{����݇�t4��_��'��F�C����q���{��!��78.����QlJ��I���O�Q>7��3I-8��6�+\�0X�ީ� 7�����.�⥺�N����Թ��� ��F�g���S[xq��;��3]��`����8_��� ��Ȧ�
�kΡk�K^�|�TNQ#i��]f�7��hh��Y��;�>��X�sC��7�~��:����㡼wt�.w�G=6���δ����̶�'v|q<�������)4�)�1&sU>��V6��;��z�;���ut�`fSBF]+��ⴀ��>,ό�)�r|-q[��ӗ���
d�Z/��5X����*���1ZΠV��f��5�R�*�f�MS*�˱չضQ2��@~��=�[��nv��܆�b��n��<�/���9Gq0�+1�n�X��aAh,�ڄ?C��v�)��N4{�e��?�Q�[��+��n��D�v����k�?k~ࠎ��2�=��A�w@Ew ������<��J��o�ןQ�]�7dg-^o�t}]&���������+R�󩕖
�yk�y����4=!<��ia�F�1���n�i]��a� ���7L�)�Y�b�V��n5�D���w74O�7�y�m�D��ˇu��/���?Ny(�����V�m��Q]�U�i��߹Q�?���|)i�-G�1�"�*�žSux���Ygab�[��]�	��@����c)\F��u�'z�Rq~O���4��Z��r����t2]�dI���f�'�����Y�_Rc��qߤ��,�w�1Ήk;k�3�"���J]�WOM�\\����FNߛxk3��;f�ϊ��Y����D��Ԕ���Z��PklOw��[��c��P�ά4�+�F�=�R���F[@�����\[�?k1AD���4عh#a�|�K!K>4��5ZT>.�\l���8�a?�`H6�NA�1�����P�����	Hsn����i�L.�W��9���	i$O�5C,i�'=Uf��ަ��p�x��\GW��l�q8����u����/B;�Ӭ�Y��	�6�0ЀY	�H���������1��e,�KNs��lw���X`r��ՅH�6鈆�n�Uf�A}��$7@���O\:z��+<0H�+]��J�h��U�"�ɶ�� �����9G�yF������90U��!���<I���\z@>������ ��;cZxN���,2o5aJN�p�yp5s}ǉ:���MA��:�C�eb\�
~�&h(%-��e-�"R
il���ղ� |a���|�G�tw�<�1����@�r�}�$�Oԃ�[̰��Wi63! �-�6�<����#��:�%��a5r.�9����R�hn4^O޺8E;��R�%�Q2_�ҧ�����_$�$(Gq�p�'C�ni�wO�2Ms]�ΈK2}�o'�_�����@�k�G~�W>��c�s�7�K���� d;���w�s4쫵v�b�b�4�,C����0����P}�*@f\��vUO����^�Mَ�hpy���[vwm�ӫ�X+$��'9n��a�c���u���D6D;o�~�"Ky5�;�#���n�D1��|q���C�?�N˦�6������I*՝��7{��������:Q2�^;���SB֪H��(ݞ���|(��y6aa:�����`sO\
����K�� ��o�Xz�Y{��O�or3����|}��Z!�����?Gz4�V �V��c�O.�ȥVcll\�шa�j�7'������|<�W�Ƅ���O�J��L��;���>x����4Oo���*�Wt�Ҏ��?Kڢ���D�&rS����iņ�:��H��	i�O�)U8��\�6����������[�Z��tڜ[J"��vjE5����iMf���XJ�{�����TT����l(���b\�"4^f�a<�n�S�òXA�6W�����u(����=(7Q�z�̋�<C�dU~)�/�e}�_'ц�=cxE��3�&IPh�R�_Yi�}��Ӥ@����+Ѹ-��E�DtrV�"�bA�(c�M
��iu�oP��Y�zE�#�I�?ɧ臺���EYM��ǏP�kS^%w[E'���h͖t���2�>���Q�F�χ�r��I�'�J	z�(���ׇS=(�m֗�IPw˺�ݘ�O�e�!ɫ Al�I���v��N�s�`0�<�@�u�e��1��}�gyr�w@:��Q��3pe���^{�Z�9���������-���P;��pL����NƎj���wN!9��w�#(lɌu>o�>,L�G�����_H&�����������R�߮�1ߨ
I���f���D}=��n�V&�#��c��n�9�"K�(����b� $�`z�b���կVf9�tr����;ƒ����LM����GP.U�=7�$Z�WWv�F�т��L�d~�hn��7�l��%��w,���u�%�����'����lX!�#_s���nn�EB�mxngHlu+ڔKu�\,yN7��BH7�E��S��4���<Wʲ[+l(����.i���gڭ�� ��&�}��Գ�Sudb��ͽ8[�r" H]5�h�=�$ lXߑ�N����'ms����¶O p�| c���h5~Rv� V-G_�9J���/��Tђ�6wo�u�vn�3���(� ����k���ad����}6��*.�-��-���?�/Q�1��(�Ŵ�=�طH��,�1�~k�����J�Y� F�M��L[a��+-|�+g	��X������k%��5��Յۮ��{�)~?6�����Yk��9?�B����{4h�q�Ğ���������`B�rO�(Їn�@Η�d'��x����b�D����*0j�yy��ԣ���[S�k(�ڪ�_�
R�r�蕣q=~Z��r-�ͣ�rZ�����8C,��׾�����Tk��
��w�|�	!��T����Y�(�c�fH��ʕ�8r����K��5{U��(�m��w�3B L�pkm���妶�Q�ۮ$��i=�n6��CP����:4�F�U�����CCm�ʨ6���;m!�6c�=��v�b�-���_ݟ7d���'M'�6�U��ԙ$��f#j3�:7�H�7�v�2��=��?ޤ{N/j���xk���0K��������,d@��sbh��F>�����n����ʢK�\������77�{B�J�/����_�%�����Aa �ғ|�S�$��E��vH�
�.Ǟ୅#27'E���ބ�����27�)Z���&�@��d��`8�e8�'��x�5z�n�JX`��S�b�-���VXt 3r�5�"���p�"&2�~��E�d�<�^~�9��kv��f�23�m2\�:�%�~୅�� ��$���qO�}�jK6!�.0�(ό4��Mr(��A� ������&��`���`�ds;!*��eM[�5�,8�7�_j�Z;g��ܜ��f���"���@s��<|�����%;�0-�k�mY�P�4.Px�+��1(��FyE[���ԉ7�f��ѫ �_짱���sn;q�/k���y�	�#�h�z���uIQ��D�]�ji/�"Ѹ�xT{�[f%2d�6+�Z%zs�퍑ai�HI��*��2Y��}�n�^T��A�#nRm.��0yV� ���X��p�X?���:Y�*�8�/$�;}i[�$��}i�O��G��.q̀E?!��v������X�q�%���/<!�����yAĢז���=Fy��ڏ9 @��F9�jF��'�(���ԁ����{\5^t���E�刄�opk��Yz��;GEir�m�I	�<M�K��7P���1�T}�{��%��p�䭻Cw�;�?���劸vw��'���X��ۿ,��1�"�o�ǋ��l=��r�,�?�Mǉ_��Exĝ�+K���; N%kf�{���[E��t�b|���B��2���	BA)lza ��w`�����<�����X������v8��i��A���;�4��/3�
l��Lz36|#C:*�xIJ�,$�����c�H/A(x<�`��\j���b���󚜱,�6i?Z���Wq^��c�I�5E�̐�E�Y�U��Wvz�b'	{<��y��UKO;�%��]iH���slR�N���jY}�
��[Qhqz���p��E"�����CRkKw��\C�)K`�2��n����/S=����x���Hi0,�����N�����/�<�P�ke� �2���^K�-2n�	��SLg���sWfJ ��G���CA�+�x�A�0��pqu�U��^�P"��f��j��LK�r�'2��1���F����5� k��Ý
a4�5u�$�Z���'Ĺ|��^4�a��!S���I������ꅗ�xV�kz仝H	�8�7E��g�/WV�ퟒ��ў�̗���"@Tm/C>�-c��~H�;��
=��"q��so��P�-�+}L�r� W*��A�����g�{M�A8|`�b]���A��R�,=�|��6w�����_�.A#Xؠ�_T����YHQlD���j�h|�ty����x�mZ�D�W���'��S��C>O��&��"�#��҃۞$5��&�?��l`A5�g�7pm)�ό���6y���]�fN�#T�1p�%3�(,9����zp���Ox���>gRxX��x��06�T����s���w�s-�UF��a0�y���&�vbD�u\�?��`�#uB�iCQ��8.%I\�jS�}E�����z;[ž��%�w-��xa;k�!\�TJ`��$3NbJVN�WZ� <B ]`/����AI���>�^x矾-�z�T�?5�{�<>;��k x���e�����AĨ��*)�s^C��10mP����������%�U�_�ݽ��x�N�_�Ұ_1��G���`�����@���O�I��&��͊��+� �,�VR_y���
2��R���h�j�.c�a�b���7l?��ʗ5��R~;��]�wz^���G��L~Bv�f{g	e����w�����*���2E|��S�dR�18��(��=��n���L6BQf�R�TJ�>�`�M�i����|��!	�P���/�0�B\C�B+-jӌ#�G�`��r9�J]�p�ڞ����[-'M=�"���#̸��U=!x����9�ap�x�������J9�@=��b�+fd����#"�z��̙����2�gD�5f�\�}צv��X�����U;UF���.�07��Wί,���<[]'4���yT\$y�r�G1���h!a�ݝ�?�>���7ގ��1?D��Xj�QS�I��/혚��i�����8�|��L>���-��t�Q�r-��}��qXCQ�ˋ( O�Z5nb��狠��;��O�X�f������tS�y��V���"�������pH�~Wm� ~.�c(��- �ȯHa:�����f��fÆ�J,֭�ԯ<�I�eε��sۼ*�e�k&��d�ں�B��'d�Y����"!+dy\疃6#u��
��5���L��#�Z���A�L��+����v�,�8�]�3�,z-��|]�OF�i(B�u)b��tu}��O7�u��؇� ֬�#��]o� 3�%��;�@̄ol4/.���G5���(7��4mc��HW�FI�8K��=���_#͞���E�]׎!�)��,ZJTZKT��Ϻ�>���Ce*~�fQ�2m��/u2m���aԉ�}w�H������AR�>��M���� �iL�*�iWS��>Ų�{��|
r�������������Du �7[Ļ�Ŀ7"@��,�|�i�9��u���� 
7p]�̫0��B.i�z��[��ޱ���Yկ����0��D�>?����]��*��#�p:x�WUS}��|V!��N��8�l\�q���&�$i���c������-��}�"��P�_��g+D���Vw���^Lj�s��,FM�_�F�<����'��7H��M}j|�K3�����DI�[���eї��oc�;=��#B��yj�1�hW �<�4�c)`	�Ӹ﬽���ܖS��ӷ/=�_�*A���th�"/���_)kn@]���Ρ�j�� ޢv������{<��+��9�??P�=8���8�~y����VG���n�^ش]����7���qw�6|'�f���H	�7v�fl�m����1��+�ƴ��%�\(G�d[@�_�7]$I���Iй��$�*�?7��?)d�K��������(&&���+���q���r�`9�M��0�geHԿ��H���98�(q�ةX���Nۛ��p�c-m�	�aE�m����%L��7��j���g�J�H?�,;�1�DѻU~}׏��f�RQb.� ���|���u��o�n�����3�a�"OO���j7����%����c�ҧ����-p�今^|�N�������2���r�4�3��{��׎<<��=��o:bŞ�׊�*�~��p�)�K�~�It�W�D��;�l{�!��=��i3��Y�p���E(�	�U�Ӈ$FM�ۮ�F�q<�`	-`9��u��{"��a��m<l!����;+)�:�QIDCL�#�D뷳O���UŞ�W�n<7rO8�c�
�}eߟ���1(��ښ{�i�����.�_���p��%-Ѷ���s��Ie�D:Ŏ����++�y�9]��W� SQ��~M"I�>��Ŀ�8�Z�I�AW����>��ܦ;�)TW1XE�Hl�X{vtd56إlo4�V���/Gܞ��6�&9��yӴ�g>��r�+�b.h�$��t�/�ݥ}i�
F��9�?�G�##-}���5C�E�Îvb�t-�N���/џ�|��ʑ�:�)RL�1xzkT��ĝơ%0']H~��v ����_�ؿr͂D�U1��D�S?�`�t�9��t�cK�N a������ �N�"�Q^�3����|�g�ԇh�}n�y�ˑ1V������ٜ�d�q��V,.C�lt�4@�������;b��oSi?�8��\��Άx��-_@>5K���U���f��v�����MW�D�� ����Ӎ�hz�x>'+�%Jm�su*~h.aG����2������_����0�=s�>8!9^|D� �V�6����l|�9c��+_�}�a���Tͫ����&��֑���ˌާ��w�Mz���j!r���"�3]�[>&�?^�ʧ��hن�pY�ͯË�=5`��$���K(��!�WH���9�OT�t��ь�*O"�f�`7��;�;�T�#N����T� ^�{j�?���%�hX<��;�%{���A��:�Tmk ߴw��^��e� >�?��&;g��� ���U
\��P�C�!�:��c����5�P�8��cڲ����h�Ӈ�`+��y���]W";��n�����Ԙ�F�����J�PY�
��|vvg���b"/N�ӧ�B�k�����2	ߨ7O����>�N�7��W�tnQ#���p��:��C��Q��Ϣ�Nw�C��X�'�ֵ�\d�Y�{�$�w���}*c���_m�N̓�"0~��1�sX�Q�^$f��L���\��dk��Q�<������$gd����޳���I�]}�=��S���f���k;��5����"c([2���y��"ޘe[Ti�n ǚ<�ä�����ݟ-u�Z'����ٝ�Χ���*ߖ��,T����Ut��w�v�9�-�w��z^�2-��g3�;�c>�ߛ[$�-��Κ.�tۮ0^��^=O2L�Ů۹Л���A�d.:i����[@�����L=�8��Y����1 �Z�X�8�M���F�����E�rRa$�k��r�;/@�C�&���>,W[���i�l��e�=��?�b��(��Ұn6��-5B"��\0���e�z�L, ���A���|8��y|�:�G�E�Kn^x�U�(��5�d�Z��C���ߋ������6�1����������.W�0�d2[��<�E`���Hn�y`~����yBvw'��P
&mwP^�3T2d�w.���Y��f��zE�E�r��yf#	��.�A|�SG�\������n=�C'�m�ç��+��>��25�����'v��������z"�i2���b.X83`�����v�nKFd>�9�X�%^�Q2� �ᷗǯ�
�{-f� dԯ�X�sKv�G^&�6�����2!�U!�3(��A��Y���g!!O�΂b��qeqK��?��1�2?�-ɢM��1kKc���r����8Il��N�A��_��<�w�L��Z�΍)��M��VߤEw�#x�ou��[b���#���h��?����76/`�g.�Qo�k��"���������g:Gbko��}Њ�y��3v�6�g�5�iwC�ycu��ĵ�ya�_N	�%�nX��U��Ix�Ѥ���c�K��HLA�1m�4���Dl=��i�Z��S��yq���[xa!��h�&~�����&07���g�;�eL�7$AFt����w�Tp�6�S����x�7`W,hk��P�P6d�eg�c�wƜX����{�������j��#�g�.�N*��y�#�_�r8�� Ҳkq������y~��jcWu������B��[�R����wty�`���!K\�
��`UNo���{�,А"'�o�]/_C���
����lR�U}d?�;�?���941�G(\���4|�������n�B���g��y;�Lrٌek��e7�Jts'�9ρ�a��>K 
ʙ���L�M�m���Wz����~yO�� ���31f� .��yg���	��HO��s�Y	�U��x�_E���7Q*���ݪ�66��{Hd]����_PI�*y�%L�r'���8.S��AYa��䣩޾�7��� C��"���M�����I�濸����3�v�C5��(g�Q�����4��gȕ�����������`&��VZ��r��'P��ښN>c	e���Ƶ�188K�����=�(Z� c����3eA���g���w&�|�50���Y� %h.14��F���~?�TM�x��{�ݳ�&��v���@ؐic2��Co��4-@k�y2m�77�IJ�hm�0c�Z綖�xB �xB(�;<��6ٚ\���
�K�B��fq�N̩���"��f�ij��;n!��
�y�d��W�ɸ�&����$c�)~�5�\lS��9��~��k�;#Ա��!p�,�ߗ?��}wBy5�`nā���
���"�V4:��E�kZЉ$����H���ѭC������ɹ;�Te�4/C��;ML�T]�����q�1f�'�omP�=�%X\Y�n��C��cV�!�Y���8qG���@:�,�,)4�\i�2�~��0|�~z�B�3�=maX��^�R؏1�I�����1,�-�Y`�e�;�-K��6��,�4у�̸_��ְ\H�����73�wj�b6�t.Qx�v��1���|{�K�m5�q4p�~HH��歋�0D�'�z0�����s�]h�Ȓ���E�� ��:(�ܧ4��]�,���J�)�d����<�AQ�j|�0���VJ�=duX�����I�}xI(x���`?8+,�s��*�?#�q��G�:�dwԻc:R a�K6���zy�D���9;����^0�3���,�����W�������{u� ��/n��.3aO�\�"R�R������*�����;jj��q�����z�'���~�Zn9Yg�`by���H�ױ���H��^�1����q���3�tyt���ܤpz�$��GI���殧;b��y�^5>�h�+P#b<cW�?h�?ք0~ 7�i!?��s��h+_fNw��H�4�r�j���qAD�/�O][W����F�����+~�tYp�9�xp��׶H�|=M����tQ����JMAF\[�K�\����%�(2�Q=��jm�8�e	��T�Q�έr�7�w�4�,#��c�J>4�*�'M
_����h��+�j|^}3E����­Ք�2j���Qk�W�9RJvz�y1�v*�	�`��{�#����s�Z��d�Ə�l�����-�²�q��ۭ>�$K�����&/s~��ϸ-�T7��a�"��rU��G�o�����_#H��1�/6}�vA��w�/ߞ9��ví�n|�%v�Dp�OO�XͲf�s�f�@�@�x�n�Y ��3Άo.I�q�%?s��U�=V��пw��5��V�,�]�q��VK�I�0t� �N��TԼj#�z��ۛg��$
h�4
 .>��V��glt��K`EMj��'��W{� �%��x�� ��R��r��13Jv�+�z�fe"���G>qy�?�T���4���X/�.+��ױl��*���h@�_�=������x]�R�P���cTs1�F�ɲ�k�z.@�B���`9:3���
#��u�[c�l!k�}��ZJ�6����!pC�c����7��EQCdX��lj[6�K������lY<��9'���fV>�i���o�)G��D�5�C;�o�����G��>^$�i�����Ûy��?mB��%�7��eh�|�Go�TI,��׫óc 0�f��������Y������=�&3�YF��D,dQ�W����n�U{W`<����CT>��R��)&/�ۤ-�t�h��]V�g㊍0���vg�x���H�I��W�_�aH(`?}+�g�ӥ�{qj�<EE�D��Z�e��goٺ[ş�a&Ӕ��,e�۞>�;�Q+/�Ν�U�G��ܲ5#�����M��e ��������n*mgؠ�T39�%�C� ���> u��N���N���x��Bp�q/4�ú{�����P|�M��b����yr�����v>r�j���^�t��*Y,�u�d$�a(A�Z�X9�s�<Xt8F�������<���(,pH�k�z<���L=�e1z�HVa�$'(�Y�N]�5��@4������ˤI�rX�:�w$.72$�-4�h|�s�Tk�N=�wOL;h��N�&��N�=\\�,���:Y6�j���ɥBY���ٺ� �׿}\�Wi��%Ϩi�i�*ü��'�ú�k�ǌ��mT�B�/�I�1�ύ5���=�7Pw�v��'���֮�w�Yp��8�3K���9V�Km�S7q�A-�+c���)R�����dٵ��g��Vg�8��q/@Փ�ZE��2Τm��ٔ��X}�kL�a_��i,���o��B�md?ѣl%�j	�� C~o@N��P�Nj�k��gn��������a7�[p>�\ �d��X��`u�,�����f���J��O�6��s5��s#��h����:���x����7��.�0>
����z���]���D��u/�]D��䓲��v�c� �����>g�'.������_מ�:���}�'z�ω���$�M�����T�d�=�'j�q'�:�?���|Y��,�*;l�}M�V1�@���`�e��2�+�"+L[OO�����~��8b�� �U��������J�:B��B�!�J9�"1�!1g��9���C�P9��36�D�q�4��|�m�3~���|���}_�u=�}?���:���r.��h�H���u�?([��:�i|皚_��̙�5Jo�,V]�O�Ԟ���G5P����,����q�V�����������=!��N~��L�O�ǖh8J��n��)��_O�~ù3�!JГ�wy�v��ST�mͳ*�S�̀�:��3*F�G��E�D�)�Dw���N��]�|�����̯w,fqQ��mw��
�Z&��sw������>G������n���^����*C��b0?��S�x(K�tZ*y(�X�ɍ�'�vKN�t=�N����|ju�4�v�J�׼�]��Y��_2�)>}�u�칦��̪Cq^Ý�5]����~&� �nz궤��Դ0�p#��ZѮ�6\�OOĞxv��Z�q�z��%��K��t�28Xt�W�pJ��锳簿�����R�/�Tl�:��s��|�n�~�[�-����[�ŝD��~0������l���w�; B��j�g-iA\>[�z�H����|G �5��q��^6�ƛq��q�)$2��5�r+KG��c�+*Ed�2=��fI^����~��%8�RR�/!��xb;���0���V5~p|�^��,���89	�����]�p�Oy�lפ7����@���8 ��cf^N��oYI\���4��tkޡ�w/�
گ��S�>}��Yġ�j�����K�g��/�gx�uD>0G���Jͷ�WF�2*��"M���B����v�L,���bs�)��?F�ڭ�kf����yH�����L7���C���R_�yg����?���TJ��&i��Z�|D�|��E���:��Hv�¤��0�v_��|�N�^ԩKTQ���%OK�H�x��$���[SUx"�zZ�ܿ�N
竒�u���0��| ��9t#�����2D��YMl\�"&#\��/v�ԕ�3w>�x��.����ԍD����.����w3R[�,i�CjW� ��[yT��jD�,[�H����;d�EPc�L7�ז0�
�Vdl�s �K3�.�dձDX���X?�H�]�N�,t�Cd�[�����"���W�;P��/��(��.�Q՘�ؖ ����*������w�*�^���}��hޅ��>���G���w�C����]4���+kz	��R�pvn�9��XH��~�\zwSC��pT�ş8S;$�V��zc�@t������?8���{�4�v2c�[.V�aI0��\h��~l�DDخ�T�%1��ދ�&�Ş�v3j�JJ�R�<v�;�׏�)7؁\�1O\sa��T������_�:�U(@��<+�,j����sȌ��/L+]�sxO]T`
���P�:�����;�7(�p���X�fI�Ox੠��fs�CTpz�j8uE�]��(��)�9�P�rlzИ*�ܪ4
TИ�}�˨������*$A>�@eˮӡ��ڝ��_�?���ԥ#V,�ވCLZ�$'�#�r��u��1�DJ���T��m�e�8_8��;粞{�0&����{�m�Gӭ�ouVv�OR�����2YUN
�Q��0Y�Ip�B9���I�D�>�>�S_y��xܿ��$HqӚF��!��2��W,5m�G��,hWk��`�+K����f���)�p�y]����QZx;�����w)��)�}Bs�5 ��|�2��V���< �����"_έ�����ⷔ�ďE�=��>}5��%;͗�����K{����/��Z�����z'
���]jǠ���T������O��t_*;]Ӌs�+��Y����N
��!@u�%*p�{��	(?dh
+�G���i�I���'6�ey��,�/���/�����Pp4wƾ�8-�����
I��S����i_�KQD[Y���V�������'�L���;��dq�㵋M~yXiz�0v_���|���a�[);,�Q�9�7ȣx�Uf�ԛ.�3>�W-�U�w�<.܁�*�Q~�?���#+U��� bm}����h'4Ya��es�5*1�!"�ϗ�&&��x��������;�dg�%��!l����.6�����<k����!�^y=����u�Z��Ɨ�����[�]z�?����v^:Up����{��$�5���?�Yǲ�:6<Z�#M���!��o�_іbz��9����d��.�x��kZE:��9"�A�r>��[�2�E/D��Fe�}�st"�Ъ�x������f�/E������a
��)첀=���#�T���c��h��f���j���!A>��� �EP�`k� q�6|8%�wc�t��w���;��Т�Kj#��ճ�7�j��1-��8�jm
Ms����%Rx�����ݼm��{�����o[;���/R��	��+3�}�^����eR�]��tZ���Հ� W���~� ]�F�c������X�������SO�"��Se����C�^	7��W�Ao�_x����N��d��<����p����(!Z$"[��q_J6�/��[P�<q)|����[)���>�&+��C��~)�`���Oz��HC#/��	�s�;�Y�q��3�q���#��d�ߣ����u� ?�=��.��2T���"eq?��@��U8�S�q	�xT��`�ZƖK�YO�Q=G�a�^�[O����=J:�tZ&N��{}|)H$Be�0x��Y���5�$��+��P4�ks� ���2i��n�������@Ϣ����I�}����b�X�B�`>_>�4�3�[��\�q��j �GG���:�󟈔bL��$�~��]��7L�Z߻d��y�j��UR�J>��ּ���4������4b{*��EB�E����&rR���9����u��w��Υ�U
�u��^k*�*U�t��:��C�d�%w��ݫ-�N5��O)�����\��W���2�݌!9U
#}�nM�W�#~���j~�ųKѐ.�nr2j�h�A�F�0��&���w2���o����x������3
�]~(�0/:+1��l�?)L�I��'�h��渆����0�)��#�KT�uh��^�;d{b�Y��$�dg1/�ϰ]�[�xU��NV �|Jk=Uч�q}�a@����$cKh%�Mt�[��駁��<����T��CM�x#ޟH�U�n���A�G=a�9���+�l�<Z�ٹ��4D��{J�*N0`��'��мٴ)^�Ϣ)���;��%gl�We���Q+�
w&�w|i�'���A!)��XZ��A�E��k����� �RaN����J�4�9JV�Mú��)D������i;�|����g8֯�u���9�{L7[@(2[D�%�T�SbL%���=$�h�N�c�8��6��8����E��&mɯ�E+(�m�,;f},�{��:��LuȄI]���6<�9��B��E�C�{�6����á;�)�C��0����;[�5��a�ȯ�//�Z�)��5S��t��K����GB_C�YS9:��;�mcB�b�tڽz�*��@M����%�8� w����C�cQW*�3�^�.����ap:l��������K�`���ü��҇�o�SWF������8�f�l9Sqs��M���1Q�3(���G��UV��!�	�j0�������{`ܽ�"���#;�pnb����PV��\+T%�N��w�az�Q-Iwz?��m(s���<�O�j�D����}��y�N8TE��	���)˗�G��JJ�3-��	�[�:'G�t.�]��j�楤����}�N��݌��ej�cq�(n8�K����ۥݲ�w�֍��O�����N,�R�F�!6,u�C���f�V���w���v���i[���8����,d�3f�RM>u%��uDPo
��l�6
�|Ta�����:�7,wk7�Q'�T�jg�.�"[al�T�_���d/斘�����7��#��A�e�lu�!�+��Ot^<��C����GJ�����4\���*�hξ��|ŝ����WP���*z�L)�1KXeH!��~|������qu/M���c��ſ,�e���v�+����\ K�'94h����-�Op��dȈ��Y��ۣ? 4.�]��k������6���g-P�9�a�����4vtF��5Ĉ�H�/k�(��*�ΰ����׽��)�G]i}M$�a��Ҽ�"Ĭ
~{���K�ym����CJ�;/�ܨlÍ���x5߳6+C���7h�P�?�6��"�B2����YP��[!�9����'�#x��ͻx
>��(�[I��9Z��R�(��)w�?����-c}�#�~	�Ǘ`�ϵ��P�8P$5<w��>�{���'Z�P�e7of�xE+c�f�9��?���F ��>��>�<-Z�Q�Q���K?*
[_��u�!B�xɩ�Q�
��)�� ���1��O�f��ͺ�휗����gPg�H?;i?OqӁO�^_~�2�r7�O��Y�Ȑ� A�o��ȭ%�r���a����H\�?�;��U��][࿗�	{�����5D��`�u���������$$.���5��� �s��J����i�����噍���i��^�-.{M�LX�a�m�Gy�(��W6`��.N;��aQn.��-�D���{Y2o���D�\��j�a�)�k�w�fO����ػۢ�.v�,�ީ�Yi�������Vu��YFâ�?��5.��S���^��_5��F�g�6[!���u�ܬ�4��v:M�J�}5��4�T]x�~�#s���vl��awH83k ���[��J.�y������x�5+��4�AR�I�v�m���\��SNJ!��0���C�~-j"���F6��ID���5E|(�z�E?J�SN��p�B.34�������o�FwL�R��Z�i��g66Մ7⛺��hH\����=;Z�x��MI� m��<?���i&���gֈ��i[���� �Gk�,-l�V\!����ͪ���;��{0�+���1��t[��<T+��{.��>!�T���u�9� Eh>Ye�7ཀ�ڡ�8@5ir��
vjg4�����S'��S�J ?���$!J6�=z��~�PGe��?���5��ZV�;�k@�"��:=Kׁ��-�^�L���9��*�۽��z���������:����f��HB^�oтO�)m�m�!$J\�]�f�#Z�̨��2��t�Ԧ��Py�۴�ڈ�*���ԕ��J%(@lv8S�&��
j�`PS����Z����a��.�>�0�� L�w�VŻ���o����d�Qd��k �Y���<�K�a-H�΍^	m2�(`oNxQ�^Ӳ���N�"�^g\��IQ���$��/�]�8��4���B�Qn����o1����Pf�E�>�X#��)���n.�>>g>5��G�%j8�5+_�ӟ�L����u������i����6vX5,���鮶V�9$��N�Yi엽_MUm�5��A� �1��Sݣ�n|Ѭ����w�jA�+���#qx�9�C���!]�C������8�8ST�:���BSC�N��[:1Vj�#�`��w��<��k^�c����2�: %(^�l�C�U8�2��	x=v�T�7�g���KlV�K�juN=��g :[�"��nOa	s��7�?-u����Y��g*���ΰ1��I���L���1Qe(�c��w�%h�"e��ʦr|ù��*�A:1����lv�'|��2�	
���l~V�=?+�#�g��"b^sg'���M16�[����a؞�*�Tb�LD�-��(3lm5C	Y�ۛ�_�.���mQ��"���Ӣn�.�>
+��������\̴t'��D�=��G�-�?��������*�:t��+aX���N�N���H����ۮM"D����%�a����C��U��=Yݼ����'�[Y~�F�3}U�^��E�w$jҕն���U?J���i�<>�������1tY-���l` u�4q�7v]�ޏwHs�nV�\� y:
U#R��M��`�W|�wkMg;���K�rn���6ˤ�M����>P����ǧ���Uu`����v�w����|���\W��c�n(���F?�p�^AHB3<��wzV��ޟV��˦�&�\Q��`ҳ:��l�NT&�6��M#R�@��KI{+2��+�qvL��Т�ֶ�fa0MG� ����9U�W������A�'
eq?J�lVH����`�����SOy��pZ˅���cט�B�x�Chk��`pp�hqR '���ǎ��YH�q���v��r�L���T�C��֢���לӉ4%����/��	B[+'�K�dx�/��g���S-s��F��3���_�/>��15�d��t,�O]�h�wG��&	��	)/��E2��R(��Ru%��s�dgԿ�?|$[��g�278����8�z��Qi�_kܤq��,���#wz�	X�J-�p���!P�ӷ�3	q�PDY�_� ��+Na��.�K�m�)�?��u�=�0W��к���s����k@-������YZ٫n�Ӳ�rj�ۑty�B�ma�X�W�XA���}۹B�>�4���F�	u��*�x"|��)�G�wS��.P�]����ԕ�������ym;)>�3�[���$>R�31*џ|;׻���CYĳ��H�H��>#y%�C��=���mP^ �ҫ�K�.n������_5�z
�Z�F[��c��"�Q�_c��)?�F;Wn(���<�./�g�YfIDߒ'��7x=�SO
">^]j�)n�����e۸}�3�%ܙ$�����Hz�1�K���T<P�� ��B�T�d��L/5�d��e���a.���Ċy�o�T��S(���#��Ƅ�O���!�~��A��c�}�"D�z��@�Y ��l`2@�|��I�j�Ә��zͬ�H��
���4�u&2���/(��nW&�YZJ����q�1�m9�~��>����	��5��(%�R�ysRǲ9wvv�`��;��ц��5�,�HD�Lx�n�B	/���!x�þ7�۽�|c0��UxJ3�.i�O5e���:XܾM�fa�<S�ƴ�2�l�������7!��/���%����o���g���p|d�S�u��c�%�gb�Qp/u�~�\��y�M�g�o"�F)��.ۨ��8�3zp�MoV�JRĳ�eѹ�A�*3����`�� 3�~Ŗ����C|����t�Nv�i�tV+ix)ᵵ�2CV��e��օ�né���u]G~��o��u�Yǒ3�fF�8������=���:���������4���_D�K�	�Tl:r��ĺ}RԻ�oC��h����3������p�%�,�L0����E�D�0���-�HX��pN I`6���*�{�y���w����3QUƔ��S�p�`+�O��m��Y�'��p)^|�G��p_**��d0r���P��N�2��ɡ�S``�ela�G�n���#���R��`����@z��;ӛO=7�1��~����r���>!��&����W�f5'İ
	�q��VE_T�{� ��4���S�A�����;ęp��c"������K��Fe�=�+�� �$����^�v�W�`�>������潊���%K�02�Tu�|�p�Qu�|*�c�3�& F���Ža��m`��`��L�I�qS���`m�iy�*�g�оU��| SP�.*��%�ӳ{9{��1�;��s�j��{�V&�Z+���?k�������A���m��	s)	H
��"j�*QIȿ��;��#�[�Y�4��{�ѧ�W$R@x+We��i4$sn��viD&��v��E~�/�y�$2�~~����|�R�A�_���� |�*���eg�՚��n�,��| ��6*m%�MR���
��$�%q����d�Q(_��⠗�׉Z��۩$&���z+x��N�}���+5rU���u�w�_~�����/Th�*n�9���'�Y���i$w�>�����΃�o�J=����E@��4�wi�?�7�)Z�M�eq�� ��	�!���x`�ax�j�EG��u .�oڒ�˪\�yv�F���N� 	�[`~����E�Қ���1��Y@v�d1�����%�/i�k��?�{�T��kK�mv3֙���F�����7J� s��l���;HGj�7�K��������tʈ�sO�D;�窙8Q�����?�e��D�
�͐7�k:Z�0���|��-G��������@f�~3zA)�O�4a�;Ƕ��!�\�UW.��ej�����9�YǊs|�9��;'U�M������1X	�M/L�]߰�[���o��>������4�)��3��~�O��������HB�5M���,`���bF��H��5����;���IW����=��;:#�>��Q��I��<g��[oP��a�֤4c$�q/��ZS�%-Oe�Z�ƿ�8}��g�t}E�a9,@����M���?�H�Getǎ�{�q��@�ُ{��f����m�wM�6����'� uȚ��"Р����i���w3�7%R͒�[��+��O:7��q�'>#��=��:�d_,4y��J�
�6_�R�I²��T�l��pAʗd�S��.+�}=�)6��7�Y�0h����>��1�&<n�B��qw�iK
<z�&`�v�񔳧�#1lȳ�0yZ\�l�;sI)��.�2BS狽X$r��u��B��a|C����/�����y�[�**ym�����E3�L����h�i�|{�|0��F)Ü��r�P� O��;[�M�흲�i.���*N�qA�L��MHN���|���0n�p��k2+�=��RR�p��v���&s�
FyIq�$�i�Oj�PJ>��Ny�����_�v�2��ۚ��3�>��o 	!�;���*mֽU���
Q�Va���E\[sF�˨�����ub%g�.�����i)<�g2;k��A�������R'����*�m�l	���'PR�jND;<�&�f���󴻧���ʷ��)���Y���񌏹z���٠����#K�mȝvg%�j3MAr�+TW]�CE�B\:�N�}ՀLq��پ#O�{d��k�܏
Pvm�\�f���nn�]ôB�.��g�YƤ"�����K^22�KR���e�8��a�_�w�`N]*�x��j�����D���w7�{`��ʼ�yO��������!���z2����F� ��}�E�Zː���t���Ӱ=�i�n.��2`Y]
r,�6��I����ˠ�d�ѪtuH�.�å����X����;r��d�T�7�wV�{�ӑӻw3����7L��O[�a�'�^��\�s���k��Z>y���mɊ��P�8�+ܷP��� ��6��l���`30`d�5��ߓ�� �#������� ќ�1p��D�_���Nj�\|:��Yz��k_�~���1)���6�������'ꤑU�)�3(�aD��q�g�:X�`�_��u,�-l�� ��iM-�<g:�|�WRp���Eˈ)3�v�`��\l�I'9EM��yM��[^Q;�ha��F<h�G.$U�G���.���8_�ž+��Snj��]=�V����>G|=G��N�k�_��nuT�;k�_j]z��dy�V)^u*Tu�۰�����,_7�a��N#��<عf<�r��� ?�=�Я��_�V�bV�:�u�ir����ä���E�u��� ��Z��?��@ΨP3��0h'@xd�d����l�U������������{ ��ߓ;�s;%�꼢5
}MN�?��=����P[ּ�`tG��/!����}%w��$�N����DO�2ËgD�3z@_[�4���y���jw�Lu�x�ܠ��0�[�8G�$�i�|���=r��爰f��h���vs�hD���.�xWo�Z��#��A���j��{��t�W���U�
�W}!krc6Z��3�ji7���&�V'Fķ[:
8;t���(���x*�:p�J:��V%Y���Q�y�yJ�"���R[f)��U����ј\g1v9r�k��TNQC�hH �v@t�l\�� F6��������I��;n%�n|tT���8�aZc|׎G��Vw�9���c�:Sb�u�KPA�<���d_�f�%�*�a5�����j��k<��������b4���_�΂l��أ�$­�u���3W��5G켊��ރ7�u�/��Q5!1 K˶kj��q�s�G�_���]�����3�e�Pg�A�'T��0��W�
R�W@x_��d�W�*J.T�P��{f`4�2e&����'Y� "��������՟�����t�s�C��������0�Hi_��(��{(A��2�V^Mȿ{��Z��!��޷����A�����g6]�CAJp;5�w��������<Eԃi�b��z� �Jr.jec٥��q�KDbקB����n:"��_������LZ'���v�w����z)�bd{�)�5���N�jg���_p�n��A���x�r<��RE�x��$���z��=��yQMk�����w���@NCi㎮��[:�Os��
�������2�`꫄QF�	=����IC�����s'���j�� |2�ɺ؛�$"D%�E}�ll.����¼0�w�<���6XO��(�-rDQ�=h�s�-v�W_�c�T9�jQT�5�l����O�2�B!v}���Xk��Զ��c�q���_9�+%Y�\t�9P�˪�m�lTI��&�qGL���j���6��¦tDP����ڽ�?��<L:�I�Է�j��oBu���@ ע���?��`�7���k�91@�3Q�Q��y���7�ئ�����+��#�D��4��ƺS�x�A/�@��+c�3���K�F�&��-���O|�(�Ձ�Ҡ��V��"�o1�T$o�jM���E����7�T��Q�c��#���w +T�?`�[���y�C�Z�����Sz��^R҉��?l��	�/I1A?7��Qt��i5��U����%`��㻌��V���q�΄/¦�}}V����{��;�C��J$�������(�e��"e����q�V��d����D��J!�HO�N�'Ա,�̺,ٵ�f14op����*�!�pcF���ŃkyO��UQy��ͮ�F��.��BK��Dl<���>j�cd9+gW5m�"��fl�wK��=��m����Y�ʶ"�
L��\S��I_��rh-�/�b�Fm�S��/.��Wld�{˹�i�~�	��V���=ۺ�X?�Æ����:�L�!3�wj�����*�BK�֬�hRs����e(i���W]Ew@\��������v�|��nZqS�985����1���[�K\(Qĩ�����)�֗�W�X��=��7��m�ˏ�Nq��t�i��k��0eƺ3�&��5��Z���Mf	e#(^�3�H�Z'yk������3��|��bDo�EE��6Ç>=������&��*h ��/�V�`1>ۀرk+�נh4jT�> v�)�b����[�[s���Y!����ogk���ߖ��`�}�z�-~y߫�Ϡ�U��)~��֗4�}��_lYZ�vo��k_3��	^��Ăٳ�N�w�r�t�o"}�-o�d}Ŧ$0�9�0�IMx�9a���䙡�Z��!P� y�+d��4rS$��it�h�Z��7 �,w�Bh��º��w�-�'ڕ��1��:�@�������"���[�5�����9��Z���8��8~ߘ`E�"WV�Sy�����_9�c`W���'����7�S� {�*2��N3�\���֬�SNR܅�������Py���G³<����|e���3!�]��C�
�u�@}_~V��ʯ����KVV|�{sGɈ�?ø7��K���0r��n�Uc��!�1q9GU��35�ӡ��%��#/��>�:}��ْ�.�%7��F:B�ʻi �Mn0Fy#�����ɳ:�sM{�0���������c1��]���GBb�ƨ�[�ϻm1䱔[1�����	<�8�~���on+�E�MU3.����zڮ�8n�3�N5�>n�1�N�Ɓ2#H	����������Cp����i�붥�V�]T���m\*�/����;K��k�u�LV�o��ԜMU'�D�݇5����L�iM��xp� o{Y2jqK�D��X�p���&��(�����?���"�X�,K� QvB��B̖�Y���3j˅+�B�'�TP�+�B�Z�O�C"�L�H�>�` :�U���{�TX��o�H�3_}	�|�nE1���Y�JU���_�`~��w��2{
c7V�`v<��ּ�J����l�(9]�o:1�0��\q��v�_Y�������d޻��J=����s��QW�d�j�k��6�V�e�s�F"��z��/'�ɝ����ŕ�&ↂ.�0֏}���ܴz�r���3�8^�����=�����H�=B�/��@n�9ޘ>�!�e�ޏBG��S'x`Uj�=,��AZ��%E�W:.߫4�et�V���3���)��xW�J%�r��M�P��Z YV��Y-��y�S��	�&.��p�?M�Q��P|i�B�T�/tf�k��>�[.7XG�1y�9�����}���i=��#+u���Z:ߕm/�xZ�D=X��4�v6��i�NU�e���` �b��G��T��ӊ��{W�XQ|^�p:���O�ҹ�-�e�~sҪ�鯸����銱)�Wc.�����X�G$��(�ιCqs��I�<Įj^jd���b�x���wC+�'A������(`����um�o��h�iSՑ�cO�PYt��SdM��>�*:��E��O�f1�s��1�7�^���l�dU���,�\.��G��d3p�f�jڌ�x*[`uJ�S�v��]PM]����L?a������F毠�e�JGU��X����Y����z�mB��zKsӐ�ܸ���JN��!���Q	��'4�[w3��[���e��޽��'�[�_Yj���Xf��7�F���R�(p�q��I���z�����
�v7�i]_7Ae��4�!|f	L�����1Q�}��Y�I�#?O� ���q��׫G��)���i87�0��$W�_;#��R�
z��]�\� �}���ZP�4�������nf��XV�w��)����F>kX��s=�,�9�(�o:{�ӗx����}����"���e�ڇ���C�Όu�S�^r���+O� �~�c��0b1�v@���*�I��7�.6�)c,�S��gR���E��/$D҄ޕi��ێ����3L�߼�wz���E���&jT�f��z���k���KH-6J����W#�S��)(o�$[̚7X
oL|,�s5�Y\O��ܳ�
M�\���b�ύ�a߃�#E=��!���=�)2[����^/9���S���\�c��UF��4�B�'������@u������t&g]rH�I?첤/dG�THm��c'�fԧ�FA���Yd'��-�8��J�2�h�$��h� �#c�Ym#�"B���K=���Ry�"��s�+��p��/�p���b鍄�k�,.��׬����q�g �w)�ї��!Tp�9�t�T���%���^[3'�Wg[�?pAˤ�-���V:Y�b�_�9�lZ��3-�u�M�l"�a��ֽ"��LG�+���͌��?��C��#*��Q��'���w(�P�vܑ���%�U�Z���]M�{�e��[���8�9�7n�����yrW��;���A~���oB�0`A�I��a#��3e�;8Ů�|�t�m�}�	P��>��4����
��J���]�V�R��حѬ+8� n�2�lv��%��oY��y_uY�b�'�;*�"k{E���A�G���������m?/9~�`��J}1�͎$Yv�r(̞�Ң�����f�Y������߉�<C7�@�Q�Xi��,�y9�n��S��p۰���,��f��t*CFS�xK{P�l�#f�>1�2|�鬂�|�A%�)ǂM�S��b�� ��ڂ�
�|�ģ�!���茄�3F�����Ґ#+?���F�u�1Rd�Z;�������;i�Sc�S�.�7�M�r�����g)������O�M�l�oƂB�[�'G�2L;�U0k��5��`��L-m��#X/�2����n�q�����s � �Yh��0�֧8��M���%��`@[+ڽ���j)�K)�g"�2�TܛQ'�Q�8�vz�SR�QdMM���Hu��;۪.K3�����{J%���	��9/���.��ԅ�P�����0�J̲�Kؕ)Dx���萑�Ƙ8�E�'�.��{�H�(����k�x�x�g�����;�s��
ͥ�]��t�f[#�:�]"����6"3��b?"�λ��� 2�)��m��+�F~>K�F�3v0o2�]R�����L�B�ЉɁ�����&
����ܭ���i
����]5\�R���9�0�����KfH��Ս@����u�vP�!	NPU����-�\Z��G� ��:�J���q��
�){r�Q����{p��&�N|�%������m���������;CP		5�gM�U|�O)���<2���4�V<ߟ��W��+�F�t��ޛ�+W�1�!��irNܢ<2�_��+����4�����Q�z�6��d�#��(�S��`2[<D���/��>��|5"9'�M�3������,���f�כuG����:�W�z���Cj�����kb�ɰ����w��۹z��{��ٌ�k�՘�D2�^��"���\[����eL�>���rl�	F�f<kD�m�I������ߞ�oZV�'�f�y��s@�T�mW���@ J�_d��q��i&����sh<�f �u�t�cK�S��i������|z	�� �;簃as�����\R�ztì��Y�t[$G0��.y���YUd+If߉��U�^Jѹ�-�����0���l^�JX�@\�Ǝ�烴��ͳB���a��F���Y��4@��].߼�e2�rdja���Q�3���kr�O?ra�W�9!�V��������\0К�ш�p��d�HGP���JRO|fi��\��4d���b�&2��:�F�	>����U�l�lf�Ȧ߮:�Ca'&7L3]��2�\��E��YQ���NW� zr]4����5 K
Rp�N�/��@�v/��q̸�.�����Z�Gc�<W���?��eJ_�/��ܰ^�ǰM����{:x[�����~�N��X�\	
��ݔ�:�!j�ƕ�^Z9|��1l �� &G�*�6Dt�$��p��@Y��-*0�犲�HSg�&���7~������	��/���!��s��PuHu��ϙ�й��B�+���|�!Í��C��T۲l�z~���f Mcz�<} �ݿ�+��>�#�+��q&,�)������R�R�4�9�ݽ�jV"�{'̆����m7�'����){�O�.7�;�-�J�܆��y/�+���L�aE1f%O�[7�d������!9e�O����/�E���W��F�ީFT�`O]��^�S�]�TA�*+��N#hD��]��"�!�e�9�.�l�Fy��n,_��!������əOi�W���M�u[Q\���K��n]ۚͰ�s��S�gEev�#������졚���Y��BW>L���o���9\У�-�>A�Z9�=h�ͪa%�����Lg����F앥�0ٳ�^���9]�5�~�TV�x�4`�!>�se5�0�|-�nσ�����2-gX��%H�dܖ�TەZl�tY�-��D��v���қz œ��`�/
 ��J+(�I��Gx2)5�4�8~��n�!�����5�"����<���}cFWܧ:�1:N~����=cqfo����0� ��z�S1+q�Y�H�ל�{\�i5'��;Af���������I��&�n�V$SRh���)�tV�qtr3�j]�tuN�*vyy�Zf��� ��.;X�Q~��E��5~������yp�J��J������c���2�z&�E$�7G0��[j �g�#��N�vҾ�ϊg�t%V��oZI]I�UK�Y4oL���N���I8\<~1����?�"3%�˦l�)f��?���D����ȄO�/z���KD	�6� kf��8o/�`�0~�$m���V�׷�Hm��Ծ�Z�����׏:�,�/k��������y�v��%.���	j���c��XhE��o��I���+�����M�?,۲g֙�w�e�Y`S[J����?�N��|):Y>�����|S��m"�!��7g�V��m U件�����?���LGP&��STۙ�ڵq�\F�k�>��?��"Zt��ѶE,\�~�*�u�h��'k�!�p6��sݒtX��޴��(9�8M�WB<�5���d��s�Mkr���Sm�/�f���nv��8��Cp6��,�N�����Kk�Bs�W�F�L��"il���1C@b��ŵ��8
� g�����i��� �ٍU��)����bb�H���Xuxn��H��>�w٣lo9r�� Qz��sl��PX$�`�MMӊqu��Z�3)5�К����= �I�H����-F%@+��7�pp����O�n�}�h"���{�<B$���<x�z=�u�1�/��呩���thu�W�8A0;��~�>�e�х^��j�����X�y|7c��e��@�K��F飯������J$��x�}�[o�������E,�AQQ�nP)��&!#�:d�ҝ#6%��5Bb�6r�����}���8��s��y��޻��L�po��#�M��"��#_BR��_u�kϫ�Ϸ7J�(ǽu4�^�y_�.�2|Oe�ǵ��/��E�W�`͇hlW�Ȉ�M��~XJ����1Wb*��qR�}�\��@\���\����Z퍆��nj�ԉڥ+U��Nu�c���Ch����!极�8�bƘ�����8 ��fζɃ�����ʋ���Ƀ�G�ubU+�G�8r�H���QS�����h�{k�k�O�?�?ZX��H%�����|Z��H�k�	�d)dF���SI��2$����!	� +�ke�����V�7|���	>ȍ}BL���%��o�{�6q:C���A����5��<H��c��rȜ`v����琯�̠��9�~y)���?��q4h�ˆ�I�/ӽ�J��z�Ǭ��7�4^6`Yf�n����(�[s��<�k��Ik��!쐶ͣ*u|�N�ڝ)2�r�"�N�����;W��tl?�;�6۩�SⅬK�vNC���=Q0�J�q�K-6�q�`:��W�����~�@��sJ$n��话�9`��4�C`c�J�QC�6գdo8�%���D᯻����[�3�J���Ux���G/�̚�8��In!J�D��s�y:E�?��>�I�_����v��tx�z�S���lu�Y��S@�4��Z�%�B����:�����mt�ʧ"l�X�����N��,39�S��L��� �%���=�@�+W�)&��rD�ڸ�9}ϦR������?R�H��u� �i>x;�)�'MB�zB�E�..�.���;ƚK���[�SG?ɼe�46թ��� y�G�ߖ�˳N�ћ���<�~ƉC\4k�1�Q%���! ���^��$����ɆL0�
*M"#�8����gG�-�:d�j�����������Ⱥ�����M_7���냷:R����5w>7J��%3	[�.fL�?Ѳ�I?�YJӈ�
ήb���S��[�5l���2�}<f0� �ͯ����B�Yr���p�]�S�74�٫BB�E�Yū�M]=a8#`�ekv�|�&�'d��9�P�1�BN�n����@�V�ѩΓ����V�i$Ef���;7�w�_��W������ T	b
�1�ݚ�|��	�J��eUi��Bi����B��N�|�(���->���ŕ_�+��c�w��fE�+�S,�'xLڮ\�����r�/S��n�|t��im'���;d��R?K9��N��W�-	ׁS�6�P�n�y/�ʗ��Zc�Y�=1 �Dt�Ovs"U�̃����6�궗��	�,�\&�r�o퇯 �uF�9��H��pM��)8�j3�ԇ��]��z�Ss;��X4J�HM�sQ�S�bcC� FՉ��-�R��ᨄ%��!�T�S�?�>�Qmb���F�5+�Ӟ�T��<
�c��B��\�jH�|4�k���o��館?;�ψ��0["7O�y"7��/�@3�7Ȧ�rb8U/�.�{y�z϶lENI�R��g��~Q���v(B���Y�m��m���,�D
r\∯����'�z.����;}�5�lQ��L�����s����!j����\�9�t�\	3�ie����������j����5�5Ե��F���Yc���d��*�t;Ƣ�Y]�?���*n:�����p����%�)��'!F���U��p�/3%F�o������.��c�N`gZX�nR�lfvnU$pYD0/�V\??�;���S��p+ؾpaJ�j9@�>jes���6�A�d��Юu�iHG����OD�T#��[bCg4F�&͘�U�G�2�5�L��-�"��*��m���Ut�틫�����Ix�se�SD�*�N1�8�i�:��R�]�Q�3� 1\Nb�bc+{�WX1�"g_�~&]?<ܚΔT��B!FS��*.�y<t�.�~ޟФSj���Cs���p�祝�QApNJf1 ��Xm!%#Ο&R������8M��kdDF�qT|��f���ŋ�����\�@@������h��*Y�9�G�8ŷ&�y� �+'n����L�J/�X~y{5�Q����"wD�u���tJ��I�pg� pD*�!�G�{d��d��Lв���"rI�����wg�K-� ��o���f$� 9NDo4�p���%������H�G���_�/"Rv�-HY��v�÷P�aX�Uv$��&�@�>��79�_5��B#3����Ő�/}�FQ���"�e��><�T�e�v�|�r��L�J�C��(ֿ���(��~�����,j���Ҫd? 7�w�0�:l�R��WrO�̢jw2�;�U��\���G2�z�&C_Ԗ;�d�d�q�a���w�a{P*�~�t��:=�	~ �o���zTN��~��w9�@v���Y&Tυ�ߚ����Z����~"Z)��\�	B�6����r{T���O�Җ~)9p"��@@z�$��U��@oURH���~��N������^?��y�F��Χ�'��=���*{���/k@�s�h�{3u�E.R\�����}Y��n����0A2"�p�f�w��R��[Y�*��r�s*�^Q������hO�K��J!x�r�@pc?S!f�^-�4dD�+�GDD���K��(~�:p�W_�#H�s�0ǡs�i�g�؁��o[��+�u��C�h��:���\&�[����kY�ҿ�18*����[bp+�+����vq�|�:���8b�)����M	�DQ���A˒�s��J�j���˄�w�����;#�Uդ�ճ�G�}�aY��C��H8��9���и�_M9~is5p��@OAE(�+����rMZ�CZ�����g��?ǯ�|���rCM��^WPA`���7�`�!��{.��,I����L�L�L^J~�L\_Q�MnMʙ�������ĺ��Wz�򉇔�#ǝ��,c���o�Cv�s_������k{�MK��P�>�����h�h�	G�:�+9�~5l�#_���}�~H+n��7i`V�mm�ep#گ�L�(	H��J���ɟ[pt-u���� �!qY�z���lU��]܋w6u}��e�>>��������l�$��ex���?�o)WO�S�<��HF��t�۱�$�旡��m�R��׍F�Z���~�x�7�?�@&%��r4���V��iur\���PF��u�x�P�����{�F'������JI�3�G`:�w�f3=�@�E��%M�j��UՌ��������9� 3����haTNڏF��9�<�RS�3������%^w���/���Ì��x���X}��ʬBS�*,�(,����̔�$�
�7���ϴ�n�V3��|�G�\)ܓ%l�h���O��D�9�?���Q��8J���-@<���7`�7�b`��`ݰ���F?4-Tn�g����(}4����� ����7�ʂ9�{\��<������	y���m\�ۥ1�F\��W������z�2+\MPe�����--�f�U�X����J�W��,���U���w~.B����~_���V�;o̾��d����xC��3/����r���4�h�k-O5��&��5���h�I7��J���n�����!��mkv["���^��|j�"�GC �w��Y�u���I����T��C9��l;�k��{K�<�[>���|��R3~�Z��=�j)�c���_���G����2Q������?���MF&���'iH�m҇k��݄�c.϶���-��/�k�-���v�\y&�y�� ��~�1ۚ��
ƟB����>��� �!o#DH�-=��>|�V��#��8��i���G��o8�O)��J�v��{��R�[�%�y�:/gWX� {.��p,���Y��z�4u�ca"���]C�Vwed���Le�#U�Y�G.u1o��|���1���ˠD�� J�*�?�eM�_��	�o�U=��,A�:�c�O���l)�����<E��HW����\�O`.,r�Y����ϵ �C'35a%��/��I$���/����꟮����n	���u�Nc�,���"ot|#6��&�7�W��W�s�âT����DH�}$vM^&X���P���)h��IO�o�l���4�ܰ�&BP\��uw�u(؁��LknBZ���Hqd����Jx#|�8�;�KIB�HX�wܜh�{!�,�	���ԣ�v�x����U&�(���t<H.C|^�	�������^S��tޟ������F-b�'��m��N����Ph$�K'�̿0��1�/HS3]�t$U�/�]��|
��7�e��ل�®�T��,��U�ڳ0�G�N�92��'�M�' 0��Lk�T�4�]��j���&�߼�W���B��o�k���.��!��Z�#���Р���/�Hp��m�����'/�}E~����t�ooBʈ����3�&���X�Uv~�8�h��T�t��e%���؀�����A��	�٪]�y95��g&W��U�j���0��@��şjTe��cìG���o�7)Q-�ؗL2?��}�=�PxF�&2ٲ�q
u9��m2�^��+2����k�ը�����^�P�������^�otޱ�� ��|:�]�4f�$ nrg�3F�)�*
�b^Ec��s�Yf+�
�Lε�����T�8w���+�P=���	����K6`U��׉Y�-��7k��=�����~nq�z1�K�����4�N�c��o�3�JC2_��ϔ����"FF�ƶ-E%����ְ:�����Δ��= c�1۲�8vJ⛥ii0>v���&�7��7����;�e���O��v�a�r+�B��\��Si�������R�������:YB9 @F�B� ���%y3���C��Nx<�x�Op�~ �9��{o2��R�kf�V��B�۵� ��,�8E`v4r���f����qX��)���Q�%Wa�����ŚF�pRR�X4@�t�ԅ�7�Dn9-�E8�n*g���v���Vw-������V�̢�̋;��4��"x���aY�6��L>���t���[En>�oPv{v��Qnv̠�q���,�\vC��^d��ZtJ&ǝ�w��]xgC���ٷ��?6*�vs����j��6���q������:�5��F��D�Y�0��ʭ�`B7횄���-�G���d����]����p���,a��8�����/4�!��2��Z�����!w�$�O�����M�)�4]��{� ����ɔʉM������'z\@�t��M��=�],���h��Gr�s%ݜLvu<"Z�(^c�3[��i^f��px���U惀�O��+`8ʗul,�y7�6� "�C�r����cN#�b(ZJ���$����[�l���;7��v!��/��y�n��ն�K.1_���Qʃy�Rw�����R�J�\�����O:��iI��[(@Ë���0��ĂNk=M��Ѵ�Y<���Ľ��9m��b>��L�{���U�!��)����$�������T�J(�u`y��Xm�(���v�6f}N���4?@�Z�=j��B?��ضB�����A��X��v��+���}?��H�"�P�#sI�/rS���F9Ъ�}#��LhM�hs�)>���f^~�(�T#[��#�}C�=��~&|_�:>Zjkp����H�/|l�}�U:K�bd��9Qu?�0��5r�;�P�H��"�USR���}���
���<�LE!�79�#��15��`\dq3�����"T�%��4�����I���<���J�Y�^}��#����0�%Y���Pf��@�2��GtA&f��M69-�}���}h��P�+e5���6�e�Y�#�lj�J�RS�e�d(�Vd��ϢH�d�8[6zp��w4&���1�_��?n��_?�4�9"ZA���B�������p��F��-��UR��(�̦�0��ڪ��y�F9�+w���= ���yy��I:�֬4��dqR���!gwu����6ã� x����l��2x}8��ܷJ��m��[����"W5��F<r�#��0i��FN�l��+G��7V�m��va�)¯�T�N;�fz�-�_�VK���ʵ��V�r+�F1�GC �b�	�4���D���Pt.aC���b�Ǡ� 9d��È�n�_��Z�������6�=*9;��	��o�2Ί ��i�9Id]S�6��\T?���ea��Zh�e�m��9�W-��t�L���o4����B]f�B���eQ�[�M2"�'�R�Rqgל���%�����j%򵴎�6Wov� Nx��q�"�f�:�v�ʭ:�u�Xi�K����a�C5�):��T��O������]-)F�"9I�'���2�b�;ƄL����ߡ�^��I��V;��5�BEf��%;.����TNT�n{Q;V ������@�e�#M����N��(;b���eU��7�49wr��#XAs����nٓ󺎗���R����pKAR�Y�i��[�K�K�! �����Čs	A��������p��r�\pS�~�����j�����N��X��ȪN�����ڳ)�_�
A�c� VE��fY=��iE�O�59�C^�0?��'�S�r�6o�d�?�G:�H�)5i�W�����[^&�89����x]�/[0�<�S̒�߸-+OU��\^wh����Z�{�}8y�����y�K�]���m��:�J�URB"Ap�^]l7�3ߗ/��l��P���3'\�������7��\۬�v�~���2��g��`c9̷�]i�J�>k�&�Se���+�*=��KN�8��hZ3.�6��&�n�]��b��J���z�c��/��N����?F��C�ٺ���1�|y�_ܜ�|64}
����r���>(�E���	+��o�V�v�Dqo���28����?��{�у�\�׹TM�Γ��}z��>V�i�aX~�$��w����Ss�^��L�߭u����!-���߆iDvj�W�M�W�ǁ2�S����Ž_�I���
®�5�O~z��_9X� �O�n4�կ� X�\� �EnoU��K���3���m ɴ���xǁ��=��:�ʶ�2 '���S��!y��,��N�a�maU�1JO5�f�Pؙ�p�\�-�ֆ��mH���kͱ�>C����yռz��V�z{�sd�{��49�iL��? �Ku �i�|��9���r����|���@$W4)<�ݴ;f6�:�����|��e�=;�ȥ���[��E#.��lo�{H��WO!�[eJ���-�e:2"ͬu<5��Ǜ���Y�\��>i?~?���po�n���Ї��C>�%�_���h��{�󝍮�Kb���/� JAs����G@��0!�k���Jnf۸����{o���ع!l��V�{���}4���H����*N����΀L)0���c�7/�<��2��(eR���UWb��O�h��{3�a��[+�l����6�N�5cShX�d2؎���ZQM58���]�}�D~���%����S��ɛ­�pe;�W��9��6�������_ɒ�0I�K���V�h\T:j �E6o�i 9=I|�.0h.ۺ�^c��`tf#�bBI�x=��������a�P�y��lM�s<����E���{&r\��=��*��9�N����N�y�o��ZVd[3�[[m�:��p����N/(�c�Z��p	�d�|U��:�:"�I~�J��Ǩ��3����/=F��JV^�>M�����IPq^���6�5C0q����&t����T�_�����5�1�O`���kwz_�2Ɖ�_�F��Jn���L�����M�L�s��݊�#XcAo��h�j��/0�(A|�_�j^�:{Lʚd�z�r�,�(}��bo~���ね�Ge�o��r�{4����k-�jqs4���T8j�g�;�=im[��t��}��d���v�p����zu����8ҰMҢ���Hz�߷�%眳��Q���/�<n/��Ҁ9	�M_��}˯>C����M��t���W��<�^���Pu&(��7��p#;�{�唦^R~/g-�l��^� ȯ�N��927g=���F�N�ӳ��R���[@o��ª���K��B��:*;��u��<2��1VG�(��Ŭ_�5,C��T���~6Ee2�����p8����ٺT��^.������K;`$j9!h�ѐ%������\@���P�,"��VW���۸�B�th�}��H' �K�;����N��:o�'��?w<X}�t_�a��]����u_�P����*bL�E��2�Z\�N?Z�8����/Ff+����
$�O�"����Z�IE��zi�P�z�z�6��O0��'��/H�k[<�x��Ŗ)�1	G`���^��qd&0��72I(���X���h 0�6	'�|����F�oB8~VDJ[�#�p��6z�3�h���O��O J1��'h�*��@f�x�u;��@�I�|[�C\?�/Cձ"Ԥ�Hͫ/7����k��"FK�n��W�J�C=
�3gTTj,fNM*������8Ko����gW^<g�Nݹaxj�"-�j���
O�x�5^��|o
'h�G��^4ى��L%t�_���%"��hSȑ�ϔ��������T`���.U���0�"I~�Hܵd�z����1l&��j���W�[��{��-I5.b�l.����j�֯>V~"���3�8�ȏ�✥}լ.�3aP-ˈS�|��y���T�Lo2���t��@ܼp�a��2+�1�L���З������0}>��(�M�3ɩJ�����A��78~�A._0*�t9�#*`�S����N�/V���#��d-W`7,^��2���}�c~>C���T�}{���>7`���� ����=�s��BI*QNa��l3/��jN���@Ff7�ٷ銭�w���_F3��D!IE�E�.��>a�g��) �e�2���[���R�wӽ��>�fY���<g��z���߼V�Ni!*l�6�t,AƪeͲSc�C��~��f���պ�����6*<�6�'ɨZ�r���Ő�]@�Y֎	g�Q숰{ �V*,V�3x���`#Z���wyN��m��>P�[@#��Zŭ�[��R�f�+L�;�Ti�:2|��� M��/�|�!U�g�M��_�-�\����I������i�?1u�ʢ>͍l �r⨾־��%�S�^[���_4G����Zz�y�;��ka���3}����Ȭbh$hQ�Yq��L��ei B�sK9������E�=�V{��o>-�
� ���F�l_v�o���ž�m�A�c�k�\�%�.c.�m�X"�� �>��A%��H�	�;sb7�^`y�I�jyZg��2���(xΝ����Y�p\H@9��=٧L�xϗٞ�3�_V̩��ه���%���|z\1Y��s�<��x��g��_��}�}���t� ������ߔl�671��P�� �����v��xO���D�5��r�;Ǆ~!rc�8߻=!��U���H8��̝����ͱ�Ά���te�7�F,�,������}���o�V�]��s�-��;pc�n)ŬH��*�����xX@�wn߸��*��=`���%��C)b���32�x��}�����y�{���<\�2-Y@�R�`����i�V��5ĉ��=��ޓ�Ϥ�SF��l{\��G����o0�*�����Vƚ��&f�R��t��P��1��D��������;�(�+�+n�)aYf$����wn�l�tރz*��(��	����_]a�a��H�9��-{l�Ȕ�'�:�>T~� a٪H�.������&w���12%x���m�����ÔA�,ȨZ���&b��_Dr�=���MD�� ޫ�+ºp�����0�m��ul*��ꚹhhPP�Il��EN>���a�Vg>��쪌�?��������I��5�A}��f�Pv��m�i�uwܡB_��I�C9�5`�*ﯡ)�m���ŀ��Ï�������x�N���KL������%\z��qF#���N=S�6��z����s��r��d,�H,m8s���I|z���$��|���޹]��q�+A�����5�i�:x:2"F����P�l5�I�ǵ@^���З\0ۜ�p�,}J٩�qM�K�
P`ԃ߲4%]�Ox���繉��%N����ҏtm��<��+��[ps{�ȷ,� I�Gx��3(%�%`��
=�c��4# �!�e�������6_c!�=�y�Se�$r�k�'oO"���
�+Q&D�^Q����xM�7�Ĵc����ODc�a���D�������b�H���;�8�!���@�H�6�]?do��g� ʌ_���pih�$`����:!=���A~�o�	)��QET�7�v���<��E��U ��V��_���{؍M��5-̅c�ܑ:�� qώɠ87`棙�WD؅�Ua�U���R8F%��w՛��q%\����++j��]��
l�R��N��ӗ<�W���]TsK� ���?ʎ��=�X�l�&U�]/�MjH�'�
�"&F9@�p�����8°)�h�P��J~Q�L^�7����6o�/�r\-a��(0D���� l���۞���ݕ�wk�H6�!��3�=����D�V���c��p���ᕈ��G�L�����ŃrmJ:�>��/��N��X{9W�.4]O���2S��t��6<��t��qNF͞[Q#��-���ޕsD��D��U�Z�d4W��_s�W]�N�|��)� |�8���u[Y=
���S(&���Ig\��F9�:��G�SՂ�Q�(�K���5=��k����z_�E_�����&�#��C��XT1[��/c�*n�������7J{I��n�ulP�,��F,��OJ��݆;��[��x/y���E�J�_)�{���+ �al�=ʱ�O��(i�_�����S�bi�q�Y��[������g�We�Wn�������`��.
����`�P�M�h�o�,�'��w�Wl��NS�� �]�|dp?]�����H���;�k�$���i��D9�yĚ������/����c��5Ҧ���F�C$�k�zѧ��#�5Sݪa;-��TK�WW�BmNt��e`�?����}����#e��5�p/Xsh���O��V�[���s���Pcp�7��8��A���J��R�9�#���0�ۣ��s=��b�,��UTZ����@6|"_ ��'6$�mv�8��e�i�w5K��*B�f;�]��Y���@��[{�d�	B�V�%ڠ�U����m���^o-TNl���	@����p�V!̘W��5�i��d�?��A���}F)?2�bJ�:��[�2!\X�Nr��劉�n�`VO�*��/�U=Q,�C�J-č4����0|�OH�v{M��jh򆇎3�]�����ӻŇ��x0�pW!q�u|[w�a=X���+vS[9�Wž�xcjF���	�������а�Z�y�nEe�Mۙ���฾�O	q�ps��x�I�i�#�v^����M��U�E|��j�x�Q�����1���MI^K;;����z���4�Cr��މ��:��<qx��|�^(�Z�,;h�jĀ:u2���s8M��"s&L$r?KZ��:�Zak�ZQ�<~���s#S����'�"d��ޅ\î�;�!�롂��0Rf�x�Bf��_�c��D�vMFM����ťQ_����m*�7@9G��=��[
++:�v$�~�)�D�~�zim-�����M�Կ�yH�d���6���2S���uC"��5���*vξ=��G�N���&��T�\~��mI%���''gǭ�o�:ȳ"�ȷa�~���Ο-,�ޚ��pJG7��3���|Eo��6��g�<���2�M\^}�mx���<���<��ہ#0"W��v���{�Բ�V?��X#z?����Q<�*�C�^�}��͆(U:�k"�;Q��8g�>���Bo5<ΖL|3)j�r8���k���L�Sp��u���4�U?���. ���$�p�'��\��M_o�[G�ס~�F�!�8�o����{AX��b�|0�)�+PLq̘�ۄ� ��W�JC���P�.Nw��cÕ�[)R������#j3;��|�jHǪ��#}��_����_���p��� g���|�n_��q����X#1�U������;���u3$		��&u��.x�G���uQ���Q�M�j����D[X�����K�l��(�;�F�&)ɫCU�i���˫�6��j)Ш7��$Ie-fQ�<&��;�6n��佪�zM�Z��?4h�fB�{��z%f�Y���~�F[$���R^g�<>����|���-?�t�2�J���mJ����h�K&��J�|�0��b��7�y��k�`}1�f��N�6\��!,Ck��ŭ�H�t�T��<���=m���:;�>Q�D~9�]�0&+���3������;�ڷ��փ޲�İc�G�)�WA�����+c3��p��2�GnoJu/�>�s
x�ђ��iwἰRV��D���p�p���D�/�\��:�&y}�y�c �1�c��%s�uثХj� �E�E\2k��]qܓ;�TU��/������;��i��E�6�/�-y��ɵn�B��wy��?��� ,�He�ٝw\�ϩ���z�g9X�&���\��uKUYb�ǯ|v��1�57�o�;2r���M��t��ޑ���K�nN,n���~Jva�ټ'~��C���(J�H`�L�}�tL�:��!�k|I�Oj�j-a���`Õ9����4^��3|3&��j���0='�ѥ-�y��(��ZH
���4��?=�g�ũ�/�.a���5.�@,I�"q��((#^W݃��y�/�4�@|0��(t�m����{f��e�%6``؀k��u�R3�N5`x��\|d�8�]�C"�K�u��؉T���ݎ��{aϘ6`r��W��$�F�Ϋ����'i0K=��A8e�^J�H""V��1��2�/R H�Q�YWO<>Z�d7`��_�
�yƃʗ�DV~
-W+9r�C�0=��[����tf�>j���q:A�]r��{���������3�����Ȓ0���j<~�v=O�z�3{��x�����{�`I���M�Zu�+"7_�����>9��~�`s�d���_�������죝�D�qII�]
�?Q�n��,��KG����.[����?�i��oT�:�+��-w؟��"�ȡ�{?�]������v}��zDҡ������~t�'g�P�k{m���#'M���k���4$
��å�>)���q2`g�/	��o!�.���Ve��0���Ua�`�	�Q�IC��s��)�UĐx��"y�Q�(O3!h���ȿ%Oh×�?�����T8�����'�-�$������9��V'Hr��������[�ј�j���� jj�#V������<)ZP��m3��9���8����qi�)��1�����s���w�X�͆�[α|���N��>0�+����m^���cՐ�"rg�;��6�'�~�P<�����O�.Ь�Cӹ�"��^f�>J6����;�É!'o��~OdaU�@n�����(GXq��Me��&x|9��Xw��N�~���?�G.�,�z�et����*��sP��tk�W�xǠ���s��ږ�8�ZE�&�s-�3�up�Y�?��63�p�ٞA{K_�_�@�w�lNMi���=y|�]��=q���W���{�E|/������j\�+�͏�l��׍j�&;�/�)�ڪ��'��,z>H,V����Ik�����-��OWp=�36%T"�[V�h*�l��8�D�R{��ÜM�@mTc|�c�D��{8�w���t3G�
�f�A}��?�<\���$��������]��i�P�c�$��_��O����j8٪1�^|o���)� U���^��7.R��>4������f�X�������T�-��Z�'�&1��;���ɘSN�x�W]���>��;��z�a�_6.8���>�:���a����d��OW�6=��3��
e�D�K]��������98 m@hb �x��Ѻ�u3l�ְk�/# % ��U������Ӓj�Ǽ�4"w��@�N�����XuU��a���F�:�#�au#���Ou��K<Y�?���5�|H5ݰo��N}wK�U��L����B�t��Ɂ����j�����p�P��A���P)���'eB�[����O>5���QI��>���5�o��x_+C�pB[y��/��Oϰ�52�,�7E㼞��%�����^��;iݕ�(�+�H�w�T���K6m����UTlyM'�p	�+$3ݘQ�}���\���ږn.��y�ʈ���g�w�f�N: 9p%�f�3�,>�~���y�1�Ș��D4�'�ߴ����_��-�`�8���p����:�H��gI	��GO��H%
 Qw������n|�ӹ׊���L��Wr'���<�J"�d/`1�+a{�]/���B�)b���>#�k#�*Š36O���8T�n����e�����έ�(�W�S��5�mR��7t��x�� ���J�v��m҃�u�8U���wIGG�!��g�_Rx"�Oc�\X!�BE�f������F'��˩ec�@���a�ZL`����,���;��c�R9Y6j�ʾ޷����mR�������2�����RGL~�:������)ͤ��\5E��p!fR�I%�sNAv���Á�c�|#>��y��K%@T�!�\��>p?�\3���f���[,��������=�r�dn7�R��R(�O��EOl|X��ez|��Фwt��Q��ɽ@��8_l�u?�Bp�?+g����"7G  ���޹+4B�9��N�J0�j��W<�t"5�Zճ?F)ޏ�z��{���~����A)����J������b��\̈́	�4>�Ne�����	��|p�k��{'8ݵJ;^���j�:~�ȃ�23پ� �>����Z���-~>=Y܆����H;�����V[Y磌�iu����IIo>���=~E��(M���"���[�j$TkD�:lݠ��2��5s��X����苯(dz�OSYl��S�xV&��n�������;Ɣ5qh���<�nXײ��e}�pƉ�埔�c,Xv���ԗ~�%���)A)��U]�;)�5��σ�9e�[�T;�V��,
�A�nqi��CW^� �`vy���U���kw=�e=�m��G�lִ�B��n]�[G������{�aV�FM'���r�WWQ(���_m�����lPk����!���+����,����<��Uc�L`�1�����[��u�q"���_�ƈ��>�!鋆�+S}�=�"n��H��F��1�[��t�?p�Aٞ��Q���s��9�v�aR�6`.NY��Z�S^��U�8���hLby����d��bjQ�O>���45H��]O1(�mаZ!E�:t�18\��ؚ/��Qے�P�KEF�e{��}y�?�ȹ�su:7�>~�7�%���K�W��L��Ν��9>�8{gYe��ǔ�ؼ���W�۪!4�^�Eu�1�P�a�T�2�N7'���D{�S�J%߱�����P��6����\�(�+ݍ�S��7,�-�L�{�@Y��i��nk,��b�j&V�����[�V�{���|���[�����5w���=�
�` �h�(M����Q;Fu9�$!�҇�f)/�T�@�o��doǲ�8� XO4߇`H,l�a#}ױq�"e[�4�^"��b��]��a��M����)�T��iT�dK��?�;���8��};|HD=Y
HM�1=�7���f�b#%���i
�";�)+"�p�%� �gt�|2���Pdh^��ԁ��q�x�����,o�cm��S�XPc��F�}�~��/S�wҘ2��:�#�Mz���`�(�������,�q�������|����%Z�9��)��vq�K�����\/O����O}�_���M	$*���[����������?<���6�bŘ�A�eo�1"�+��Ēj��#��[�GQE�ͺ=�-@��o����~���;�LO�J�V����)wL�r�K`0�,rR�7s�ȳ;y�@G#!�l&��?�_B�1	-����-�q;�,��P��)�ii)E�-ڱT �p�O��o�U�Y�G��j�!��ڥ�;���Mzz�-��)�����*����|F�@g�����������RqR��ޤ����*���1�pE����9�� h��!x�G���K�p���}�|8�ۋ#䐦��G{����Y&�a<C�U�|�ð��b@��'�<�8�鲈e�v�VI��)��?�}�ks��m��bU���z�=Wm�Cj��u�5"�}�'�y�%��*	�'��p"O���}S�u?��Dƞ��d�3�H)%��B�Y)-�~�߻�/����W������_d���o\wptX�7�r���q73܂�h�};2�$eK|	��UuY��.�y���:������,�iqWxg�I��+V�����m�#1�x'���7�#�(�
j"q��V��нx÷�P��
��i���ix	�70:���'2�{�2h�&1�c�[�0�E`N&�6ְ�?j�앉��hxǈw�J$£���c'�m�>0iTgQ��%�Z�z7��T=:I?�����{uO�X�0za9��:�凿%��p�Ja>�#�I����8��n�6"n�����	vl���K5�*5ty/�-yrA�ܪ�Tc�[�#ñ�5��q��q��N��3��P �Y�F��+�z�Κg����3ˣ����K+&����S�s��ḣ��2�V%�IV|e� �l�s�ܻ�06y,�[��U0����Ыe��yE���Q�nJ�!��30x��u��.�����ީ��_�Z|���P�QQ��� � �R"�-�4J(J!�0tI*%%H���0�ЍHI�C��}~�^_���s���=j�5(��.������(\c5^SF&&w�*��"�/#�6�o����(��f�^�Չ�00v�lОE�}��a����������S���L��5zX��Г�^=�F�|l��+�#j�����$!b:2gџ;��P+�1�4{�%�mkrk�WF�iT�N�*��Nb�ٶs]�s�����cBX��_�}�xv��9�W8��Z\|��Ml8h��qϭ��{�l�팪2w�#�&�|񿞺�z؅�2�:|�?= >�D	uĠ:�8|t���7Ζ��Z2�ٶ���W�3 �۴V,HN�bw�����Z�P���	u;:�l�я/�7��!�h�a'u�'^#m��Gr����=Wj�.��s$3���L���eb����\���Se�h��Y�cO�1tl&�Yqr��^he���s!b�A /�N�)��e�5�>mk��$a�P}�ֲ��/drO�"T:�"����<c]4�?K99#ј�z�)c��hi,�ơ��-JN���R����q����(�1�8}�;Ъ3�O��\	Z#��1d�	e�s�ݪL��mݬ�m��^�	�#�,��1���+ ��!�5\n>곑��S�34i�.}�%�����콱w'8%W$łe�v�&t���7�3\��5�}aL�Ò�@I�!?�Yt(N�p޺,Wq�?���a�{Il�Q�]L�����>-���f�T�/;��u$3�)����~�k�=��pV�7Z9	�d�u���s�#[>!���P[�m=�r��F����T�S��ӶMW_ϙ��I��a|q��o�'�̹ٵ�I��4Q�;cJ��7k��u�B$�M*yV���U��U#�P�ϧ���L��.��pIi��C:��[~��9 ڇ��[���,��V�s����}��l��r�v����;�F�L�Ui���9L�Ϲ5#� ��8���~�����y�Sѿ$V߅��	�l�Mg��{`/š�A�rX�㮳��tx_�Z���R��'�~��l�S���TCk�_�)v����sĬ���E1��M��u��}������A�� ?����[Φ��Vͣ�oF��^����{�,5/;���x´f����O����o�X��*�O��g"QL�������gK����1<�ױ����s��I#�r���NOڈ�4��*�;1���@������l�%�{cm�4�<�<�}F�~}�� t�qQ�B���&&u5
1Û�X���ف���Q��PW��B��T�����#>��(�P["^:���1+�G�4�F�������&P�zQ/�p�=����M��;3���Vûi��:/�;���v����A�h��VKC�%�9J�C�V�����+sg��c;�/��#��{�A�Śih�]��-��o\C�����KN��'��F���?�����2�ly9\�������w�'���3�$o�f;@˭Em\>�]V=�﹵����A�;�b㓸m��ڲ�\d׆�S(��l^�yfo��7n	�8� ���
`ڗ��R����[Ӏ��*��ο	y(�ld�������N�Փ�/����{�>�8��^|8}$=�v�'�"�Mj�@��b,�EL�nI�Pi����x��On*fM~���(���Z����K�qv7��~ǹ;��gn|krU,�<�/�[�5o��;�O��}M"�Q���nw�a">���l��t�x�>�bC��G��Z�U�\��s�����k�����͜?��~�!��i��g>��K�r���:F&^�[B�2�7��54
�	�i����J	8�݆���d���*i'j$ĵeZO�Zj~	�{z6���a�	n�w���u��$��l����iJm���j�
��J�!ވ��i�I.�W�xw��`�{h��?4��v���YFz�M�W�F#�<�&�[�;,S�h�q���]�,s}��4����ߩ~M������'��7l~I{�3�
7ȭ�|�y'�7>a�n�fw���z�L8utB;c��C�$y��5����_����Ts�ZzcY�4{��L{�֘x�&Y�y&h�y���SO���GxV��MXp�B_޻^���C��r}.A&�#��|��Ŝ����rň#T����1��vP�By��$�O揠_�)��������M�_�?����1Y�Y��k����?r^����wOk�^���L�l񷩕r��9v_���`�&��a��`�e�x1#�Pt��ʽa�����8��.�x�����)�G�֣Tԡ-�� $듕Au|�� $^~��ȓ$����?������|/�Zb��(�-��"��9�&�	��'�c�_�h�	�f?�$)j@�pWV(B��F���
�Ю���x��n+GTRx6�5Ο2���3��~����}8T��2�u� "��}�}*A�A��,�}����g6#?��ha�{A�6�a��`5D��Zcy�?�M�f8}��4�ƴ�!a�EУ�2�,��s}�
Z#�`_��s`���w� �N��נs�vAZ~78_WE
�ˇ���_LF���A��cd_"��d���i���ﯳs��A�ɬˤ��=��#m�-vi�掎ͬ��a�ۭ��;����ļ_Cz���������V��7<���E��>����x_�ul�S���LR�K�ɶ!ݼ��㦲������̄��SÖ6>��9���T���[�gd��x�8�&�{��1<۹.y���RB6��c��$���y�p{�c�� B���S����a��UZ"�UdhەK{(yO��%�T/�^�b��v��{4����՞����+�t}^��
��K��oqlS7+7��"+b#*G.Xb�N����ݗ0�:(ט�P����{���6o���>lY�j�5iP��[�	���7��jܛu9kk�P#����z2"�l���������P���Q	yt:�����z-���	{T�-R���?�}��������'�YW���In,�`�z�����l~����������a6m/�����K�."�~�0.코d*�7�{�!ҷ8sL3���BD�&q42WR����
s��{�Y�~��ȲD),O���on��=vXeb���kI��|��e���D��ew�+���#�87"iz��l��\��K��SM��Dl��y�xySMT�uE�4�.�Ӭ�{Գi�ګ��Ɨ�Y��z^���j���y��� ���bs�0�"'-�S��3��ƨ�,��z���s������(�������Wҹ���5){O{����e��-�<���b�,��#���:�����.`y�����!�Ћ3U��z���(�Ь1ص�h%#`��d֍:�x�T�Q�T�����X�����[�I��B��.�f"͂g�FnL�D�m^D��wQ����+�d��-�hک�� �NK|�I~��p��:}W�$�nL �lY�.�i�lBL�<��a������Y��H�P����׾H��7I�塥��>홰��,z�W�hv�-����q-���8��g�9G��<�Jnu��s�t0�>S�"���f�R����3��8^���g��^���`e��p�#�L�Z�p�	��h��O�EW���^K9�R%�YUb�"�j���i�k})���x�2�>6Λ}y�� f]�y���	j��H��\��[�ְ��3�O��IδDc_��D��⾠�q����α ���\�����?"�a|B�Cl���Nv#�磣���k
��ѽq`����ƃ ���H��2ׇwpg(���_;������~K�nوt[}|+U	~r�b��SgfW[%��k�,�X0��gS�)����s�p�m�7�ĎBB"�z̭&��o,�x��pr��8���V��b�:R�N7>~5QjPv�p�j4d'�����F��&�뵦R��jBa4w�O����_R|�t��@P	M�0��>}]�E�up���м+k�3F�x@�>�:��w�*c��kQ��^�HX���rf�_D.D����c�t�%�c_I��!	:�Kd��R0̹+���\n�D�H�3�/�y9��%�軍�nw���l<�=��K����9R��G�s'o�M�zv��܅P��>�� ��a��_;9��[�5�����P����͞��Z
�M5`3��C ␻�͡�-5lK�ȋ�����ʼV���ȬT�/�q	m�0g~��g�z��&��=�E0�;G�^TM�y��!j�����+��u�f�n� �5M�F�N�.t-IC�̌�5ń)w��4o8�J�%$BiY�&��U�L6�N
�Xu2[�oB$�&GF������|[��a�/Q:��=� 
�`^G����0;���#]O9I
��Zԗ���P�?�U��7����w���0&''Q�v����\�0�v�H�a���wL\&�m(�K�5��ڹg��q��)��6���e%�B{���c2�[::���R�2�)8�f�>�a�_j���c��ٛ��l�[	1�?�,'�^�:�'�;��nR���ެo`���U�2���;z�]����=و[��R�P���m����(u��2���^�K�!D�6���Ez�����K�� A���QW���Nu�{�d��c�a�1}T���1��n�ʸ�E�D��l��w@�����0^T��/>�+�تƍ�aj7�r.!o��ۣ n���#�4��[�&b���gё�'��w�ܴ"�2�qk����	FH��wS \XRoo���ۍ��kq�'�>�e��G�o<�T ��,����vYa滋>�ׯy����h�&
@���$�����t=�a��JSB-��,�y�~@�_�ەD��|Az��x�e�nP#!�x���ԍ��O�ufA�Ɩ��p�*	�&畜6�N��i�Kj+���X�4���]�/>��o�M�xw���c痩&hX�����D�N7�l�G~f���2RFդ\�������:�ZY"
[KNҭ���§)o���"��M�/���@�Q0q��*��j�@x#�:F���B���X�t�H���_�W7-��HDF�10@� � �^%�=���'w%�D��\E�H=�`S��Y��~u1�;ܳ��t�	g��/E,n\�'
�^�6�Ab��`9V��&z���T]���v�Z.�g��G�|��q���Ty�:�i��*�-��f�G	����z��]|��8�
�w�M~چ��ۢ�S��ax~o�s ��#�)1
%��W��yu���vF�"k���b��F&��i������VmV����&��Q*�γ?g\�����y"���iˍ�l 鰰��<I #1� F�\�r7[:��+=5��%�E�)>������M�ZK�>��v��W�̼b�`jc�X�Q2�iߋQE��S�H�߾�a�3������z���՗f�_]g-Q�n �7f�ū�� ��M��DT� � <;��i&�
\��}ԭX7A3_��G��?ۀ+¹$�EHQk�%��L�kT��nB��9`A��c��'��7��Qؿhc����!�r�t
�8��Īy�� ��@8��<~�����/捒�j�#��6f��@�G�Y�%��4l0a�%�E@=+M����s#gI�B�[I�w�&�)�+�������[9�G!�-YU:_ŚwdP��C��T�
����y��'�z�>�Dě=���3S������C+���N0X+�Re��5yM8�d����+�4]]���z�f=0���x��̽���ϊ�~c�ӷt1o8��3�J�7�`iz]6K�C(��RjB�u��\@kߩp�<�"A�$��p�_VSBlX;E����a���o���� ��8�e;����ݕ��a��s'�B"�]�f�F��a��ܝZ�g�r���]�2"�.�RK�ɘ���&� r﷢�$\n\���p׷|KN����c#���%FY|���g|��@����#S]X���H�9븪��a�"��	�3�1��4��ɀ��z{��޷%Z���4���b:�PEϵ���aAy�X�w}K<$��A������R�;;sVXd�9�����>����8J]@�#9�-�^�Hr4|>���s�-�G�.>؊Dܳ����̱�z4��=P�Ǭ���q8s�Z��@�^���	j�F��~8d�4v��T���(ʯ��')�҂�~O�� 0���Yhw��/�Y�o�M��޴�Ąs�&X�ljF͎;�jvm�h�Gr�*:�o����E!�Q�ِn}:���%��O;wW��%�Q�
iי�c�&�s`Ȯ�n�����̫�&Ő��f�cii�A]e �v���nQj/_�6�2b���'�a�Sצ<�H��Q<C���;O:���p�mh���v���T���|M�����N쫞�}޸F�!��� D0�Y���7�ﭫgVU��ܥ�4��"j���,hj2sc�"���1����eQ�{�����Mi&���{��b��(kl� �zP	�d� �k�Y3�q�	�o,��N`�E
���1gy�2�?�!]��V� V�L�s�61�� z��80����0���:��7�D�cs{;��{{�,���� _~�Y+���?�����
�X{���w4��3��3��;}���Gh'��U1��@�-@ӗS�a��Z�^ޙ*7���u
����s������gt�uS[-}�����6��9	�^(Z�Qj�y��n�b�jfW>���p8Y��u�����L��ϵ���{��:���g	=��  ���=&�r��m����g�ǳ9#��$���}.�q�����8�d��ŸŬ�u����D�{��%����wHnH�������k��뵁��L{�����7�"�z���+��pu�C�dc�趄����£�$��A�!�I�~x�MӔ�ǉ�YK�Or���޹U��O�-k���:�ce�Q`���>`�
#��s�9g���,i���`x��簴�+��. �|�z�ǣ�O� ���� &���ݷZ3��	�>.$u �tgz���dg�m���sf���{�-��4��7�I�j�/�\��LUᛴ��ظ)���%�|:sMl�.�b==�����Tra"DڇL7���ۣ���bll|�gk8��r-`g��=��]e�:�����u�����iO�	���qjg}4Q{Y�̨tN�"}ǼT|Ǎ*�6��a�*
7�6�0j��E��d�q���c5�ќ��ȝt�����(�ܶ��	�!A�Iv��v�a9c/���(������n�(�&���b<2B\��^���=Ҍ��k������x� o����i @���$�� ��k ݤǮh�=8(����(�MN*��	��a�Y5��j�0uk��e��o(&�/rl�ȗ�x��/��Z�y'�g�.Rwdb!!�+�C!�γ�N�oH����1_�� p��/9~�Y��j��8N�����.�W�@c4ǻ+�N�m���`iCxǔ�n�{Ev�ۓ����� A����,�P-���x����Q�9�~�����\J=&a/����7ٺͦ�԰ %ſ�V@���Ҷr�l(_�M䨆R�=�~Ni���=��>�mYʚ8�s������2 dl5�N�4��/�r��)�P}c��C�����3�h�(����5��������4�x���pϿB����GJZ�j����%���/z�g�)z�Zs=SIy�	��[��s9e����2�Ł6P�+�ɦ�G:�|����{�s�_.:������?���=ʤ�P{�r\���h�Y��nre�������2,7��a�A#��K���xH�����Qg�݄�^a�#�Z|��֌5E�����A;F�H��wD�z+#�5B^�Χ�
���c��]��1��~����9�:e�CV�L[~�խF�aj�g��ck& ;Q��n�ӑի�Q�>�մ���2�O"�+��sX�<ｘjr��>��Jׄ�UX������\V���ˀ�]`���*����e�9H�0����?"��SHq,�ɧY��E>8_��z�'��]|����-]��K�H�h�'�0������<I�r���wԤ�glp�|w�pZ���ȧ��C��ݰ*Yi�n��<�i���E5S��L[?�Q����i;#�ϟ?];��d���𷷷�<��3����)��$��a��Ȧ��]-ф���U}Ҁ
[ۿ5�S9rp����z0�Y�Ko�!��ԬS{U�y����$�3"+Z�os�N`�A�$�ҷq�|w����L���Y��^踽AZk����\Tdd�ǆ6���W�X��w@q�/5s��Or�ij�&[UbU���N�SƖBW	m@7�|�Sl�)�����ᛊˤ�}���Y2�[�YrM�$kq�� }����l�x <F���>a�w�����; **���OR
��<F��z'�]��R�e��V��G�
Tb�r><���ZI���'22�*-9-R���k*㻴���hBm��I]��� Z��|z�<�@Xȹ�'�.
�/�jG�c���,Z��D�ƼW�-�H�.�wjYx�m8t5�Wx��b��f�@{mwAY^S� ��:�ah�^���i�ݢ��r>�Pi4 �)�c�khT"�\�q�����hGO�v��Kǅ`|����H��hn=�"��/	���"t�fڱ%�Q��|�9~̳ܵ�� ��8BxO/�b����[*d]��ŜkQ�񰴞�!4��ss�ewj4u��u���h��{Vwe�$�9�E�X���>�9���{�U�hC'�R�����q�����6������{â��}�.�P1a�ȳⰳV�x��Y�H�;���|L3�����y?�W h�'������nf�uML����Ff��p{����P����ř<��FV�C��ca'�&(����p�ɬ�s��7�ϑ�8�!�ok�LoKP򽿪q\Oz�C�:���t�@��?]Ƹn~|s�˻��i�Ա���.`I�z���	���]G\�|�8q�����B,r������Gu��B��15�dt�K�|@��Y޸�P�d�c���,�����VRڿM�a'�y��n go���>���(3}��A�-M��#� �k�!S��U��r)��R�\���ISi���%���Y��@(FY�rV\���1�$�ت��(��y��霢�����v5�#2��~��M�B�~�q���4�F�,��� �9�����'~�x'8�Q��:��sV���TJS��v�p�sUd;����޼R	؝N!�Z��G��*ρ57��u���Kž���C"�3m*�Wh-�H=������\J�Y署�"��3a�x�I�h8h�7Α%��p3����[��t � 9f1�ٔ!�g�vvܨ;3(©��f.�+M��~3غ���1񖸻{��j��|�%��NoG���M�b�c��%�?�9a�A;�PXaC��
��.�p�_�
B��M�Y�Q�1�-����AGIEK����r� l���&^����B`��05���.g8T��l����j�ȉa�?10��@~�q�x���C��5�Q���O�ݦ.IA�IȽ���|.����0ʷ����h��U��������	���gѮgי�Y���KB�W��[��&�]4Z��4����(�B��^��w�!XR��������p��n7y3��m`������IZ�OШM}XPc^Q�GHB2��]�i�^�3$fz�"�˟PK��a��[��e��ȕ�kԁqQ{'���`�Uy����h~\���G�!U�UV�$轴 P�{�T�>�ٟ#:a>��F��:,{�f.�|��l�a�L�g��z�F~0b���얆�8{h���q��L$F��22�������2G7~��,��:-E�vJ<:�s�C�>b���j��j����+������z��m��T!9��Ea`��7�yZ���DU~����o�Ht�������]�������"w-x���̺��ʶ[�� �ӌ5�\0���	��/!����_&"�q}(0�,5���_���	�q����H�����3���XX���ĺ�Ԏ�ʄ��S֔�;��A�3���>!��djEF��/���@�1�#�o�dZ�k��]g��p�[wh�ZJ�] l���^�P�E�9L�H�Ѻ�ސW�P���[3�^�s�������c�|���-���1���0��'蘮ʝ[׻b�>zm� h>�V^��a�J�^���:�s��[�įu�,�'e��f�a���9ˆ��q]�,i�M�@�8R!wn����l�ov�;��z��TX��A�
F$���3��T			� � ��c��1���j��T���ü�K������up���CJ~/)�V���(��/��)$����}PV��S��s�>a/���g�ȅp*��oj k!���/��w���j_�n+��=7ί��%m[L @�����k�v?�aK�=�����N�ؠ�����v+~�
�3kk��ʾxFiR\�љ����~�}:?#&xC4���%��
J49M���xƂ��U5��:�0��K�>�f�j���5P#Ǎ���!�<!�mt��C�̇z�U��K#7^^Y�Z3���\<<�&�gF��bmr|U��?k�=0 ��&ۋjXr���Guu�*���q�??Ҙ����wl���e#��*RL���C����0���h.6�0�����@4���[�h�02�g��"�X]g�Q ���l̘:q�&B έQ�_����/ӂߏ��j�	 +d��lw��
�߯��9�7���n��u��k�?:>Q��7�0'��:�u��$y*P����n����C����g��a�<!��4�a`�2ԮDW-�'���~���t�|��;@�Y �ִa[�����Yom:˘)+
F�S�90��e[���F��b�e�6d���@>�G�e�bW��;��4��`��a���̯� �0'�l9��/ĹJ<��fYf�w�!u��μ��
n��`�~��l[����ՌG�!-?`�Q�>?�;.:�$�+98��]���vQ�3��T�z߷.����N��OTSْ�'�mj�?��9[F����C/����!	g�����ub(l�70 !�����g�����cD���m1.)�cM�������JJ�.�Q,Z��li�#�Q2���ђ�>ƭE̮z�{����VG�f�����V��x�l����Ą.}�!��-����VsX�}4�W�w���5A��c���f��hGƇ��}5 {�<�yC�̀�9=�!�`:`��sKj51�8��l�~�h�=Z��xX� Cͮ�i� ���n�4x2��"��-nd�Y.F�S���e{���?j�\�B�c�E,Lt��X�0R�J�����.�!=�|�R�`���9��Ġ�1W�+e�"�\��ȏ+|ځU�����)%w6�i"��������{l�z����}Ԧ�$K'��qx������̣�cz��(&?�����g�֘���Y/����rI���g�f��Rj(".�z��%�s� 2*
P:/��@��=3����(@@�l%'|	\�n�@P�Ls�nK�z�yۭd�i����v��t�[|�橛x��n�v�wX� 	�TKu��4���v�..}��}n@VȒ��/z�&���Uv��Ӗ�EZ�`]L�t�]�P�>����Մ���w�H�4�$�!���Q��j��c�ȵ��R�9�B�2�����%*
*v�%*O�=M���b7��k�}�2�3d (���n�3��m���v�b`a����my{�d&-Dؑ�>3��91�!��Î^���?%1��ALgko߹���d��km-��Ty���N5�D��4>?KQ)-]�\�~��_el�~MϺ�1�� x�vBO0xem Y���!�:<.��X*�c~K8LW�4y�T����:+�;Z��Amو�MiRI��߆�k*yټ;��e�0�1R.|Y����[�p������Q�YU{�'��6�Oϔ���1r�����NGz-wF�l�;�:o��� ~�MQ����7����?ޔ�n���X�/ފ��NS��b f#;;{s{[QM�
���`���C:~Y�r��>�&힟&4B�Wq�Mu�-�˭��n|j
��R��!���h&%�k���~`+�e��n��]ޓ,�٘ʸ~J�!&�h��|{	򿻸�<ۀ�o�՜w�.#ro� ���rFF�M�{��7��y���vd~��|�����"����:�"⟹v��	Jt�����B\	��07_:���P���ca f��g~��'�G6��kj����<�����v����j��$v��s�I���@U뮯#�?:��CF�#S%�טO��������q�c�L�Mo,��V͏�V$���za��/9��
4�6�/z?w�Ċ�v���h�Y�2�O������,U55A99����";HB9�ϭ����2`�l�
�����Mc��%���y�w�okk��D��(9Z��Z*=##N(ţEv���?`JPv���'�f��-HʧO���sXo��]�z F ����T�уl2��Bw�3Z�����I=s�H�Є�����"��J������Q?�d���G�!�U�Ѫ��"���B��&9M__I
 �(= }��-�)�{����.ˉjL�&���{�(}��	H��&O���!VR\TQ��bi��g������R�^7߳�1|rX���uf���gxQ�8�-y�8���.�xF& #sX��z�Zp��t3R���n���ˆ�:*<0�h�@�{�V�\ ~���SB���&b�?�W��3�贐���Eǝ��M���n���9�1`�m���qt�n�3��'+]��y\�	<%��7?���z����*��@ش�Y��{��*"�15�o/���X����q=8�x�탨�ܖ��kd,?�1V;�Lw�P�X�V��%�}'DQ��v3��E���A�P '+k�f�@.�w�bo�m	����t�!��-�9�iq8tu�	L��8v������*�׃%Ա�v�^�w.>��k	>�PJj*
}Ξ!u������S��ӡ�m��^�13w+�(�
LJ4�>�	���������f�\>l�szv����//ޛUl"6
- �[�*v�U�i��z;���j}[z9��yʇ����d?�)dlL�z	G>����qſ�:��WZZ �8�iUE::I`Y��	Ø��R�A�旅��υj%���{^�@�7θ�w��:�8��#��oO�r6!�~?o��/���U7%,0��ծ@��ݓ����Ɗ����kh!����<-����`L-��
\d5}0<b"������NQcx+��� ��.��s�	��v�-�^�������R��}�z�ñ��Hb�gX�ueea�z��3ҁ�:�)��p�ߟ�k17x��#��l�M�3NW�d.�!�K��Ӈ�󀠛=�q�镯�����J���n}M�r�曱��:�h=�L��8K���`ߌM./�� �m{�\�,�c<��be�y�r�C��)&�Y�����ʼ��6����O��+6� �w���t6��Nϖ\V@�zѵ�R���p�
���= ]`�DH���6���Ug��t�-�*G�2����l	���|�[�m�7��y`�]�fl�=9��/�'����e�/aiD�eDǝ��M����<J�5�O���+����Q�d=���� �r�t�L��H�ï�ľgVY�|�c��D̥�l"��!��/ pn
��-HU��gԳ�~������8U"Q 2�׏��Fo���i����� ƭkcu��7��B� 2�+��g�QFei�����T�j�%�����4E���c�t�RV�������Ys��ÿ13�8���p��;�	�W���/�S\��R'�C&�����9�3�i�gg�Zb��2�#����2��)�T[[���N�f�/:�Ќ?�� ��b�����*��1�v�(��]����<
(��Su�B���ؿ�����]�����#[��Q+��?/��O�ڒ+tGe�!�y�0���gX��20y7�|hHNE�u��Vr�/2�&���n1I�K���F�g����"w�ܜN[�%r�K��vF���+9���+�����DC����w��=>�,����ʪ�k���q;�[�2^J�*A?|��S�����p��,>A3��o��IJ/C�;��D��ٟ#��@�.p$B�!���l�pש��t8���kM�]��a7y͠�����V''' we�:X�)��Q�n��2�Qds���.٤1f8<T�<�c���`�
]9��J6�##���o�.���lcNT|���&oGϞ0�z6	�]�*q#y[~�C�l�HD���}���DRNߧ���
��|������������
�nE��@�����U\��*��sL>V�q�^Q��B��s����4�غu+)E�x?œe
-�Y"J�}㦦�<���yï�܊bsL�Ē1�H䁜;��'nSؼ\�;���Dp�����{5����Q�����7*�N��Ɋ9�6�ea�m)K���Օt�pN�^�*m���P�0��'ŀ�j�NSJ1��}��1��y��
�a'��u���V8��{^G�^7�����P�ii����8�$�ɵ�9�[��h���s$5�A�"W>�g��?׸p�³خ�pq(���U��\D�I:=:�8N��?�z_&@ajk�]�B�q��|Kjii	H-^C���J`��\��ѿ��1���A���>��6��=&���n�����M{�j���\��A����.g�e3�I���/q���a��aq�7��Րϛ�/�#
���[h^�`9G��;���!	��s�gE�r�\/ (/S�j��5�,�����ߛA�}�$�z1�0))����
�4J�fB,���Y�?��&�d�E��<�ш���\���.y���`j���"�NU4G��
[4�tD<m�A%����QR��3�8���|��3Ab<s�:{������pZH�#�ٻ4�
%x��tȟ���3����o�(n����oPy�����e|H3�]TRwݣ���}WT�UW�����X��G���~����I��KX�)�#�I���{�}e��SF�����E�?��1M��^�1:�3텑���<}��9�/ƅ�yY��}�
<���o7�vE�!�A���5F҉���%N�K<bf��P���N�;0���*�wۘ�^S�.�妙4ʗ�.m��:<rt	��Jg�I���>��,�d������\%i_=��� ���4�y��3�����|���x/���h�-�I� !������S톁-@�GG �z���s��B^��u��z�;WgA�=io'�<	�k��ГAȑ�[�B30�3ꀩ2o��pIaFE�����壩�� !����0u|t'z��,���xM���"�|�)�����=*6�:&f�G��m�_�.g���H�n�m&��&�lV~�!������=%���s*"x��2��ߘ�+<����c���e������Y�rߏރlLDk�ࠋdu�#�F�.�x�vʽ|����A5���M[�4>=N6��@Q�� 韲a%Gg(�C�p�I}r3�q�^L�iǲHMH��m �{|O]��y&/nt����˜,]�'	��8��vj�����cofNf��%s�"��n����.=_usb�{�h����6G/�q�.����RzL��m�Qd糙u0,�(*=@�fZ=�k��v����^�s��>�'��#���d�Tj��<]��:����N3S��uŔ�/ßLv~[z�e�Y�T��^v����Է>�<�<���U������;���Q�{}�� q�!=i�jUp���������hh/�WG�|]_��`�J̚�C�o���ҒxQ��3��V`��C1P컑�	e(h��W��}t!K^rX7�U�&Q[*�->W�g�@D�&�{o.�������
�3j'�#��yqjm�g���SW	#:��Ej4���3X�=��w;kb����2�MJ�߭���}#�H}��iY4�bz�7:y�Iʰ��H���ёp���|lb�!4�q�[AnKwO�#A�V�
�<KJYF׋���Օ��@��ä���)����#d٬I��ԨA�jXtv1���L9�(�������O�c(w�6dF�+)�h�����u\7g�^.�)E��y�N�K�V���/<��Ǿ�W��(Qz�����;�(ʻ��8m2I�\(�<�:c~@8�w
r7���o+�_ׯ s�8�ҏg�O�u�4Üמ�z)�CR/����s�	��dk��a]�����+湳�܆�Y���$�h澩��4�ݬ8���nҜ��>=u!,��Bn#�3�s(�~t<4Y5�.^�uv"W(�cֻޅSآ�~���{����X� �eח`n����*\�É$PouP��c��?��n|����@����Q�.b��}���r���|��Q�����0����a��2���M3k��wE0V��G���	�b�lS���b��&���TI .Q9�������J0�Qw��&^�/C���Ĉg��",�� ���2W���`�U�>땻����,���%�����|}d��� ��?}�Je�)<R�R�Xt�0�x�)	��(e�^=��� �p?������-J|L��Q%F���?�'І��������'���E�����*h�s�]ٙ��� f=®�q�8j� =0w�[��ӨB��H�C}�	��љ��~���|%>�<��Q���������k�;���n�HiҤ)H���&�w%4A@�� 
R�&��� ��Ih�BI(A�=����˛�a�F��{�9�\�����ۿ��<K���ht.����"	QN�*��p��)�����՗R�ݽ�$}���/�u�f<�����c*4(��4�6@�`<##E�{08�Ϯ�$r�Y��Uc���;�l�'����%���_��^큳��v]��n���g�Y�>էy�O�lSW��u[i�S�zJ؍l����p�l���g�޻�8s&�[����ZP�U���>�񪕭�#;9[T��d�h��Q�#;���`���>zT�W������������o;d�
aI(��(�6����U#30׏اo)ޛ>��;8zfs��"�nf4[��Eӽ�!�^��M5!讷��.�e�h���6}d����� �+ܷ����%���炣�WXnP���gJZso���}������η�����=�rk�������7�,Jݤ�ކJ/���������b�nBk?�X���o��j���}�{E˭�� �`ŋ|��F�2�u<��ci�-A�t3��4^O�Pؘ�;N�u� fbW]�S�V��8�6��|����+_���wmxO�}�2���>#���Cj�0��F3ڗ�;lV���:{�����\��R��X���3�<�uc�nX�)}V�
P'��՟��C�ZGa�:���瀑ac�sw�p��k+Ò��	5 �`G��T���K�����w�]�6�~��1򼆌\A�f���:��׮���
{c*�3`w�t��EbG�]E>�׉nN>�~ȕT���	�_v�zz�j�>c�*��+��Uv�r���C=�8��mb����6��+�74S8f�M
˻0��o�����O�)����ɤ��9��9�� z�l�����J�a�������}����K��a���x�7����)i������Wb�+��"?�"WR�14�G/y��~�D���	�l�D��O�*�D�������f)��w>��
 ��N�~��nc,������$�\��$�R�
ѷm2 ��h����y�Ω����W2���z��-�/{SQ���V�+~v�bշ�d��\^2U��JR����(���\Q>���T��X3���1p���aER��d���x�8x�=��A��J�R*3�7˻�ք���<_PO�sMX����X8#u1��������P��OA����͡򟋧x�%�ºOw� �Lqɩ|�1/��wT�uG�ֻT<��>�z2K������-��z_�pڔ��I�)?�E�C���'W˰����%�y��m"0 ��hg�N2�6d0�X�uU����<���2`�6<����16�F$#1�l�#�;�lI�h��źS���K��K��Ffg��S�; ��u��`4��N8j�<�i��C^�-�O�X�M�n�OA�2�\��x�a��-��L��L��zqV�xH�x_ ��@��W�^��'j�����g�r�m�bً��eڞg��H�D>��ޝ]9�zB�(y�5_1�I� ��r#�~��O�#ۃ��������T��zߛN;�˳����4�����C��CNO��`Yœ�ĥJ�$B�3[��\{�g��\����zE����6F1`5��4,Ai`�_�+�':���p������e��1����ѷ2���X܂��'���J+j���Ey��{��U6p�B���t���y�~\�\<pށS·��" �w`LޙM_�
���X�CEa�òp�c�[�xk��UP�>��qv�N/;��O;�!�L;%0ڑQMC_���J쏨K���ʹsڻ_)�]�ԥ�N���+�J �*�0�(K����L��#5%���V��L�jn�bއ�[�#��s��Zʾ�ʹ#;h�߿"}~pɪ��PhO�wP��s�I��UOk��.����V�zaQ4�iַ�&�٠�2��Y��7h~K�m��G����W?�g̈\��y��-ғ���؜���/_EMkc9t�Hi.@�7����+(rܬ�`�(�Au��R=�,r��ҤxX[����͞=��7��S�}���4�Ō׾d����ټ�y��� �Q}Z��=#���U������O���oayQy���dۢ�[~�q�=<�{y�0[�S���7B��!ݦ1�IbQ���p�&Q�}�0�9)ЈBa��� g��v6;��0���.ϰU���o��'?�/�?Q�8M۵���b�� 84��P�AIz�tj��f2�y<x'$ȱ���$u������_�3]|����f�ѭN<��xl�|�s�Uty�}?+��Pp�(dS�ЋM����^Rq騏K`�5dag��h�����c[�לa�Ls`�P�-��Ԯ���3r�@8�B���9����a���/�%�<aS�{'����P-�?�)(�L�)���̦��@+����g�	x�����T@n8m�����k���ƢΉ����:��&~�GA�KCd}ξ�i�{%T���e(EN�,z��}���&O߭J�?��O�4b,�������������7��p\�mmgƥ�s;����\�^���0�.`��z�x����_>oA��n`n.�t���y+l�kv�萫?+߼o��q��?�G��ƭ�GA�A��g�r&��?tƋ{��T%����߈)�ٮ�_L٨٠��Wy/�y��}�pPab%L!�Q��/U�n	f�}�5�q䟻��x�+�<�q;l b���`n��v��E�b⻏��t|b"���j�Lup֋>�s�N�Y�nЯ��i�.pL/�r�B6����2��@�c���.��E���,���������w.���z�{�,�Cҁ�FG�mUb%�O;>��kb �O��犹�`��BS�k���k�Q>�޲��9�j� �߶~�Ŕa������ƃ:U9=cɤ@uѤ�/�/k�����BHݵ���#TFs����=��������/�Bq���ӎ����Kh��/#b�����F��ſ��]ئ���}����uf���%�˄�i���n���-�'�(�R���7��NO�e���b��rZ�	��[=~�_�I ���Z�QWx��ٳ�z=��|넘��R�t��4d%gw�"> �ʹ@�9�+"�z�C��7�@�ˉ�*ǀ��WTQ��Z���ѯ��5��zZ2�E7��[�}����-U;��'D�&hd�KL�˳[2q���1��|B��0�|���#�Ώ�2��JG�r[^;�怡���S�ҕ�#}R3�q�	��Z��ª����n���ɍ��d�PV��t����6:��z�d�m=�%���y3��X
��z�P/��51Y���b\||�p��P�$��
�j��7��^^c{�u��u�ן�U��d����yDC�#?B��X�8���!y�L��$�ρ���s�3x�d����?}=Uz�,P�\��#
'���fl�ή[���{��޴T�O5�sr�@y�;!�����s���@O~U��� �8���{���=/�H�RÈ����8���IYe_�aT��cFe��T��ߊ��A��~X�����#�*��).�c��JFl���2O�\m�ؼ1}☦�t�~$+����8m��?/J���1�%�p1�Q�E�Y��~�Hv�L��囓������p������ʃ�[*�5
�Ъ����pO�������Á�K���>����o�
i��覉UO�3ԸH�_[s"�D���wqw�tM/��鷃, o���@ؽ��XZ3�A�U(v�y-�n�pTOg�U�����o����w;���jE@�!��U���#!?o[R���m���W���^
+�*VQ�H*���T�zl�����R�Q'��nE�(�ϩv���>������<�	y��Q���r��pta1�?/K��j/d�]��S����YzF���ě�ra&҅�5����8G
�׮���خ��>k|�;,�u�u3Smm��)�:C��7�fX��Eg�.�4`r�<-9�~�L0�my�z&����K�M	�n��&�#��G�Zp[.`�ڌ��|��2����_�Ug�/:}/d20� �i�P�M��"�$O��(~��
�~|/,$���"l����6Jm���!�X�Y��^ ����]\]��������{�	[卍���*�~�~�2�u�J�ejZ� 6���JPȲ�s�r�]*�3+�J=�q�ڎ�0�K�Yuh'~�F^��}Fɪ8^)
^��o�a�^U��;|`��6�������V����:|;F�v�
�V���z��a�i��P�v���fc�*eea�'�@�ח���O�?�pO�~v/@���K�;~T9	{~^��NLL��Ɩj)���j�h�%=��U��𐰅�9��b�g{��Y�:D2��
9�~a��k	��p�X���g��+��oVɴ�=0��qP.E�ĥ�l�%v+��_Y����������j�=��;����6|������"
��\��o߮�>ZDJ�Vb)���p\)>`����d�r���CӢ������]�t������s��y1�'����Os�ӵ�m%F�!�}⯿2�6a�up���Q�:�Ϊ:M�f�iI�d;��lX%%�-ۄ�F�(��?��{�/J����b$A��Wb��@��E�fHx���eѫ��Z���U��B�ߓXo�e���V,)�d���q�G�����2�fdʚ�"R�HǶ*��x"�%N3*���>  A����}R2�0��~��Ù��s�r񻘬�N��2z5�t�ׄ�'i����N�Ҡ�SWS�>@��φ�_�5�	{"��E��b"�i|�Mu�`�C|����s�W��O�j�	�q��ƭ�ǀ��#�w�)�r�F���)���-���k�X����Ё\�O .&;�]a�^��3f�#x/�7.�<��0x��e���2Z�х��b��.�Q�K���XWOT�9]4�JI�����U�$u�#n`���w`j���y�vx5+��ߴ���(Q�"Rc��ܐ���Ί�=�\z�&�J���6K� �f���1�斣<��W���;�A	�>�p���*qCr��IP�6c�u�fլ����ũP=(��я�{�7�QQdȌ�Tcܕ}��~���85���Fأ����	�f=���$�H�-������n�Z��!�C�����{�|QO]����/�H�����ϾT�_d���-	�=���q@>r��m2�e�Ѹ>�JSx�mKES|'�HM>������)����g���`��-f���:tD�_lCq����1�эzP�@��gkgl#������
ߪ�/���b0�uj�����H�C᫸+Z���o: iJ9���HʓjF��DR���Oڻ��hC�\U�g��$��s�H+�\+��j�I�[���>�]8t�]��_2n��X���,:��-Y,�_�r���1�C���r��{G/+�u�p���O$7�����&%r���;��&�~��/E�\E�F���y��Y�t������lve�z��k��"^�zT�5_��N�xXW�ib��]�H1p���|�s`�O��1�-�Xxs���8܂�Ȍ��O�Zƍ��5�J:"\���ߤMW�.H1Wq*�cp$eV�U�+Eè�T�os��h����eq����O�fm����s��M�2��������d҅u�gjs�T���t���{�����m2�J[�	9*+�s#��F�,���b<L��CQvC�J�k E��le���۠�m��T�<��:ܨڶ�g�a�ߣ����< ���L���D�}z���������#6�S+[ނ�� ��Z��Na�9�����vp�\*[]L�A�6�BD�^���Qўch1��t}����\&���5a�od�9�G�'&T��Î<G�e�@_��&*B��n�
s�z�.��n~�Ӓ?�1F�q����-p74�n���:3�mz�#��[g�?h�b��\�$l�*q����¹�����ء&A��$�iE)u�����k�7Nῆ{�Eu*sf���F�iO!<Dd\�Y�$��P��n!d�u�WkI+rtl�㠄���������Ϳ�39���c��=�þ��\��	�l��]x=���-ʑ��
W�,;��Y|zRx�sy�;6tug,�p����k��~rT�>L�i�� G}��S2��3�C�Z�}��*B^o�糮3�>��/1�x�c��c�C=����$�� >rJ���|��B�y��ؓe���6��6��D�?{>�<��`I�ٙ8?%˟��ė�/rT�i�r�BG����*�q��2N��;[�a�߈V����̓�k+��1Qy��_�	�ȥ# �räʖ$+�2"{�7�bE�*�����k<��f~_�8
;E��v��5�^.H��t&P�i��\�Ou��ؓޔ����Y��lz˺��a��`c���.,��SK{c!R(��뒸.m�����D����s;���I�$2��e�Ӡ�úӘ��V�m�#.Ц�7`� �E�����>"�a�pP��#BPb!	�:}~��"�r4��*�ĉ To�ՙ�h�hrD`��MJ!'����5a�p9����sKTX���>;�ep�FϮ�1mt»#ۊ��5�5�25���m�Q�#W�b ����lo�?�ܶW@5�� �O�٩���|o_�&��^T�2���dU&��r��.|�%<h9��'͂��IV��f���z`�`9��&�l�ÝꙌ�f��&���i#�Ĥ�횓3�v�}&P��u@7����"��(��.����O`n�N�[�u���Į����0�1���!-.oN�D�Iw�s����gҊ7'}h�^�=�V&�F�[�u�~�_�|��@e-3�0�(x��]ce����P9w><����8�Y�����nt�����,b+�Q�8OgeB��������3��aZ+��=C�R�zۻ���b�>A$��c����#�O-�ñ�p�\S��u̅4o	�~mִџ���G%o��'hC��)�p���`X{H@9�k�D��������!�/��[9��(���Ї�z��`޽ۣN*!�磯���0�i^��#��p�(���W�_�U�}�l����u7�+�0����wu �7Y:��C�[' nA��pWݱ�2rpڗdr�o��!��6e#  �Z��z/��{��)�{�j��p�'���~�;�ၮ��;����b7�D����1��=ٞ(�P9�P#�\���J���5��_P�q��ν2%�1��+Po������0�x�	m��z�I*=
����3��7�y�I�|Q����X���ν6�D��)�uI-B�A�fu9s;GnIs�C':X'��@G�z#�E�ŻQ9f�j��&-#��LR�8�y
��2�j��I��#��4% T�nG'az�O}~�@�����GO���-�`��3Vv�磗��'��[��bʑ,e�Q[�A�3V�Nv���}���(�!�_	KоF�q@p��ȼ�S��m�%2LeK�������9������s�m�����M�|��(p�NG9~�[�dI�����4���3���#G@x��1����������4޵���C]�x����Ɠ��!Q!����$J$?VB�]��'D�j��;~'�xa2܇���бpQ:E�#��J;�����ȼuʙ	2��~Z���ݓ��̱��5��cIp�PNп��v29��o;���p�_l;(�LC�b���#� H�Z�ke�=Ѩ� �~ӿ3i��a�p�1�sӭg���=4�O���e�~:��ީE�������W�rX�G��|/�,gi��G^�[���H�3u;4���>�q���	�	�J��|���j�:��e
Yawm_&6�ǂ��u�����kD׹��G�\���`��eF#۲���J1��FG��/��v��.v�	��z��H�_�b��_���T~X��e�����*��&� ��m��[Q�4RG=�ܾ^?/P�l*p^���A�v�J�~�߅��^+|��[h?^'$�SJG(*3�k0�K��_�������󌽆b���XU�`�VL��%"����G�
`s���f�>.,(���sO���҄$ �`�b���S3�Yn!t{�|��dUs7_Ʒ]��Z�R)�r�np6f�&���*�&"31��f� �����#�\C���R�� t�@L[k�:Z�l���:����fΘ�	=O�Xr/�&�vE�����/nG(������
����e�����9�æ�٥���e_9��Kpŷ����w\�*t��_��"��e�[��N�1���h�//�.�O3�!���=�݇x.���儜L�H����[v���.�a�y�����G�'c �j�3G�t���r®7�3R]�P+�m�ܰ�����8�@��Zt���i��o=,O8��҆mZI��Uo����$�����:��|�\.;߀�(�@-��"����Կ�Л���Ϧ��Q:����ޏ�P�C����m�5�I�`ۑy���`հ���w5�Z~ƍBӇ�<j����]	G�Z�cD e���3�eb��=(���F��zj�"���w�&pI
�J-���[�q6oi"��U�`�i��ӱՇ��FB�K���Zܜs�Iћsc���U�`��'D H	�kΎ�$�i��#�$��B�4��=OT�
$��a,���i_���JVxh���'�������=�����IT��\57N��
D@��=�#�Q�UU�v׎�?V�.33�i}��gC�������n��q�?��a�qj���I��#�b�ښ�X�[UT�A�Xd���`����-�~��O��$�Zb|��9(\�p���s�16�����4�{X�g�я����D�%pe��,���w�;�K��H뢁?PBNB�Ph��y�+�޲Ӄ`�-�B��r���M�+c�Sr��N3���EK�!>�}}"�l q �+N�sJ_O釳��Q×��
^�DP���p+.���)k�HHO��!j?�IvUC�K8�t߿
�v�M����#:�}	�?�@q�3��9�[����֙@�!�U�r~>Ȓ%��'��G��FK��出�:�E��g�a�.�m�p(B���z3�U\ѹ*g�0ɛ crT��׈���G�$8O^���T���>9	��pa9�j�<��'�`s\�|���)�Nߓ/GO)e��L)����1A�h�h�S��fbv��5���0'|��ݔ�"U?s5�=L����}r�a�}A���S�v�H{F�Q��ř��O�"$�,[Sx���������]��JK�k����d9�p�h(��fn��A��Ĭ��0��⢜��-f��d]ϒъ�&��@�s� �����U��
�p"
8Ucg$��@�j<�	�&�Ɔwn���Fjp�5ֺ��s*҂�@/�_˃@̏�Ӷ���	���5��8�?w��|�z��.-�:�d7<��Mϙ������C�F��(��ef"��	)�$����e�Bh:�?��c�l�B[F&�
	�mW�2Q�|��[_>��-m�]�)Z�8W��z����yu_�84~:�d��T�� {������4Z�%@�D��x���>P_����J��D�V��c��3�@�W�n�S~T���6	�o�|`�x�/�0�GRo�ձH�q��?\�"n1䝜�_��g�9�;���@�I��� h.C�3�|�!b����&�������m�$B����>k-@��V��n)l�u�����^'*$Z���Z����a*-j�޶�([gM�3-	R ��bB�L�I�lB-<�m_0A~�.�P��!�(���~�gfˏ�7��n��j��?��Nd�'�*&��A'���DpC2���,�/s�a�v<a/�WmNhϗf�*C�0F;���O�`"?��9s��.%)Y�yX��x�5�r�����!A껻�����Lo�j���(	 ��v-�����dL�F�^�rjO}�;&����j{3�z������Qh�=i��*���f|@��$q�]�/�L:^��F�k��i��=���>���U�P�)>���9vi�>���Tbz���R/�`s�Oq0#cnۣ�!鿇�6��OWk�휂C9��*���Rw ��7��6g]Ź�9P*���C��$�_�T����ɒP��ż=��wͷfB��y�����!�/��yd�6�� G8� H�:��lM�~���=a.�4��@C��_�m���N/;��%�w����aa�ax��������q���0�)�"
_�g��G*�&9-8:�]%��-��A��?��n�=����0�8��S� &V��]�TZ8�la�=}���}���X|�$ՑK>��6v���_���3��]V�ҝ�n���F@�7o��;}΃�]��M�-T����?/����T����n�Yo%Z.X�O����Z2gcj���i�A�q;T �J��� ���Z�C�&<ƼkTG�K>��g�>%mO�ʏ���0Ki�2_�^�2t2� D�a&r���ڞ�R���Gf�s�4�H}c��"�6�=ˡ�Bc�j�L�� ��V���3���^���_?����!/O�`��M��,+A�PU���2����ȏK�Y��~�[�/��sU�o�U���K@6k9̟$G���9Z�ԓN�j���.���ٺdDwW�xS�@:�д̍0m�4��/������\�|P�k�C�,����uo�呿�P"-P2��"����$1��G�倦;���*�iH�pzjF �3W���3���7Y�#K������i�lOЀ@Fd������|��]����v/VC)6hY���I<57������mqㄞ({9��tPn���u�������V@��r���=uG2e�_�u ���=��E�*�K���!V���ݽ���]j��^|DC���\����O��+.��t�"���u�?�����mxK�v��!卂�Hh���C�����_K����7�=6^�ݿSU;��� |6�\k�;�Qfx�_Տ*��z��;���Jh�<'�
G��ٕ	.�Klβ\�c����iw���Rr9�ٓ��1��lA�B�6�b��+S�j�B�eS^��/|�X>τ�>�9��+��5��y���l��$J�էy�\Ϩ�9%�
�n�gA������>-�7(��Y�b���W6x�+|��O.J���
�j#^���"��o�L��f0����|��q�"��vK�F4\ѻm�م�ﭤ���:�g*���*�&LpM�M��t������Q+AҲ8�%��lm��Z!��V�b���>����*��&/���T�'���'y�>�ܩ����gg܍rp�W�M��f��hh*�8O)��]�:n'bg��WٲJ5&��±�)s�N��oy���X�p�
E={��6��kȖt������O�F�R��M�hm�_O.�
8��{˦���Y�OG�d�F�vnxa��˧���/����8��={DP�u�eC	�Z�������i��!%��ϪG�(n_T!�V߽H�i���*з�zs�[P6G*T����HH����1`c,F�k�a�F<���!r�]���ӆ=���[����!���@�����h�:p� ��=��3=4ؒ�ɯ���R^��=�}�]���?�|�{矘��|fa��#���cÌV��`�� ��|,PT>���y���r�/�fɲ���0�"v@LH����Q��/�厢ðS����l�K���B���r�� �D�}:�v�a�r�v�L*؅�J�����:m�������h�2p8��p�Ds$˕=�ƌ�!\w�z]d|Ѵ���Y�5��i!!	�e/L���:��g(,E�y뜬�ւM��8`݊��e��3��G��	5�3S��m��礐����-Q��H^h0}�L�_��cC�H�U!(�Pr$��K~���]6��Rn��-2u&\~�$ܾxثU?-�]/؃c�OK���^`4� <�K��(LP�V��;�� �~�ރy����Q�.�N�C0Иh~�����D(�u�Ҍ�U���:�$�}���D��~��Sh����J:ˢX��(���-4s]"K��A�⎃�����m�����b������>����Jr�P;V�$JQnA��wjo�@��tGBWiCM���e΍" 1����i9�Ƥ.����od4_�P���&������>�'De�Q/Կ�8��d�� <�Huc�n0hEFu^Yh�c����!��Vzbp~��1���ُC8O��Ƿd�MV�f����뻻w�k��kȏ��@ �;/ ��lY�_4�$K�I��V>>�k��1�\��ɟGv��q�y���fO�Iq��Kub�l+e��C�P�,��\Cj�˭N��K�����,z���m0�� P8���M�c��ٙ�C��⺡���,6���E�Z�	�z�3�N��3�oU��X��f��v 5��t0��O�a=����EJ�ƨ�[js}��E�ٌ��8b����p���)"��It��L���*ɭT��yw��ن�1_VQ�el�+#���.n�6��L�E�y���H�^���2��#de��CѡRI9HfB��Ԁ���į��E�{Q���P�b_j'�t�y�7z9���$o{�n�e�	��V�rO�I�ݓ5�SůS@j
?u�@���{4�5S�#�-�W	�ک���mIHhU���}C�s o��z�ߍtF���y2�:��/�D��f-�c+�A�m���{�g��H�~�m'/��_���L�����9���JH�R��y�}���5�~ ����(�>ʖ�وݷ1%���� �y���" �1 c��?xY\���&�mk�c�l��2��0��1��*Ztt`�*K�E��[�O64Ft�#{� ÿ,1�5��;T�ǟA���	�j[D��F୭�gZ�^m<(���6��OY�#��&~�z<3��B����+���lWIp��p��CR�ukX���HC�L@F������8���F�n��.ش�!K��kļ��*>!DUW8Z���of���̹;�����(�`�
O��>�Ͻ�WhP������F�<tJ,e�龰]=����$E
L� �����U��aJ��㉖mMS?�o�ً��-�vn��U:߾W�	�.��:QpHk�̘+��#�׸�`=ق�.�L�P���<p2{��Y�S����QlL[�B5螎��t��X�M�ٵ�tѣ��p�S=�i�����?��f��<�Suo��"$7psX����H(��L(�&_k�C�[݊��q�k�Z"��n���_El�\�����-R��~�Z_�ңs���5.�rYL���i���5���o%*����]CfRt`�m�^�\�ㅟ�<���n�R	}ڭxߝ���5����?e
�S����"�%��I���a�d��ѣ�Ͳ�����*��Y�'��/�HJZ$���S��(�F�s��?{K{��
<շ���x��x)�5��һN��E��ٿc�r�=������tY�����ڬd�K���UZ��٨3ӕ5"US���cC��b��U�j����7�*C��_W�4D�￧B��d��6��O�=+�ƶ�.�Yy��H�	)��q[;�>&c��66Iy�w�ꋬ+v`�kj��L��&r��VX�U"/���m�ʜ�9��I��
�U�:2��	+��*G��Lo�a�5��U� !�L�w�(����k/�� "*$a5��z���C��?=m�7����S���H0�����iS
�2\��F$>:��	iU��a�6��ѩg�5Q�p�d�����"����u!���
�N�-O���7L�kS��`hf��}���^�QآNF�j���)/����iw��П�y>�9[)0 � ���?������)�%e
����84����x�a��~���y�CH�8���a�����!�c�߿taD�=�Z��qB��sC�
F����d��E~��?�����|�[���A�{s<YJ�F��v����5�_���D>��-�'@�j��m�����	����?�a���q�!t�<�����I��Wm��,�`����͓����fR�Zz��f�Kt�ɣ���픪6�=��A�b���7�>�o{o ~�����$�t�$�y\D^IC���-3(�\g��m�i[�N�0���2��m .��y�����́�|ڣ8څ�y�ZTIY���`	者��`c,�&,[�#�{줡Η����k?�B4Qh$��"D6ꃩ����|�o�@��V��h�:�y���uO�#��q��RS�$lf�I���㞔�R�YT�����X�y����u�fpy���0��0�$��=�2�>��W
�z�F���*�֍t���&X�,q�Ϛy��	/re�(E������U��6ݭS���╅��W�>����YTgnh~�!]��GR����˹Ļ��vv��Ҝ�����Ø��p/��2��-P"�'^�ί�	f%�6
A�A�<�`Vb��ҀB������,�I���b�����^���U�(��C��8����o�e8��4��2un�ˊpKa��.�5��h���B
���O��\�QL�v�o��Kp��I�M7?HU}b
�_?a.f�u/|�w�b��xr��E��Ժ��EX`Њ����d���~V�(�_[pzKݠ�)��T�`�E��-nO�Y�咦ؖ\�'T�+�1�9����,9!��b����	�C��	R�j~%6��>=g�@KBW j'���P�k�Ï�\%d��ǹuOjP^d�qXM�ڹ~/�b�lY�&�c��sDs�%/������i- �Ì�6�c��G���M�I��Ւ>ߝ|:ٺL�d��Kn���t�"�<{��b�镐��;m�5�z�Ny��iN�iBrS���Qwr7�oT۸VͰ3��:��TO���X!���nݵ�t���F?�9t�蚤��I���4���	�:�Sba�����������)/	���lZ�����e�Ƙ�Y�2�0��R�JqD)�i�;m�=��f���2)A�W�v�����һg�T����M�ͧ�nd`�ϱ�	S\q��IG��I�x��j�Z���z�e��rf��)�-������0k�-������[;3C�������=���I^q����^�lҵ� �!����i2��(dў������4 (H�_a �v��5:BY��e�BX�Z�ZS4��D<)�cx�Vz�x�T��}3m�t狤��]wHj��[i��m����L����6����'�͸��"-Vc��c��(���, �Y�,��p޾4u�v�@	**��i5N=ywK<>�����q����E�hm�c)�e&�����̇)[ˆ(�iZY*��,��)QX�l���Y�O?0�p��	rݕ�{Dx�^�%��G%�?��{����=�����}�_����YXNy��j�A�z�媶�PK   �X�X��_�  >  /   images/17d126d1-8a97-48c5-9cdb-beb53ba7b71c.png�XgPP���:�PZ�� �*"U@@z $*B���ބЃH/�� �{���ޔ�q3��~�����̾�y�;�����}1&F��@
<<<j]M�;�|�cd$w�Qs��!�ձB��qu������?��dCjY"�<G8������<N��.b>~�Y�J���!]Mu���=���v�/�����z[��l��։�Ll��BHJKu�9P��	�P~ۻw�����&2��D Xj���=í��¼�E��D���(���\��l�_4�(U�qOؿQ���;r�s������@u�$
��P��a׈~�KfJE��i���3���tL�OO~�����~��.L���(�,x�����Gy-�Ō�*��4�RϿ''�����42b�j�����-�<��v��ZJF��>4z��/��z�F�8\7d�&���>���ؼ�����		/���s���@<�fa#��	����09�z���ڵ�P��lI����a��>sO���72=1��SI�Y��'���哜i
~(�#Z�pG�<\���ssr��`�����B�)��(΅�����Hj��Rrޓx"S ��Y��]:��CΗE5�V���m-�"�ǵp���eD_Oh���\��V��B�����I"��u�X�i藻e#��D\�(�d�s�I1��]^Η�N��v�0�h8 )�37�+q�o�F�U��x��Z<��W0�\; d�ھ:�m�gN.�+��R=r�c����MZ �	��3Go1j�֩��}0Ä�"��h<\�IO�뱀�"[/��'G_�Oj�t��������u����J�s9�੣�2���]D{^������i|L�M��eW%��w�2�
���0O����߷�qZ[�B��,��@�Ǭ��ۺ�{mG�k,��0ZA����S~e���X��p��d��
]]y M��1^?Ν���e�e����:t�w��ۋ�5�ψJ7�N��՟юmB�A&%�$�4Z���Qe|$2 n���9�Wmw�����[��S���%�z~�9�T����#����W������ɽ{X3�p��1�j�I5}J�'�*���X�9��FFZ��ɓ��J�0ż|�̎��G� �^���j��O5^�z��iz^���Ky'k��bYJUю?�f9ϑu�����2$�busK��=(�|��n+��*�u�R���񎔀��w�_s�b��#d�?	\l.+��1IO5�ɶ�`OP�(��^��eM%,?�������=�i��b�(��P<kk����ż���`�	o/�Umqnŋ�_\�iq췪���b�yh���\���][;)�9S^T��k�J���$��jo�r#if�fNj��.��N*<� 7KK1�N��V�d���,�CZ�,�es�iDԷ���EV�~��C�s��3,�,x�Q4[a�mg�W���@IA
���Gޢ<��w����i'\}}�0_ϭ��?�p聈�R `�Ǐ���F�PPo~\�2�B����d�.�	�
|-���I�H˖C�)�wl�9��zwӼ��_Yy����c�ZsV�dn��530�dtv��8��"�:ZZ2�0��r34ig*p��&����e���3�Z�"0k5.�+���IР<-Н67]"��Ȗ����z�8m��eD���[� ZJ��F��y�>+=\3')�_�(�H�9:	�iɉ�18����"2����=
�t��G|�(lc�Ÿ���A�����s<��<����e��z��Ht>�MJ�!�-�CL$߱���G�;��vӰ}B�'���#�"jY_1��X$�ˈ��ω�U��Y֔�I#s�nAl�($J���ޣ��i!�#	Jm���h���j<�Kg�Tɮ^������������*0g�������'���_O��
�6�ҥ��i�>����5 �\վӏ��Kz��ZH4x�h~�s<!i�F$.��#w��;nO��h��4xG����^�o��a�����\�/��EDN�q����$��~QqE���4�&����⧳�RQ$�ҹ����\o�r)�P���4[.���HR���Ie�h�g����J����g1M�В�hK^Á�kG�7�����)s�������-=O�<Ɖ�^d\��.N���u�0�iݲ����`ε?�8��*1/�o�?A'�p��a���	�vV@���\}�$o��������K��\���B���`��ɐ2����ᗰ,�*�ow�u�uT�c�RA �M�e$�2yt�l4��Q�͏�~�>���R9���kU�^*��xλ(�;��z����vf)"㕫�g<�������ϟ������i�G��#�F.�%t;"����v��k5�EE$%$$�$�@��nS��f���e�M���ө�ѹ���gTvڒQ���=r�&Gt^�3��s(��ok��͆�R�Z��,�1���,���B�KYo����2����|L�l���U�[^��O^����
�����2`�Dy�0rQ*%��y�Fs�K�`v9��/��MLL����P��3������͛���)�v�P��)����>XCDȇ�P���i��'?:��z��Yu�����Vz;~\�D��1|��o�s�4�z����3'�D�Ga�/څ�g��~P)[v){��!ejjj_�GWf��ﲯsY���%�'��_hSnN��7�+���$�ak�
?����<l{#WG=<<b�Z���;�IgcY+�O�W������o|T������o\U�JG���pW�~{�Dbv-���F�	U-zf{�|a�/����+�3W�<Tm�p5Bm���-�[�F�Tra=8�/�%���}�nT��^4g�i�L�8���h7Br��)���B��ާ�ϷV�5 H�}��B���q�
���-Թhj��7Kv������
�S�^��	�!r�<Y�\ �֑ �\�x
++��Ly��ց:]-�8}��F�i�`Q�ilg��˲b�{k����>��C��>����%����2��k%�:�賋����V<mm��g�ƒ���J��h͒,��h��"4�� �P]�(������>�}�'>?���ٙ�J��	�o4˳���{�v� �rl8�A�$����-�,�]����(��T{�_�����NOK��ėj��p����3���]�d����fP'8���Mn����&��"#EoD`D��B�Q<"3���$[D��a��^�S��eïI�ES��y�����\x�Ѕ#����^�
���O�,Я��@&_ ���9z�G�-He��恔'���]Mm���JϪq��^�2�yJ8f��SI�+��XHN�PD�-=���o��v�"ڋL��I�A�c��JKu���0(~*��,[�G����
v�:�?�p*�T`��dwpz��o#���IM#D� �C��y��,G�A�b�QR��D�M�2��&J�����C�� �:�>jn����=T�DD���&kYiW��	d��AXe���k��`>o+ATO�_OTĳ�|�`��(�S�)6��$�1�T/aً�,��$��K�浨��X�e�L�j�é��x�[+���V�@��1���p=����&�S�B�z|�N��ږ�J�YL�?���J���!�A?)EV��+HLo\��'2�f]e�4(ZL�;��0�|�q$R0_���GN�9#Z���"?QGf�7ǉ�+�O�+D�o|�/Ҋ�W�N�p�2`�X��~ֹ�&�y3�U\��Ա+�w��D�6�-�!H���k�>��/��V���АK�۝-���j�J�>�Ւl����s��������ݷk}b�v]W<��}�يo�K��&�W֑�1 ��<����/��Q܆�=|�ID�a#<<��7ZL�1 üTFg�*��75�f��p7����5븥��a���˵����q�ڢkT�y�ۇ��M�-A�c���g�D1Ѥu?6=��ϱ���\��L<����ֲw��
,��l�G0�M�j��/��ޙO04��('}��F���h��j2�Fpǘ:X�L��'�]V��NN�%�&����	k0�&��u��}��wA�}��\{�����f�do�F��A�j�RbC�&5b3I���R	c���himݙ�hݩ/�A�,��S�X	F|`@��nH�3��_�L��2/۸��%����v[-�?�Zݟ�&zapj��$͘m�!{�M���l�������{�?�$;I�x�oh�.
u�7�!���Ѥ�b'|s�zg�-�e�H:`A�^����bk�u<�꟢1�,�볤�s�0�P���W����^��Pi91����_�g��m�X͎|8�}��L/x�(Ј�����A{w�~��5�N��Yv"w;���>e�(��Ũ|6�h��(`	��W��s��|z"Q&$��|I�CqR#���W��C�cYcھpw־�ϛ����O&o�٫���k�k����7ׂ�c������F�}_�<J|6n�ls�C|�hW���e�]�	TT���$-�!�3+�r�ez�8��8�3��ۙ����7��c����'�ܞ��� BP��;2d`�	����<�Y��8U��vt�n!���#I.���I�u��H(ueY{��k#�X��|�5�9|��y����P��>
G�U1"�E6��Y7�~�IP�� lBy6'�T�m��Ҹ�}&^�BD
��#�d�_p4	��{��� �>۔�o��렡��������+C7��س�?�q�/�O<K&ʷ�	�)����*;�.�q�aD�ב���~�K����q�o�rF�Nܣ�Vsx��XH��������?�����`�s��%]�~t�U�y#�磪Q�Fn��!A����!�x��=�)ɛ��dee���2�9�+ �����W��'�fzqV�.��j_:�6�Cɜ�&�[n3ע<�S�P��d;�0+v�M֥��9��>?�8Ra�TЎc\�����M�3��vH(	�������dy�>��R�u#��&Ʊ���F�8���%�t����l�^6;�4C�@�-�^A�4�����?`0�XY��ʡ~����@~Cߔ7[b:��գϻY4�{����+��{w�Xgz��D� �x��K��������^��h\�[QCC�a����0���sħ,ߌ:��h!>�^��:6��"��*�,1�<��P9�.951Q�iiiѥ��i�X�ǙW�y�I��>-��g��nJ=��Z�����t����AX��W<�kA��*����l=���� �	4�ި!�$^�3'E>zN���MP{Eu{&�����ґ�_l�ߓ�����,���b���E��|����$i? qU��H�[�#��z���'�'��U� ��n�T��rx��l�O2EmV�SQk�$)�����A�~7����Q[i{�U�0��&��5ʖ+`�S�遇���ۨ�6��ɎZ����Uq�
W۪��N�PN3��'�8��I��������)�>[�x��*ب��i�}�V�vK�5�qM��{cr��Ud ��)�^끕^�'��i'b�ӥ�� ]J�F$�tn���o�t���b'�.��Ï��%1���c"�O�K:�J�/�<��o �� ��\-^2�7��)���%�Ա.K��ՓW������*j;����m=�N�jGI$ɇ�tY��uf�J:�(V���*��'�b&�̈́�s�NN$e��9[e��J��R,=2e7��lË�T��T}��N��U��>i5�1+��W�X��Zu˿�\���ն��"�c?
Oq���^�|n�~qz�؁�ӛUUu�0/�Ԭ�``=G�#_u��E�֝AZk���8�&�O�6L�a5��'��%R#����s�;�8Vx�-�%��V�J������V8��i'���ȹ!�*S}�`�1�WM<|r�9~����rTYq��A�,q8��j1�G@p���W�;��o /�4C^�����8;p�!���W���C�Oo�REӵ�}ձx[�o�LI��;U��ə7ޜ�.�f?�C����Ozi4>����>�.�XhL��|���V�n�nWf�l6���Ǐ��ӈ�#���z(�ǚtݝ��E�E
IYeq.DYC*��F50婻b:22t��ITi[K�t�ƹ�}�tFdYt��j�"<j�g��#���5U��}6����ӂGR��τ�����ʭNx'�,��.���$F�tV4���Ә2h17�D�Q��ΑY������t~���������-�A�{�x���u���T��q7��S��ˢ���t�����W
0Ƃlf�G:���/Z*x�:�!��_^��\�u�I�)��{���� <�;�"�lɺd3��$�"��>zf0<:�+�]���<ARwPDR��&�$�l�����OHiD�o<���xw��e���8��PK   �X�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   �X�X�z���o U� /   images/3076bb86-a585-4cba-b1e7-fb1a193624b4.png\�uX������-"%�t+�ݰ�HJw�tJJ��%].���H,���H�o���{�q���^��9�U��9gb5��q�q@ ����6�����1�o�T� ti%]0�
����vU4� ��������%������������5��Ǉ��������5���m��85��$�J�7gw�/����ᖁm%ԣ=����K�,�f���s��$V�̿>k�^{��a#�Mԛ�Om��������s5�Ua����8\��:�wU]y�9��[4u��lɀ܍�`�@��ʝ��ӊ�%��䫩�� -A����YG��49-qme5�
Fe�p�+����L%v:f����J��5M�o3�����QW6��.������^
�d���Y6��U
i_�����(�9JvI�#T'��2vJ�Ĥ5Ȁ���T��w�����<�L������C�Nxu�j���x�"�6�c�'��.$������C0ܘ	s���٭;
������]g��&ϯo{{�W��C�A^wH�
��1f�%�5��D ��4=�q-IP��eu�v��B��X�0�!X\!-��ş{��e���+l��H������V�e��lazZ^�,Ӕt�ȋ��	Rǟ^|4��VI���د����B;z�>�<�x݂חo+h�wT�䑍���� ���6�&�gu��ղ���[Vk��E�$��&x�$ ���G�B��Hy��h�C"d{z��s���{z��H"/Pe_f �F8�J�+AH��g��6�~T�.G�<'��>�,��bFlh�Kh�w����k?.yQ(���
�2����,cE���򜴷��ȁ ',�Bï�S�h����ْ#P#H���yg����4:��w�����Nl&���e}�i�|��������Z�;T^���^a�r��E�p�,`X����i-	�y(<&������&����`���D��<�Ѥ���w��1�F�����r~
�m��#>��V�]�đ�]��li�P(������!�}j�Xk���s��`aN�ϰ��"]��O
��J�&<%��*��py�����^�f��{\�|'�N辴�#�l���
w���GY&�J'`�R�����d/��z���L"�L:��h�w����/�^=�WbgE�xܳ�n�v��䊘a*	�$A��y���i��w�h���n&jX��x��埪S�EJ�utV�JFo��Ǉ���fk�ȟb�#���%�&���/�U��^�kjgc*�-a�fF�\v��߉ �)	��N����L�Q]2k}Gq<��N;��X+#3��0^3<�� ���>�oEլ��cǶ��-
��J�(�p�b�/>X�E�I.?�Ŀ}�P��A(�������5�[R7��;�-�őLڑD��ȿkE1�p��α�O���g5w�a,Eu5��k�bZ|H;�c���r}�t�������U��������;������q�"T�u�#�����
�����o��eJ�(�W�A��s��\م8��<V�������N}---j��,��戏��Baȁ*7��(��q� ������C�����ع��cd�(p��������){�T��ңr����Cw"`��PQbp1�^��C�$ڽ���z�e�i����޷�C@,Lo�8��!�Ȗ|��6/o��q3'�O�fׂ��i\�	sKá�o
~y�3��R�5حB��-���&7�B�#ݞ�N\o�ܶtpރҋ��Ǿ�u<���*����7+���--6���͔�g�(�D�B�����K]��c��R` Oq��D&-��pI��2 ^��)���)�`�����eC�	�D�@�^�J`�3��T�sB3��?�Z> �o���l�&�d�f�SbZݙȹGگ-���^yt,�ip�梭���䀯�of?�lx�e�5��b%��
Z-+6�Q��ҴkȬ�ƶPXm�"s����ޠ�`g�٠hV����y1r ����y8W5��eZ��Ѵ�5�*�K���`ň��T:�Ƿk���~D�w�8���mP��O4�ѝwl'���7�3mo��,�ļw�_y��/�/�,���NƳ�LDy��|n��'�zз5>��Ҟ��	��^��p���:�KKJ������"�jiSSI�)��ҏ�A�SZ�\f��R7����j���d�:��!����Hi�̰������}�-F�!*ю��=�����Us��&)���������;W�"��뛖v��\�ORiS�Dy[\FZ}��@���F`��K?FY�3�����2H��~05þ���ȶ6W�!�E�����n%�K[P2��n�)��.�	�|Z��Y�#���ʲJ�*ن���@� �u#X]��xډ���I��}��f=1���U�~f*6u��t�|$ѵ'$d���he�;�40������^��8ÔW\�
|���oW��h�y��#��ÝG|��`�+����r�S%o�Z?�O�mք�vxB�i��O�V�^�`������-�]���A|�0x�d�rhhJM.����P���4kV3M\i^��k����0�_bf/>�q��ɧcQ���C��;��1Z�2#0��Y����{o�k\x���Ҏ�A�E��x��xιݮůz�J5e��1a/��4KoQA;�nSR��k�m�h��i�y ��O��[썌�ڦ"���#KY�r��l����6�_A]N+�!mZ�������H���y���$�{�U�?!��킷�	������*�Z�3����"m�V��N���6�E1痯��޻*��~��F�� ���O�@7ZZi��f.}�,@o'R�4��;��Z�{e��~�)�	�ͳ��S��M|+�cl�	8��K��zӲ,q��S�8_�MF���c�ge�<_� 0e��ݡ}�����������iA���Y=��ʁ�Q/t	[8��|#�PI��'(�\%�s�j�b%�}������}Y\�"@�������z;Om'�M����J{���bV�J���L'����sH��u��Ű�I�h���" ��A=�/Z3�EY�<���on�� B�F!*�h֬�6E�~�<�CJw�L�pP�A����g9��<!Q����M𑊩��̩�y�i�~u� ='0u_f������t�'���o�P��r����v����+��7�`���M��y��F�ݖ-�p9biq���p ��+㙑 d�����zt�lCL ܒ�-^�2_ZAӞ�:�V31�$ā�za���hI�#YVĿ�T�r�a��-?+ퟗw��ێo7�\�J��璇�<#���R���Wq(����9��ڛ{�Aˆ4��5[ '�E��:���WVV��|}�ǋ	\��Q؀B�
D�$D^+m��B[�`R~��a��[*�.�1싹����2�wY��*�����6���)-�}zFKp���X�}�g��_Lb�uq�$�d=YY�ރTd�f�y��+��Q'�b��脱E�A��'�-)1�`�i[c��~�g>pH����i�afWo�����K1U�'�!p���_D3����L�\��v0�|�'��T�k����k+��m�"���,�g��(�p��J�X��q�" ~8�o�r�����'�.H;n�V^�y��=�O+K�(��p�N�<�Y0x{wtm0vq�Do�c�H$GyU;;+�Rw7���J�kC��p����K�[����� be(�g��WF{h
pPC>	%
�<�r�n5�ai�9lqj���-�E�,e��e�R"]�^?�a!�8Ը+�ꬴ
K=A'}��^�"t�-�]�<�׽W�Tl��ތ��g�u�Y<�|&c�[s"�����;BQ��Gz�9Ȱ�mͬ������N��VO[���DS�N{��V����k1/��agv�8�c�IIM��}�S&2kǃxKJ�`��ߗ71�[=�����*!�J�!H$����/vGR�mU�wp�@:����1�>���{)�/{v,"?�V ol`{#�p�}\\�o��&�y��Gv�DZ!��L��N�����a�0^"<Lb����$������=�VӚ��kַ.f�����u!c4�m�:A_�!�����
i��5���ƿ7��U�ӪżSە�B�Q.���v���׭�P���"��E���r1����7�3��ŕ[l��Ԣ1���xb[����#@I-#��'d�<Q `�V]�?C��G]�Z~��'�QY����'5���� �޾�b7W�~��~d[��q'�4��P�SW�6K*D��V84���Gu�O��F�d%⊘�����@�=
p��)�Sj�Wؤ���&ˆ�c���}_Z�L�?Y�R#Sò#��@�#�����dW^Z�6j�&��^s*"+w�x(�D�߉����v��+)���V�k����+f�����p�Z��A�,y�|w��L�g��������XrU� ��#�����G?c�� ��i!�F��x5��֒�Ч���P<��Y��" .2kC�.�_�Q9B|��,�Bj�������Q{e|x�'S899��Q�3?�8@I��<���1���U¥VO"I��x����<�jSp�	���bt8ćn)�کʬ��Y!駿�#���׋��h p_xH�.�Y2{F{��#�g����o�0	hc"q)^�\�^nfWs�@w^9a`
���M��������� |-W���՛��&X�]�E�Bܫ]��D�}��j��3���#��_�c�,��{v@6bi��)w^�j4�B-{a�lcVs���/�q��M�e�	V��|R~{'p���-
jX�i���T8���J��?�4F��^�
�B���T���X�񹹸˓�sO��M��>�\5�I��|3_/�:����0���Q'V�������^J"#۪7
U/y?���D1�.n��d��6�E��;
���6�`XL�<���_W�¯��HZ72LOkC�Ƥ�ŻϻV���B�z���N�������c�`P����=��6 ��7F���P�v���5��L�0�o6x� ��v�HeA��Y�3>m|�/��W8?ߙ�3��%
�˧J�<���Z\L��'�e�� S�b��_N�C�"��sn�����V( �l�-u��6Rj�?v���{�Λ�kp䚉���wn�[l��p�M��<����0/��@P 
���,��~�:g�;6�l�\�P= ?%�Eo�&�']h��R�o;���z�U�g�rA��'��8ɿw�:����&]��.C�0F��T�s#Ft]���]BSz�@� G��B�҆��o(Ͼ����5>���W���#�tT�)"M�H^#l<���J+�/A����g�:��/�`������4�'����E�3K�����L���(��\��\��MJ�z�>�^j8�\cL��Ѐ��1�������!e2�P�]����[��LK�p����<3���h3��y��ѳޡtN�v}/=*5��
��*/޷s3	�Y;�'�o��%0�/M��G�h�H���p���سKS_1evb0:A�����N�|EG�b�/�LUb��ܿ��5"~���gW��dN�Q�=/��?c��rD���x%/��/�Ӗ�d�iۤ~fX���K��꼻B���-����6���@m��K�����vsWZk�j�،wT����?�����,Pjz������ޜ�͓;��+�Kґ.�@�ٔ������5���_{�OLe�����Ó�i̍~J05�ɪ�pdwx���<V���� <�:a�U^S��=���ٲ]�Δ~��8�A� {SNˢeP8���snΔ������=s�iQӪ>IޠL�&����&o`��}d��Y�۳�M���vߍ�ܙ-tvo�Q��;<� �����/#��5�_s}�>�-7|���8�	���}�M��m9��nZ9@TO���Z`��g�}vc��2���$!P<	
��p��#BJ#�{�a]"�-\��51h��h9�0tܔ��y!�����P#�/hm]����gǎ#Bj��lɲL]fZdiy���`aZ�=�(H+�e�s�  A4�z)A4�:J��?u������GĮr�j���BID�mY^c�YaO�A�����e5�'	
s_ə��-غ��O�|��J��s�P���R'����y��rw�)�;h̸������ ���2�[F�BH��sf��:M��DB�J��Si�L���	%���V�h�{?>ߦ�
Y�1�RH[�ѡ��O�h�u�sU�D[��	��nw�����Gs�r�����U8a?8?KQ��Z����}�1 /ZPʏ�^�;�7����� ����b�"�e:����X ]d^h*Kg��T�Q����C���8h�M����A"m���y<{.+=0�\\\��m[�+�(77[R���7[	�B�x(��i���5R�%c[�_�� ��Y�&q���9⎭AB+�����f��@~7lue\����.�,��!��t��_�(�!� %����.O������BȊ�����E�iR񦼭rMԞd>O��	Y^JY6�!�����G�=�tܙ�V����������X��{[cX�s�Y$q$���$�6&�{,��}��7uM�p͝;��AZ	�l\�tk����Y�	��0���d�p_9�w>���7q�G��Ɂ��Ô���ڡI気���B�C��}�ye��������fO�MĪ�t�UWW������ԝ������0.WQ��i���m����^8,�}�8'�-� p*�dc�2&@O1��[�
���ˀ���SjOk�}�����F�bol��V��Fɯmk�{!��M�hmM6y>�Շ�|��w��-����7�g ���};]�$�x���"�[aڻ��9e�Q�&ۿ�)/dנ�J�uQu��G����Qzy�����/G\֚�f0$��I؜�I��u�x����k�^R�ԋ�-����(���lUa��@�bnn.�<l�wn~~|j*���8)ZvwemmY��������E7+EWb="�jV7��.^����K��sNNһ'�w5�A�?���.oR�rW5��9�_cb⋰���.e��Qg�W�ؖUR�Ff��l!��,��B.f�
�l����{ �{�;$�����X��p���:q�"4�����I�_E<�����Zg�9�ݵf鿋b\�9�g�U [\��^�s�W ��5��_�z��Jd�=�L�Ř<�Ծt�S?���K�Vb�u{�4�"�5lb'9s��;K@��*� ������Sw�c��㧀�L�	�����j�����6)?W�y	 q~��<E�S�]h��:w�y��F�v�^�qv�qDh![��^P�v\�� �g:|x�{�`�Q�s0���P�ۻk�7�6@����=C��gn���s��MI�&��,=#����<�a�~Y���OP���{�Ş\;�⋌fSH�C�j�^�":ݡ�|��ϕ��{.-3/�^�x��l��q$�	���v>Fc9�W�6ՁH�T���,�:ݳ�PQ�.�L��/�
�w�Yټ�dv���b��[-�UQ�H�
(�i���L��a�k�/���Se��?E@��^A�5���v3/�,���z܀4���R{DI�	��es{�)�ۚ�����z���S����o������t�J��{�.{n7�斫0�#�#me�0�<P���>��߿�&v�YO�;:&�e���Oޝ�y_v7E��#�@ r��
LZ��gyɍ�d	t|vS�y�#/�l��T��N�Z�t��0��,�gu����c���ڝ����!��x�u��{@�
��NW��m�.K�UF���d�� ��*G��A���"�9����1S�J�f���@��B�-@d�~H�O&Z#������؛k6lq�C^�[H��t���_�ks��ֵ��[-!;�(�<
C��7�
V�����b�Sa�`�_KKy���m�C����#�k;��*�98�s��Mu6�Ƌ�so�>
�m:y*x��H���H��d�oA5W�ׁ��ӯ��&�g�Tʳ%�H��^��!���KNo�z�#�V� ps@ɪ�i}���}s	�5N*�{��J������c�\|��8SZ�mM</�Z!�0��F��j�5�8*�YP�Ζİ8��9E���U�L�k��S���mX(��u����s�/�x*�Jckjj�<��N����V])YXX��y �$9��V<$��򠛙R��OV�+>OW�H�,\hir��j�oI���w�<y�����&*N�n'� ��yQ<��{VsRn�����F\a����`�������@Tu�w#��Pӫ?X�e��G�N=�߰oH���+���F�����`;���D:���jzB������ن���\B-��^�.D@��J<��3_G��f�O�,?C?�먽����%���!�O��׹Kd}||��V�T��&�� ǉTMJF��0m�ؖ��^������A���w氋�$M[WR��a�y���*>(��}��;I�d{G!�3�5\�F���M�c�<~�\���:�c� PKP�u�bVv�� ��ʔ��@9������h�2{=A�y���}����U��'�r�K��  4�iǸ���	�(�P�����a��
!��l��1�iRͥ1����_����:����C�I*n:���r��zB4���l����7�8�Ƃ�c�ɟ���}�R�B�d��P۫�R5��#���,���G<Q���L����ZRS����${��.n��� 4�?��:Z�&8�O��5��=H.�m�n�S������EM?��<	�f�όFka쇊�=�3%�+qz��@�t�ǅ��p@ىĕ� �6�>k��i
c�p�d��v�� 1������%b�x	���,�u@M������F̣~z}�>F��e�b��*���\����Hf�m�Ӫ�UQ^Ii����p0�Qw�kc6��|�o�\!�˾����P�&���}��u@%���@9���\RpPs[_�U���=.3�U��y�m8i��2�Ho�
uPV����<{ft4@Qx鞖N>���g����O��T:�ȼ����!n<�蜢�hQ���u���kJ�b��'��
�6Lu��������o�b�:$��L���f�s_�	��͏��u������50��*f�֝���eX��Pe���q�AԦ�"ނ<���7�������P�t�;bWkYco��|_>XT���j���pTNk�'x�ǋ���y��&I��ϒ�J�����!l�|�mu��Ӄ�`>]M�ߡ�\� ��(�'A��`����|� �oo�AMCc�2�!h!�]Z��ʰ��z~X&u��$��e���h�Ԫv+���R���Y��6S�*+��x�ȹ]����7�ɲ�)ƌ�_Ƌ���~������ *:�o��.���������hJ���I��izE�U�,������G�uV>��X��Tv����ɼ�}g�?��{��j3�Bfku~@� ��;ѿ	#K�/����ȿ��c��dq���*�<����'�ӠX��f�Xx���g��.���Т1�"��d�|�>��|�T��D���qjW�<��kϚ]���{��~K�I�� T���;s�cJ<c���";�kA�$���|�8�3bbrdI;�,�>k8�oE
���=�t�S�)u��h324L�#���ꐟ;@�7�V4֌�R��ZFݚ�ez0��t�{y��~o���\m�	 �(���S'�Y[[+��|�Zea9Jd����H�z/rsP,�\���z_�q�Eؼ�xZU��cȦ����[F6/:�m�=�&����jY)����u�{}�=�e�T��`����}#5L�u����6��95�:��yP�.au=��ʢ��/� ������@��-���BK[?q�.�<����|���F���}��G^gŅ�|��%
=�Wz�`ZI?����ʮn�e�~I}{z��i�*j|b;��/=N䊧()5K�K=���P2�&�4�OE|Y~s}����^xw����}
���D�'d[��KHdZo�%��'�4��i����t���m9њ7ރ�ҳ�}]���>W���F?pJ�t�e>�;�@�}K�w�舟X�b�����i�:��
� ������~}���`�v]8��{�afY����2QZ�a�6�Z[�US9A��9�)���d�������;��X��P��*�KM��g���U��#A}R�`�Хw��y;#=��f�l|i[�������Ƨ����sw,.�~�e�w&ME�ᙜ֯߿�ed<ڝm�"?����4���@�uQ/���oK���'�G��Q�&�U ���z�s�4����������]r��v�}M�r ���Xy�9¹S'!�wM��@�w5���$N�p|�܅�/N����6�Rҩ�]/�.��W~;C b)���1 �j�������:�D�c��/�Hh�?�&�[+��\k�Y]mζ�j�"p��O���HM�
p�m,���m�Xsg�>L�Cq2���Y^oٰ�� r��u=I������Z�v0\o?�W�w��` �oR6���?��6����B;H��~���e�˼3�\�����L8wTF�=�՘�%�>X���,����>Յɫ�|;�@}�����k����cr�ֿ�����(�V���r{�)ǔ�f���YFH����AnV�l�DK���/�\��1���SW��`D�W쟟�>��X��\Es�W��6��o|��;9��J�\l��Yj������f�����ph@�}�D�@RL̳u�VCƒ¨]	Sn
��m�" W�P?�É�^���5���ZQ��_���qqj���tO�2�jQ�mi6��w��>�Q�����������U���i���!���%���X�%�)�˅A�]K���\�SMv r�ŕt
����eu[��QP(ޥ�]��EH��m
�I@���&�_/��\�u���INy�=����k �b����aS��Y:��~�F�y��w�d8,�rȕ�D������,�Y��|�^?3m%"'��z�2�����F����(�JBCǊk���:u���	
 zgM�����W�Z��+hb��++����ahX�8����ι�I�J������v54����>��S`"��
�7(���uҷ�#�HTGr!�L�v��p�*���oc<X��XW��ݕ����tK�!����5	1�;�R�
;���4ٓ�WG���(����u3>�+�dk�@�|y�[11�ub���'$�T�Sa0��$��cX�aw���q����Y/���F=1��h[R�))��W�6=m���뙵IiR��T�D<Xoo�X{sKQAA�7M��*K1v��yŃ�7Rݒ�#�����F�EՋYTgg�_Cn����؉hY�}�[��'	�@�����´*��e�.G;���r/��nn�R��8��Hʢ�DJt��~��� �IăҊ�7�ed�1�i$!	M�,�o+�����;�Zqg��?�r�!�_^�{Rq���_�ٯ�
� ��y
,�;�P��Iz����ٸ�G8[�n�dJL�lն�[C�D4�n�g�����>�V<8h�������9��G��<<F��� #k��ay�y0�ς������/��C?g�_��R����gE����s�f �N�ƶ�O��<L��&aH,��-�����K�(�⊿���X�#,*����$������_�%
��9��. w�������p]���J<�&0����*��D� �Xq��*ɧ3` e�	X�$h	�Ib�H�v�,��@c�Qsgp4�^��u�ѩ��'n�����4�e,�]�>\�ܛ��+��d��тP�-�6._�E�<�U��-D�6�+�v�u��tg*2�
�O��%J���a�iriMYLm�����"i������ ��ʰ�݋o�.^"*HH?��V|��{�B�8b'��J�1�OA�q�"^��af5xsm��V+VxJ�v�������O��ȪLٲ�7G����TPP��8��NK����I��Ly�V|���V�1����p��~�]��C�ܟ�h0$R�tܳ}��`��i��˭���[�u����p'�y�`���|�WA�kK�)��ٌ���AH2 ��,�:y&���-)�V�҄���[�Ҏ�Y�)� v7�k6��}����͔�cýqz&"����� ÿ��,�~�i˭�dҚ�Ɂ��Q���6��/�HBn�{,%�78��C;��k���MǼڄ���}�A4Z\����8��Q�6Ӻ�=���XY&�m�1�k)Ѩ[���U�JJ�*�)=��
��8wBSn,�)���(W�wl�=RV�n�����Q]�IL$J�#u�t[	t��9QA�sIA`O�
��zI�ܰ(}2r6���j�z��*HǣE���ʩt����N�5����wlD`�:�^U��[6k(�@�l�\u����!Sˬc��Z|��싟Y��n� ���<�G"����Hub񡏴Oف�J@�r`$�,��}�\9�3lv����%몧# �.C+p�~Z�ق��τ��>������Ti8~�Y#�77S�Me��:ZZa�
IO�6���q��R�p��i��{��&�+���|�5Xn������+�N��K='�M����<QP�&�=\<� �����v��|�ׄ֫&������]�TyYY���X�&�0崺YJnpB�Mut�/O����o�v�j�2�\.WaJ�j�V���9l�S��l��%r<W���v	a������9��X�P�|{GWaaݣ����BT�l|@��
3}�����BNb���[?zr�M.���`�U�@�EY�~!�+��K��f`-�����B� ��J�P�(�y����%�̒�.�TقN_��9�o���4���Mq��~�oy~n����q�����=!�� ZQb�D�k{x�9w�n��[b���:���I�<J�r��r=�s>���{� ��X��_�c�9�Oj*b�]"��V�AX�����+��*/L���zØ����:�$�x��\��D�j;?z��SS�S4��K�V����}�#�����E�F{�����g��/��p���4���E-`��/��^��=lar8� &&.�����NV k5�����b"����o�+� P(-AQ�	�`7�&�`7���d���	eUH0's=B�q#L�n����õ�g{�:��1�L�x̫�U=���+-=�����YS8 ��E���l���y��({w�UkǏ���dVb�RV ��i�߽m��̆ȠE��O�Q�I��+��7O�n���}z��8��ثQi���T� �QvίCw���Ɣ�=�5�
^N�KX�֬Oa����MvĞ���C�Ѱ0�����e�m���P���_n �L'���m;F���mNem-��^	 ��r�Ќh�I���t];�Ya��wj�~��e��#6�u�[%��/���횶�,����&�Ҏ��(�^u";�?h�ht짮��Ը@�D&.�)����T��6a}��_�{�X����6��raa��Z�1�H�����^F�i��nlb2���k/�. YGY�T��5��Da�H�uv`]���"���N��>�<�n��>��f��
���tokp�U����|��CB
�\Ac#��X������Υ�w{���`n�?�ʫ��-[^�Fà��M!W��d�R�}���0�[ANTdD�%��%����eUω�w��_���9�%Ch�1�>��b>��N��O	"�n����I.�#���n~��-E��©fÂ/_�S�|;����UqO��8|σ�X�֛{w�ywH��_�j��Y!NxS)Y<�)j��5�`)V�nWk����p��)�]R����\.˶���l�!�����/��˗2��&vސ@~���pm`n2����ƌ��Z:�N Ɨg#SV�
x������ql5�n5���>())1��H�ܺ��8ׄ]�_��TC<eR��V@N�2���:q�i��ڷ����C���
]O�G�lcK{Ȧ��A9-^�Mզ/_����'����(�!M��=����U|r+�,Ѿ�)���6�*^E�߅w��=(�b[ZB>�!)��FB��S�C��B2}����h�(��IJ�L�͔7�QҌ��"oΗ`3]��*��"=؍��2�?�QijE��7�Z����2�UC~�%���-�*��j�`�M~���_2��w�n�>�G�96q��j��QG���s�z����;�m��}l��d�.B�ޞ��f�w=�RԳ��K�h</�َ_��s@t�M���F�T=3�Z��Ek���YP�`w�^nwqM�Q$���X����_SS��~��V�IUf�:��}s�o?H.�557��1qiъ�?�@�)k�%Pp �ͿWaѤ����0����!-���\�78�)��ym�(�7��<��'����=ح�W�4�%�@�{���OO"BGPA����v2�g45W�A!�df���S@��[���R8�a4l��t���%��u�!�	 AUj�1iA������UW3�`:�m"<�䚴�h�A�����Y�虌[��~W�@Ծ�Ѽ	��2��;��Y�;�����*R?s�'�D7�vS�����b�E������Kw}8�T^���Q�[���?�r��s�y��ڝ��ֹk����_Z�UA�6�н�p�\���(�B��t� ���q����FcLa��MԖ�[��11�� 3S!��T���l��/��x�3������B(��hn<OжJ�
�[��׸�V'������Po����GjikX� �����F�ep0z�O_AE7�Nl�����pv��s��	�Q���C ����g���<�R�5�9���ǽ��kX� ޭ����@�{�v��g�N<�ͺ�_����3b��^���Y=�?��J~��p�e��OU�>� ����3\FV��-`N��^A�����xq;�pE��?���kc�o�����Nx���y��zړ~i队)E#���N<i$$��)OS�������vjs�D>EٷM6֡mO���C�rZ��yY?��F�_ޜ�,���X+�GY�n��ܢ��>L��Y�ט�M�������=�wn��~�5�{����D3o�"�RU���O٥c��k��]!2y׎��O|��5@-�Y6'����� 20�;He�Ga�>����IA37C�![}U�)#�T�~n@�L�.��S���#�*KQD/�ߜ����1j�����Ҩ��Q>�q鯺�S�@yYpn�f����_XH�E��(��1�bъ\������yK����޷B��R�	�Y������j�w��H"vD���g�E3b;L)`Q11@:�zwp�.�(�����,��m�^�˘|_��"����d��|��^�v�jt��@v��/&�M�%�� �c[*Qv����6�{�JJ��qɨ�)>y����fl�w2����ԯ��D$��B�ss�T0���V�g�b��h����Ғ�� � HA��� ?��_��V��h�%e}=�`�z<�ɵT#�a��,��\+_�ww70���ac3�p���::���Bl_8�-�EEe%gV�ļ
�C��z�@&z�Կ�]"s8��ꪩ{�JH5���+299i���fԦ�訜���:s�<h�=�>b[h�x�o�;�\[=��{p	%/#�FG;V�jݓ�D>z�u�����2�ʍ���4~̒���iGBh�����\�ײc~O��[μ�3�*� �Z�9fj=8/��ʵ�y��	��J&��Ω:|j*2..�
��wr #9{�7 ��4�R̵��7;�-���ۂg9܏T2���oj�E �y�[�}`��.����lۯ��WN�	�+~��N�e~5O//@Jo������W����[�i�%��z)��f�h�L49e�rյS4N�|⁜�e^BA��dU]��A>�2�D%����H׎E��p;���}g@�x���)Ǿ|�Ɇ�2�ۼ���J@@@H$�5p��;�Hy�y�$�g��[��+(���T���]5uث���=�{��k��}���[f����������Gn;<Ѱ��  ? �G��ʚ�?H�	�e�B�ʸ'Y�XqI@�(��?-s�������R�P����(�T�.˻6혊�n�����+��y���eb�7�]G�)(`���?����к�rl�����v2y�Ή���N��!����)��KĪGm7��Z&&��'
EZ��y�����k�"�Ą���}���'R{_7��[�4��m���OQu5�����^ʟC���#�[�K�RF��o����E�������y��L���S ��S_@�[��{6��� q}�؀>J�H"orj��NX�1g�i7�+��*�?��a�G�9��+l���%c���"d�L�ܴ���	��4�� ��閏��_�>t3�ZM���[=*>�X�˯��i�o2�Q�>���� L��n����ɬ��
���TШ��|+6��u����2�? � 鵈Y�8MB���W �$��a�r��;gc$~�����Z���T�w-����hՊ��'Pr9T���=,公��*���Ż�c�{Ĺ�j��'�����}1��v�2|p�L~�4j_��"��'ޝ��v���G�V������(��Su� i��9ͼu06�+����窮����ͩ��7�H�G�Ѫ���S'n.~����=壠���gI����_��^z�h�ץ~?CQ�4��V:��d���>f�ldd4*�W̆cll�\��
8_��>ܙ��j��*}����|9䢸)b�ې�%�n���}H��c�a�ID�K��˯��}n��\�0Db��w�acLW6?��#���8���n5M�{ũ��UZ�F<��)�����M����B���� lP&5@r�CG�_��<�3����"0������e�!��O3f��Q��v���'c�������+]�KHw	���JwIww�,%  �)! � ---��R���{���˳��3��;����wD��mg����AM�g�Oՙ��%���l2��%�ph��F��
���A>��kw�h�.�F8ѽ@�p��rsqY�\[!�� l��X����U�0@%��e~��*>M���ی���V�|�}L!�����a�X�s���_�~g1gآ��b˛���|�l�W+O�Ϋ?_���"�g�W���,d�,�$��nN�G%B�e�2D0X�"�U;Ŝ����Q�d�t�����z�q��f�`��̪��!jC��nxbѽ!��T�z�A񽦏:�kNړw�����Z:Ե�l�z��9��̲�%��q�gDl��{����Hl��$��o�X��lX	h)7C�p��F ,��fd�֥ᚅ��tlhH��>�?�����xA�iI�B��!iz#¦��?�ĥ���N'��C����K�U�ݙ�q
�P���5_��"B�K@��t����Yl�'H�@�<���2k3��NP�9D]=����I�~hk�����6{0=���e��M江/��8���iliI����ؾ�yG�䛛���(+>��f�	�gʝ+�� �����/~�~K�qחܬF��\{i	�-��������R��+R7\{t_#1_wa�J���u+�/}6���f��� �{S\�	.��`�=�!#�a�������J=��Uq..� �9�kGI��1FR.�T��@/-!զ>,Ip�T�ڭy�%��\U����Rݵ��|��k�E�_6- �w���цRX~V��j�3�l.���'�z
��a�?6R���t��֗2F�_���T����U>�����v<
.6$�� S���Ve(���em�/�����ס��=��ȏ�d-2/;���-�I܆��w]��w]Ҩ�F��,����tp��>F��Q� 􎧫j��C�^����s/U��5���rW�- ����+�Jo���C;s��&2`�^�q��w:7�YV�{q1sr���T��%����L��RVR�g�"I*� ��J9�fbԣ��C�l�.���pf�sG,$�����U���xjx�TUU)g�s��~/,|խ��ah����J}�d�o��~�+}a�x��3��`){\��4�9Ч>Z��٥)��&9��ٓ7*)�Ad��U����k;���r"t�[��������N�+7ql��8�\kbZZZ^�DҚ��T ��]�C�ϼ������E��҆��*���z���e:�3R�����M� 1��.�_U:���Tc �:�@��H��"S��质c)����2��rP�,�ĳ#��DAP_ �
gFgh� \��V����v�����f0��p�9I�����"Vg�)\��#�C;O ��i_6y������՗;��
퍚�k���6�Ira�(�L�m��������E�L��M�1F>�.�_?㓄�-9h���ΰ��^�Xd�&���%�����)��+�kh�Ǹ��{>a��&��t���_��Wpb7g�LL(�弍<�9Ń��" ��?C
}ann�%@��s��}|�U�)�����^L*{�Pk:�={�l�n sy����Z�0m�����}�8��9�sqk
0%�8�]� tp�=΋�R��>'���uS������Y#�:�if)�7e��t�G��
Ȭ�P��ë&�$����x2^"""���}�!�'����+[�76S�Io����gq���9�,�VT(�G�/�WhT�7c��\ؠ}>u�����qr+����[Q�W���`��Ƥi:L�vk.M4cQ���<.//�C�JE��U�f?�7ߕ�X�]�3A��L��6��Z����� ^I@k��
�؁pe,Pֽ�,R�;^EI ����<;��\�T~ͯW6���F��0a��>��?���d&�''��ѶSE���~v���c�(4:���yI�;���WJJ����/����OI(��� \���s%>[��ʐ�sћ�ߩ�X��~¶����8�o�\e�o�t��1�i6V�(����>G�<qIj�~�[�L&�#����/��!�D�I�*�lQ�n�bE�|����_O~[ݾ��:tv����zeG���%}�y{�����љ��a�#S��O;��}$���{/�^�����2�+�2�x ^���r K.fdE���`��ݎ���sv}����v������~�*�e�W�!`��{? �墽�D�2n����C�.DW
p!��\/��~�I.�85��^�οWgCFO����V=�K��m�-��20pjE5��zX:w��pxޝ�ԗR��]��)Z����`�s��ڂ�}����k
��DL�9�)=�B�eH�,�yr���0T���}�ױ+�-2h��ɽ��ꎪ��T���|����@�q��e١"��d�C�0�0���˦A��¯ʆӹ�Ig ���W�ى�ܥ�8g��.�B:)����`9)�#�1b��kȸ^��M1#�@U�����}Z�� �!@#�N�[e¦V tKo��]u��_7�*�_��;��Ã�ش��z��
l�Q���*�ku��S����6&��2j�$��T���ퟑ�<Rm ��+��ל���G�;��(�KwKB��Y���!S��k�9W��@��?��� �L�a'
����o?d.��u����M�bb5NI�,�f��]����A�t1�� B���A�#�M~sU�J��щJf�Z��\�p��[ٓ,��6��}�cyٻƲ����ɄG튌R����8�Ю1?�@c'R�B��ͷ�-�v.�$�R�oe�
�#M����j�1� g^� ��r[I+w>C����Xʟ��'L	,f������\���Jz�Ә�Xz�]�@#Xj/e��O��Ǘ?�ҙ[����v�G���n�6O)j��" �-��6�%S	i/;U�O?KHhϴ���~_��TC�q��,u��)�1�2""��m�N\isl��&��� c+��� Mle̩�U{�G��ZC��a핁�z��L�pϣ�Lc�k���?�,���2q���WmSC��ȹ~���+��<�ח�OuQ�����bcF��~3-No��
X�q �46j;Ǩ6c�~ժ�+�K�&��<�i^�L�o�X��V�QN�N�彼�ˏ1��d��6zsk�U^*W� uȂ2e#0�F�����ί�/N�@��ؚ��ku�2g��Ź��lߗ'þx9�%l�%.� ��&��{����\eG뺹��55��|y���U�Xi|��It�2�2xT��S/��l�ԡp ?eh�����V/�>)ҙjxg�0��^)Lr����a�6n,e��ajd�����m���:�0�%r���Ӫ�B�ׇ���Q����0>�Ug*�]�Gx8w��O3n�̅U���6����tY�c�6��܂��=I�W�T�}6�x���0n��z2,����PB��1\[(Pd���do�>m�����ڧ���^ڮNcՄ?�~�Bh�kr6��\N�h��DC.N(��bKE�K�Gz�B�v���>k��3�i��.ߋ�r������wQ�fg�t�r�u/_�.|��K�1]��btbЃU�[�ű��Q�\GN��2�lR@!n�n�N˾�E�
�u~����َ_4��(C��D:7�%���i�7�{_h�!�ꫫ �_9��sg�i����܂�.��l�Z��&
�P�[/�s���-4���V���:���X�#��x��M�� ���CW���}eM1�D"�&c�.Pם�A�jE5�w?i��֥Z/'|T���ݿzVU����@���LiG�Ȟ-���J�y��(Yd���܌���#��u����C�D	��k#����fo����������T>�ǥt@�P��
y���t�od��H��	�I�9q<tXlX�~���Z��w�)p^j}���P��)�����c�Yy�Y�����q�����GElFz\!.�Y쯵M��?�^۵Q��'<���ja�T��[�N����(!����N�U�J��S�b2�?�A��$��rPDZ��k^A�����ȇj���~$�Ǘ��%��Z��E0�|N�i�f��u�m7y9�Nnd���f�fѶM�bKs��A%��ӭ����ә���a_h��|Z�5����ªr�)�X�{nL��q��G>���>���z�å��٩�jC\t��� .��N䁲mU�`�m�c��^�7�Ax�ʰ1F�+V� ���t�&��!�߁��;�4�������c~ۜ�q/��՞��.S���L����Lkˉ�&���h�AbnL�;��B�"1f��SI�ʊ�%��2dC�0�Wz��0�h	D�`P�?͓��DY���>�ލM]'-�y��~nW��w�8�i={E�'mZVn�;?f���	�h����MO'���Rn�C� ���M���烈V�dy�5����v���xs��j�s7×����ySC��'`����d�ȰQޘW� ��ݨ�_�������T�O:ukF��G��TB�C@~e�Zf�6M<D7�"�U��VV�&3��[�m�āB�n������k�~U��.��+��k����<�����.G���U�x�_[J�f|��-��d�Sֲ�x4}�m����AC,O_��#薷���������
r�I.R����
)n���{��|���W���R���r)3,�aK�}��-,,\[��3;���JX����3]S�����C��A'6)3h�G�o$��!O� ]FAn���0b#�!�ֱ"�;.qK�,/G�{K]zw�x����񦠽������|s#ʬqFҹE��ߙ�Q�������c	_b��=�F�>y��sbI��"�j���������*y0�eV_���h��EI�M����k�M��l��w�������t�5�y2ݛ�i��y��MJt�ȼ�c�-�PmG�n%����MG(�7H���.��|�3QП��20!�W'��z�*�$~�V�t*ţZ�c�έ��C��i�d�Z�B{�)�?�v�'F�un�q�[quyt��׾z��-&vl'�������3A����Q�FYIv��(��/L9��~�oe�~k{���+��J�9��Z��=s�`cf��#Q�໘���VԴ<Dn�����@��A�&ϖ�.�2Eɪ��2�pX�fB�n� =U9��30`�k�bӣ��I�M�
mY�Jl�q0+J�\���1�N�,��o���_�n���1V����	�z+�������յ��;�;��o���jS�~���|���ۿե0FP�U�8H#5��*�+.웦��>?L��U�'�X�P�p'�~��^�l�`�a,:����э�t0bL�%ڍze��u�ᬅ�u:�~g�&�osv�����OJ��]k�*J����W�3�!�v�ozooRw�4�����h���y}��"�]�J��I�ܖ����_���s,�����ϯc���@�\w��nWCA�������p�v�o�6d\�������y���9n'G���[��W�6Kq�X҉��[(;g^�,C�W�7S�D�Ǖ��8<�9MΔׯ��F��׮���$A�� �F
]S��:A�AA������C�7p�8lu��0��/ʝ�Ӝ���m�!�m%���=/>r�z(]�$���+Zt4���!�˭v��9�(_��"�� j'���-K�C��#Bd��%�!E͔�66������+����շ�(�ӀĨ�:����W�����w{0(�>H�d�X����u�g��Vp�"�X�Q��n��~ᇸ�7Y������Eױ�xf%J�8-���ʌ���[��0_��hjF�V�i�;�SQK)������S곥n�N�>����Yo*Ҳ�V���^w�����fʣi`��l�ӷ%~M{�?&��:�a9[�(��"ي�Y���/�mv�R�됈?G׺�;Ϣ �i�IS������_�*	�u�ѨtI/h⭸��Y���A����i�J<�����>{��i���*bZ��^�d����T	+���{��ǭI����!����6@���N����b���.��̨]�٨_�*�r�ӡ����C3AVR�ALB"�"�W�k�Bq���-N���=7�������H��>������`�X�H*���& �'묐��,V��l:�����g1@ӯ�>�L�)��7��E
��\}(i���"�?m�>J��E�������Ϯ?	���Ю��o�2JX��;��cG�e�[��}�/eǸ���y� =a��U7>D��\���M�R2�AP��Q�:����z����i��b��o�k�Q���]�/�%hZo2�'�	�#��P�::�����zg�.!��bL|߹������+����</�#H杆X-M�U<�b��#�w:�����y�̔���ұA���[.���z�T ʀ��!�)Ph��I���͹_G�:�_���2��Җ��r�\L�q�¹�����ti��� ��\f����x26_��U=8���M����
W�5H0����<j/�sw7���/o\�z��"@S�{�l�Ep�w�o�`_z�?.�}''�y�MV����e�D�'�5�c�t[���#Yޠ��pE�*A�\���>�*�Mb��J�[Z����hJ��R��Ф�maS�����.5��u�"=�x��+�k��~��y���s�D�$G�>���q�՟x�����)�Y�K� �*�l`�P_�����GG�c�b����.&���RZ2_~��bҁ�ןo&���r"+V���0VlM��$B*�E @I��y6��������j�:�l~�,�uj�=�M
��onlZ�rb��k�5���x/ut��!� �YV]*� ұ̿(Q�~a�G���B�9KO0��y%��G�7��c���󴍿}�G��/c޾#׆�h\PR^���E��z�<(C/ρ�i�2�Ą��:�]	 m�c��8F�ɗ)�-hN=i0�i�[+ס�F� W
�C�ÇM�:3+��hY0�*����D��'���l葨[���9�n�Pʒhfq�Q����B���F�4�WUUewx݁��LI2mU�!+Ө�U�I���Q�N�F�M�Mx+��S>֘j�<Jr�vر�����yb�=�����>0���a{$���%�������y�����m�q��-8�Y8't���yVә�
�ĳ�s��R=rkߖZ��dk���&<�M�RO������PVh
Ƒͧ��*ܭv'�Ҹ�q�Or�T�H�kxmԴ#}8W�^�r�ă�ӟeȐ��m�U�tM���=e1oJ��<�6���U��<HBǖ��\�h*Q2�t1*w��q�i��[��z�t5�W��?�v!"#��k7a���ph��{�.ET�i��Q���͹K�,���J���lU�)�u�~
v�[�~�x.KCşkП5
~����Z����BCμi��K�.���\	�g
 �)n�H�0oD���Q�ߕVW���[ $x�d��˨�)�(�y�: ���*s�{����w���y�g}8����6ț9�����ڨy�w�����Q
 �JNț-�e{WV$��-EmH!'�y3�k��]��&�w��0��6�ݥE�5�B.U0��;�F�����Ta�~�����l�1̄�ݖ��}Lm������,L��>��FfY	�e_՜y�ޓd8O's������3��0<��?���H��*(��R���zr���Dv{�9�]J��
�����g��͋,�[���TTTFӿ�J�T�X0`��'ؽ"��A� 2�ѕ���O��7Jv�I�+�]9K аW�v<����rDE�����E�����9M*�4{�.��4�ͯ��j���-�j����\���TwH����n�W�'ˇ�),��r�*=�d�-����N1�C������A{IHTԁ�ag��㱚�쿝ݪ�D���I�x0B�s^?	+�m;C��i�-�v]ۂ��qURv��֞Z���I�q� j�kFI�N����%k��n��|,�����j��ž�L�m	.,p���u�>��B�W�c�m$[k�P��FHĭ��ͽU��Q�����#.�Fw	Wo:�	y�e�8�dR�I���tU�ߙ\���
)��r�'��N�r 1__��+q�w�����n����I�OZ`�8��T@[��Qm��U����ܳ���@^��@�Z�h��
(gK?�YY�)x<\�蟫�i$�H���N�h}�j0��B`-�|&��_#�@s߉n�'�Q�|ci�d�E��a��ـ���6����\=;ˏF��]Ʈt�{���:5Ӷ(j9
�62u_��|'o��A 3Rc+U�*ALK�v��ZW8$�:g��y�^�У�bc������e3������Hbw��V\��<����f�V�F�d�bj��_/E�־��t ?j���<��l�p�tvC2�)l���b'�$��i=5+�#�zV���,�O_��7~��<���@�����.!��J ��W�w��1K�7^��]��$Q�A���è�!��a��X�i>'ʁA�b�/���b��~v��`n�c
Z2z�ۉ�3�7��x��F��1-"���.��#���R�8vF�o�L���&x|>��#��u��#���]�Ba%�����/�E�~�B��mx|�fM�/�!n!�{�.��fYN|1�� Xjm\�|���X)�G�%+�Z�啦�Y�5����C��7]�*�����B洐���	n�OF�f]H�z2��{���Y�W{��vo�Ӳ�;�QM$yɿ�+��iᖕ��%	-')�S��d������䌀����e:mS	POئ=��֡�z�%�NѺ�IE獯7�(q��6
��j	�پ��`J�>˔/z����*V*��j�g�m�L�/�=9
�O^}=~ާ�	��'��#�$�`�2�o�jS�B��?)���={��^��n8-��v�E]c�G��@"��f�4���_3�i"�?�c�Q�?LV]K� ?.���y#��v���y� �W
�ݰ�¬2��6|a^�lrg�݇&j�ؤu�å���ֱhJ���b��<K�k|Ǵ�ݐ��U�������H����_�b(�����C���5݁�R����a�;����s����W˳�M�*F��npS�N�p	��ōZ}���s�777�e�z6��x٭�S�\�hpk������s��TeM���m;!S�����n��%�v�V�h7�Ğ1@�ݥ����ڼ/,t����E�v� woK� p�(���wfx�FFC_^~���f�و?���ȱ��c�a�wԓ#k)�/K��YQ"\<�<�H{���=Z��|��kGʱ`���
s�]rx�7HĀϝ���>[�Ҿ�t^�3���J%��H�?}�G^�?�:+~�$�٢g��!��F��l���r�"9-GW�\�tP޼W?�oN$}�'�\��sa�oT=w�Nx�y���`���O�
+N�9Tf��y
c#���$C�lY�C&����U--.~��{~^����zQ�ٙ6���?�U?�;澥Mh��;��Wd����������χ���8XPW��@V�"��q�W�,�
��e^WdЧb�^�����-'.q˒�Q�E�����C�Ty�w��usUk�O �r�e{�jI�ln���WI�Lu^{��
/Z_B���|����ķKx�>10������RfB��U)J.��\$GEM+�;�c���/Ӛ_�,�Qa,��#:;67"6��Q����Xw���E�p� 3;o���w���uxJp��R�g��~>xH�"��5�A��������g�k@_ ?�.,����<������i��M�I7��JZ�l{�*�ho;��=΢���K� �^︈��v$؉>Ӻ���b�[��	��y�=aL�y_�y� �m��ݎo�Eٙ6���:⒂��IV����o����/���z��2�t�e�m��i�K�)��x���D�N�Q�r�/���Ȥq>���^53�;xk��2�:r#j�R�7~7��b��KW�63��14
o�B��������gYJ��=���Bӎ�f� �{֣�v�0+掮�&���n��$;q�,]R��Z�����\T>\0���qԔwB��~�7c$�ȵi��v���RUŦӏEKth��n�j�Z�E��V���YU�C	
lՇ쯥�A�N��y�p��^ui���F�� �hѮ�|i��w�� ����799��jF�>pf~
@�����G��:����Yh ���T�dsv"��,�AM��#@�������a� �B�!@�����_Ą�ȍ��?�2��QPx��S/�g�z"�Y������j������?j�|Fm��-ҳ1��ɞS�O���O�)Z��VՈ�W-�a��<��^��M�����W:^���N�ý)����*w�c���1>�G~3极�a]o4����y��*:��g)QҴ��U�d,�{�
��ٸ�981�&z	�.r����p��=�>!_��EVVV��:p��df�*�@�����]�߹�fj�c��*4H}�(
8��q#����X�����B˚��{�V�5���V�'ⶾ��\9cw��ݰpl�Ζ�"��L,b@shЛ.���a�6�b'��/+��"25;{󬥧'��]VZ*&%��Y�Ͽ��bgl���lhN�B'����-���m�oăZH�{{ӳm���|{��sssA�����:ȥ���c�O������y�d��GF(�h���'/�(,�2�zFF��}���Oh�a>��P�{��-�Ҿ��F�V�X����/W+ }�8����o�ɼ9{�V������Wo���>^��VO�b��վ�=ؽ+�.��DG`2��w{�=\���r������=^j�t�Jn685��%I����B`�w���ƥc�|�F[[3�FI*S�EP�����s<9>vXJ����;��n�R�Z3��VQ^����u�r����7�?BZ(Pv�1s��}V�e�.x�Qo���ʓR��B;����+~^%�t��e'�"���.����ղl�qʆU���R��-l�m�p؀[^B"��lK?�ލ��Y�
'S�7�{��b�w�鋮�D�k�t�ŬD�;�E�$w�'r����cհ�ue�n�E�K�0Ɍ�S��$ ����%�'��+~�Q�1�*��L. R	_�t=X��t��'���<r�O�5��6��5'ϑ�镈��!t� ꯳����e	x��B�t;�Δ�!�'ĥ���/J�0�(��.��V�^�u]$G�%��Dӯ�3�R�,(�G��vμ`"�IM�z�Y�)o(����;?��#�ؔF�8 p]p�`=��+]�s��t'T�w)�֝����"-N�c�Z(u����5�:�R�����H��i,���
H�Lќ�όjū�_��+���tR�)u'��ׂJN܍Z?f-�0y�{]�ƍ�N�ŶA��ϥ�=�!�C�Ą2�Ӹc h��ɢm�';�C@Ǉ3!@�n�V9�M�qs1���pɋ?#����9 ����#��?3��9�`��})���5�r�5"�+�o[0����P�VD��P��O0wƱ�UV�E��OM�<�LHQ��ٱgꐴ*�H(3aL�N������3�Y��Vi��,���|b_E���rN(�>���T� ������$�"��4�a������JU�Ik�Ͻ5� M��E��^���a�2^�:��YQ����>��G
dNbE�`hm�t�ɹf�n���33���7K�CO(!��_gu�R@����89��x��t����63����bY��?��v���$��jIZރiک�B�e5��Tߴ
���N���cӿ,�4��<,k��Ѡ
�2K1�.�����*�E�������Z�3�X���s��9�nڅ|���<�U���;�ῖ�L�⹗�'ʛV�\�Z�yr"��=�Ys7��_��,�z/�+�.L�˙U��kǥ���8���:��sLڿG��Էs��]Ъ�b����o�p��{V?���)S�_��F� ��鏌C��G��=��/���Kn�ĺ�'LK2�����JuS� �����6o[-�\�8	__����o��\�[}����_�aC��K'7��B��ӟX��^����k���n�9�YS3�o�'C�|����3R�Ny����D����\�?/mF���0��kƪ� �H��G�?o�8}�hYs�~�@������;�䋲�)]��V���f(;�L���.L
�L��+љm%�O�'�[
�f�Pd���3�7�%��-�j|Z�pP�;���NB{M����5]�]]�v��1�B:s7K����O�} ��[��3�q))<�o6�1@�"^����{UU����o�TYv���b�AX��I�ݔ ���m�,��E��_]]�
|>y~:�k��>#�����^�N�`t1�Q���;��M���8L7A�9\��'���"��T<�];��?"�\7����G3�" ��X�f;~Q�+|�(�DrE.I�q蛴���';�#���m�5G���!#n�B�u,�^4�wdACő�?��+9�5��{3%�`�����r�Wl`��\�X��x'�$%<{�=�9͎�rh�נ�Lc07��m��]|�s�g�?���,~G�)�E5���J��o�|*6V$������e�/Q�8J܆ۈˎ7Y���G�_+�hpQ���:6�O{�TJ����H�:��*�w��d�;j��je%Z��*b\X�Z�r���$�l��ں���˙�&םu�����b ��:���w�oq�àu�zn��w�M��HV�h+.�6K���j�'�؆��2/w޷B����+�"n�k�h�
ɒ���Wy@*^��6��e�f^�z	��˞k:g���a�5MҜ��� �]r�������v���,�SV V _��f�ɟ�G9m��U`�1H�Z��+R�=ר��	<=�Nδ����ԈS�Xwfnp�t&���b�n1ޭ��ǽ[�T�L�g%�w�����et�Ӗ.�?*P/�[1	�_]�x�ް[o;;(@�{�ӣ��irӎgeBgꋄ�z��S0^z@7�E��\�	�cEe�(�ۦ~v����2p�߹��w�Hx�����x�r���Z�m�|u�51_�М��XN<��6�D�W������I��O��>�\x��7��4ٓ���+5y���eNS�=ǠD9��I]k�6/��>$>�aKA����pNd�^�d�ݫ�rW�ap7?�]�4��W��\�V�J�aޙ&�)^D؆һe���h���7/67G]u��*6���DNQ��^������P��X��*I1Mȯ؃��l%X���99fc�nm������i��dӇR��ε=f=�'��c����U'�$X?]40���nB���$�6Mk�M8(�˘�--z?l笸�Z�[N�I gT��Îh<�ռo�@��B�+�?����|�ͿC�`��=@ ���X��&z����8���m����ʗ�LW�r=Vn(����^��{�t�����{6�*D̬%!�I��2�f�./l���q�uG����S�{�o�~��$��^ٶ�8�3�jO��HBz�8	��� SC���� �A#���y�q`�?ه���:�H�߫q��s���ެ�t�L,?��q�ux��ɭL��v����r��	7�R=d��8s�3��VP�"��<G��D(�����D�V���J~�ȣeI��k>C�����fI��Ģ���W��s[�HVQQ��WظU@�HJ�`�<4�C�O�e���sr��&˷����X���`�`�9�QI�`'�L�'6�(:ūx�p����H)�h�l��H(a��1�)�j�Ji�(��4���	l�Uz��>�i�ٝ �^7[��?m��\hp�AD?�z�J�qO�|DP_$�.���|��͢ Dү����UGA���GG�*���6�n���OJ���G��/σ�q�' (8���D�[ Õ�9��$�W���8�n�M^�� ��h�Ҹg��`ƣ���E�y����R�����7'�;�~8��J��k��@��Zq��E���_V8'H1?�?��O���<����=���8`�GJM<�4�Iy�'~Zz����8
~�MռfC�#\s2`*��4��^� ��9a�t,ײ�Y0�%	ɨ�
	�44�-Y���E�����ˬ����׵?3��4��IeJoX9����Q�+|��zT�Ĕ��Im��"u�e�~,D]��y ̄�*:\J�D]�X�w�&�[f�낥�ږcj����\ ��_-��AN��Q�CU�OG2��{D�Ű�[�~�?�F~'���� qQ���7푼�^�ItJ0*�F���n�2�or�Δ�5�H��v���KM�2�u�ެ�>=�f�����^iK��{� ��F����B����Imɡ0�v�Iy'GA_p�6�gI"_�1�h� �V���1���C&����)o�m�KaK��B'&���j�!J:�a���q<��k�M|�^E�pXs�	S�L�x��� ����Gyޔ3y}||�⋴� Ԙ��D�zL��9u�����z�e���1:$�*Nv5�8��G$���8.�M� d;5��ό�'����w�s6���cEtwg&�����X�It��ʥZ{�E���)W��5�Wx�J<R�׀/|M�<@ɓ|�J��?�n�)hJ��#L��:q�\�Fb
		y�͎&��7�SoK��i��P.���e�T�Eʟ��Jz���2�W)S��#{���������.��wG7��WD�,��脿��K&Q*����pU�����/{��DV_�V���/c�V�m�s�[e[�J?R�x�|Rܮ8QL`�:~c�������eF,��P�m��}���,5���٧I(��԰l35������|�� $��y�B����Ő.vTO��pM���%Dۘܽu��i�/)��{mf%�Kt������2[��U$Աk47zK��7>��
[�x�D����U�ζmϕ�"��c��IN{�&�S� !���x�����tC<@f�5�0)}1���"^|�h�Qp�u�3Y����j��e�ɰ�x��#��7�/1�����Şo��}V?�L�t�،o�M�E��4���ƀ��.q%{����-�{�Mn�Yx�d���daa�U>L�=!�DH�A��jw� ������m�?r�����gE�� 2��N�?�o^�����P>��v\�s(�@�/����꿆�"�7��E��N�qub�	���p@�����S���À�L�ynY;��b�B�7C�˛�\��&h!M���5A&_�EZ�]�^��1<-�0��*��q�Li/�rqY��91bt3�D���L�]ާme��5'�r�o�,�j��<�s�����|O�x6�b�'(��
�
*�\)��q��捞��3�����u��fI *��}Q��NS����7��|>M��]eb���B��.���7��.��mek����o����|�7j�"�\�E�Hej��˹����;;r�c�v��L���Sa���e�,�y�VO��
Z:��j�G��@,XԩN��F�f2��G�Vpa{�2҇��x:]�s�.�n��K'�,��*\A�)�<I�l��e���X�a�O=�LRp�k��
N��&����z7�c^%��s��vT#�,U���=��P��E����72�F�B��4���k�ҟ$H��d>�yrGv��JGt1���7�ӒV]|6]L�^��=6���V�y�x���)g~����6���Zv;�d�ξ��^,�T���w�r��3���j�l���������Eq��uSUi��(yi�-�T��0��J��۪�e��V4��@���V �ӑ.�!�L|���]hd�GLt�����T��U�Y��O�S3ss�<v�f��{iY7�����op�H�D�-�}�V��o�����9�ײ��m{d	o�aͮ�z���R���L�|z���!�o�嬿̷��2�<�A.�;�G���e��Q�X�,l �x�\�o:���31��e���� =g\���e�(o���Q,�s��:��=F
[y�7����D��H�U3]	�r��#��R"%:�ʯ'WT��L���|��KJd�o�n��x��ԏ��g�f<�� 7�K=���U:4,���|OAӝ%F��4T����4!1��c���0����yI�7����9��Ӣ̀+�`ڶ�pvRAL�K|���S���9K�W���O�U>��6����c)~dE-��Z\_V�ܹ����Ķ�� i{����~l���T��w)��V��0P�d�\Ī�f�:����>����S����}�ZVe��:n1f�9m#Ŕ�����bU�f�i��5��6�FH�0}���d��Ȃ�-��{�G2`�i鶨��Q���B�=�wfF��=#�Jxw����o�7ñ�{�+�r�f���E��"˻�f��6g�k�[�����e���:ؙ͑>��S1�H���d��d��9�e���z,  �%}�'�X�V�4$���^��#�Z�o�({?W�E�)(��s��#����Y���P�gV��'��"Ou׬����	�"�G��*,f{ܷ�4���Z�J&���({L�*�<����w|k�T��>���+�ʳ�'��!�5�'iiYR5��FG��S5.���V|#}�G4���$����ղ�`��"��7���wc�?��WGOz�T�8�7�h��k�h�e"9|��2�%����C���,/����˙}�P��^8h>6��?y,���Vo�z]���-Usþٹم��UL�Iǳ�f�~�1���^\���M�����O͢�ڳT��K�]�5ko�gP��Q�5k��Y{Kl����#FS[���������s�%O�{]����=&F�rw�W���1��zE�ש3�����ůL����b(:)o �?~���/�#�M��|�X�̾E3_����a���M򦎀)�]�O��ǵ���=���bu�r+�E*�竂&��ZN�O���E=����ZԀY�E��+sާQ*��wW�li�d48� <�(�.�n�V��K�i�_f�e"B����sK��o;̈w��A)ݷ��X�y���-v�pgW+;�t�� �N_�qW�˩���@��W��l49�<[*�\{�&|�L\�[��r�o@t����%�\z^��}�Nѭ��޽o)����b.m�g�������_H ��|X�0�ӳ�u	r�H�}ڤ���H�@�ԪR�P�s�猾!�{�mee奸 P��P�I|&-�{��t�K������[$X]J2��c�L�c�Ah�6jD���;�S�X7GLR�(Z���%��J�>� �DIOɣr_��m��&�t�p�m��{��p�K��Yt��y���Ǭ�������C]�v\C��O����7���l�mI}���>����������+�o�wH9�@���0������\��1��80��X�9�ep��eɝ�))1���C�
EƐ]v�gIk׾!�R���S��,)�L-(}���S�6~,�h�V�B���5ғ��D�hk��{~$;������?� �chL%���3y]�9@OImk����K��はƺ �[�C�զ�4�kO8?��F��䒝�G�#���0WD�s��O:�/_�KC���wc�&x�#�O�D���=��[��XR���4��,˩���F���8�*G�����߭f����3v�dԫ���E�K<�6P�=rXyR�pj�����~�+�*��Dr���H��ސ/�~�%��{�/W�#G�-���eˍ�׾�9.���u3W!���?�Pc�R@�`��>�w�$�G�g.V޽�,�ՂF���}ϝ����=N"��<�	Ęl��5���W���[��֫���ҷ�ҷ��Gla��q?0L�V��O)�e�D�6�6�l�{��A;�[A��Z�q��^[��*!�O���m��a4q�A_�J���Ń�����xS��K_>�y�ۈ�[�.a�fB
��u������R� �)X���k�L͢�f��!�9^}n�)�o���' xg�ܓ�H���ݮ�3Jy`q���j�;�Y	���t׆Q&��y�*�4���t'��O]s�v���jTK�Z�)G����x���M^0�������d�� �@;�sm� ��"�����@~���n��\L	��-�f��(���'�w�Zȋ��Ky���d��;y�c5�{9���s��n��(���Է�
Y���G���q��
��r��G�;��������È���"�d�4ܪ�6��-����CA�mg�Y�L}��8�?=�g�w�rb�n�?������!ſ�DOc�&�^�c���������K��Fw�]y��(�7�hD ����Q����#/���J��e�fzC�D�<���O?js9R������NZ��x5�H�U�7`����Y�E��Pb;���c,�܂l����6���d]�t=fh"�/��^J�K�^��WE��ӭ�7	(ڼ���c��%1�ED��Il\�Q�%=@Wƌ:۝Q��_4���w�C� c�������7�3h�(>&�wk�&it�����9�')Y56�e�kr:k��2�0{�Z����2X�������0q�z����\�+��+�[e�0s��3�������1{{�dG�����#i< ;��^)�Ο��a�=��e^ބ������T�����}*�G�����\�9-J� ��5	~�gg^��ꖐ��I&��{��5�+T�Nc���,�:#�����ߐE���)�;�$hU�����&�l�`��u%X�tv��,�D4U�vO~uJ����w�-uՠ�P�=�<�q�y͵��k��3$��Fw�s�!]�r��*M�4��']�{�7w��~��3��7˻����)A��:=D��N�F����-	X�u��.�ͭ�ՙ/���	=fe�����FΦ�H��]j?����"4�nD߉���n^{����ҫ�̊���-Y���|9�|�j	۸eHgb�qp]�ǞK`[�񘰏{"�,Rq�az]�P�W�r�>SӞ�ն�=��T�kV�,|gd6fh�3�؏�Pk������L+���-2JO8w<�?���VՊ�EׯOu�����,�o��^�Y�����x��gb�,`��R	��m)
Gʏ�/[�T�j3q1��<�R1 ��{��N*��2<b����C#\�v�b���6P&�{��Ml�ͨ�I[�y�ÌQ<��	�Z;0$�Ë�>�-S�̏�z�MWAз0,9����AT����RyeqO�����X©���[�DM>�~�iJ��/͏�J����_E��I���&�l�k���:��!��dy[b�	�l����:K��<&��	�>S�82y7o^�ǀbӃ�O����8`�⯼�mw��'\鈷M��?J�k��C�qIDႉ�^/D��Z|Q,���@t@I4��6����/�-�-j�b�PH�GH� ���m��]I)�!�7�&Y�P�9�%?&�6���_�^sD�B�ց���Y���IP`�5ϙsf��Zt�tT��
K4���V�E�����_COI����LؓWݿķ��������K��Q�� ���W�J9��<�Q�E����w#W$�0Y��_��Io���%��f�r�'�ZJ����a�6w�f�0���mE��G��r*���5,�K3a� �I�jI�:�N~OE�G�p�=�~QL��2럩\�I��∓��,�S�^����������q����)Q��&?j,�=l_�6�ʴ�����znd����6���S��U}�.h���A�gD�&��K�h[�*�4i[�nx�_aQ��\�b�M��f����q
�<x);�49���Z{;;������Yv*q�>�������`�tR(����-ۗ��]��|w#��r�D��Ƌh�z�+��R˃��g��XM�M��zd������2�M�{��)$��E ��_��u�J&c���)���lm�+k<��4]�nLm���8�����Fq���"E�ru%ƨʽ�r,j+ p�'e͸/^����j%�c�i���Q�[u��jn�ټ��*
��v���,���b�>R�;�)?$�VJY;���]�K�!�p��<[)ںg�0�vhE�9��H%JM�IyvQ 6Bio~��I��`�����Ɛ���hB�jBt�Z�9��������Xla;q�'��� ܿ;`�S]�Z�5�l�OF�_E)��;6�EZ-�8l�8lJ�>O�3�Y[CTy��m���n�㜺�\����mf��%���&��`[{r�	���ZcH	�6lw�+B��WO�~qJ2=��m���Y����d-�+�|���6��gk �2��Wo5��b
�N��>�e�zD�޷��	�z2k]$GB(�p�(Zy�����A�;b�N��-��M���ȢG}���?mjfDճDG(�g�|��*���͆9�Bx�Ф��������,��#�r^*7ϟ'F���PɵT���l͜iǜ{=}��j	��zH�����]`^��$�����6�쳡9wֱ��I��Z�j��N������IC�v}$��D�8N({��Tʿ�����1M�OV�Dg�xj���C�#���[���4M�}�n"ˎ�9�o����_�2I�iwgU���@V�+�L�{
��Cl���9�`�wb&(���wY!#@�`S��&��oU��稵܋�9�MD8��9Y�>ק��~Y�K�4$�ɏ'�|��ud��@�j�|y9�����'��j�|����z]��#+�s��%���p�����{�3LH)8'7.<���w��MEaH��E��#�O���%��ө?�k$�Y�-b61���w�W���.Κ�/^����i�2�7���P�:�~Z�Ml8�������F�1P%?�����v�y^�8����4�<%#�ՁTc��C��H0z����`|�t��yn���v��(���U_&�_��P�89��M)AT]��͠mu�oKc)j,Q�ц�����	�Q��ӗeP��rN����n���Y�HŨKu����"�N�g�n�=������(R���{�BV�>���"�F-��%*,��i�3�\ҩ�#j�f�js|��A�1���S(YU��T��(;�H,e���i��I���rXK�	=}�ۅo��;������>�1�
�5q=�N���mmjV�=� B�X���d@���ܽ{[>�EoR�.��2������?.�j`˸�S�WW�"g�o�����E������D�w�_�=�Uż�SURX�3Ȑ!�EA��!k�BX�ּ0����%�>���$�ro�F�^�j�6������Ĉ:��R�%1�F?�+�_�� d��8�{�W��v��Q�4O�Z��|�4�G�m<���Ttm��p	_�{��$W �_�Ú�������=���ublpxp��$��3�]~(�m�-90�
��g�Z�P�$j�dvihM�g��~0�! >����`� 	���L��!�V$�넂t�]��/��U��8#eέ�I"�w�!k���6=NBu�V��k�9WY��{���Ϧ�=����x2v� J��Ǆ�r�V������cL-͜T�$d=��NJ;Q�<ӻ�{HDt)W���Z��AU�Q�R�v�����l31p�v�w�s���:�q@q�q�g�Wq�m�HQ�4ۍR�X��6�g���[��kU�is����x��ں�I��;��_�r�&�iS�5%Y��a@���=�3���ɒ}��}�|�G��p�jy�&c��
�����!��\� 	\�.4�}E��I"�Uڑ�g�8L'P��`m�(���h�[\��ҽ܉U�Jd�.w�BF7Lc��'�#9��ߦ_��CzY���,����H�OJ.�|�d�7�񟱰j��`YI�в�wY�Z�أ@ړ�<�ǲ��˵�@��S�	u�c�*,��$Ļ���u��tl�>�/8�K9Yk!7=3S��4}���k�� mȊK�Jw� }��3ʹa2px�nk K\��_�[*��A@)%bx+��X�H9���0�׶r��'���	�v�V�g�y�;6<]�U�F}��e:}幋ژٍ�7������ᅌ�doЙ��^�~)�1��O��4z�N��yy�3��j:-GE����]{7���9i�c�xzFm�[Xa��d�1�gQV�V�������K��������V��H���*Ɛ���dGG��)��Z9�3JX�8��XT�Mވ�_��{��؉@_���R�eS���Íx���>�G�e�������L�^���߀�b]���c�R�m	�@4y[qܵ���m.��,r�e�YRƸ�5{���	 +C5%�-4�N�$��)��M�,��������r�Y�����)G�7No�(�j>zH�s�����+�S���]���}VH#X�}�������U/�B��!6ڠĮ��A>��
�~��7\��1E���ش�hS��z��ʝbl���.��I�+m˫�b��y��%-~��Y����E���g��3T�G��B�[���
K�~VW�w�V~w��e9n�O;6�3?赡���.�ʳ��EZ{��%6B��I�
m�T��߭��j|��p��\�=��o�=�������?%Ρz���'���N7J�72s�_%�I�,��B�U���>0�ͭd��ܪs!Ʈ��$��`̍,�����þ�����Kc�ƞj��@F��>j) ־01�^�I�*{��uB�~*�,��d���{l'b�m�(�
�\��Zx$�<��(�5�����+l�HxA�@�/B��N�%P���D�+�K���0ܣ�w4��1Q��@�*��XCc�'o�Xl{��e�'H�-{b����l��*Ч�|���1�PE�2��4��}���1��V�<Ixl�sK�B�N��f��Ϋ��l��VZη�)��S䄏���zY�0J�rp�HE��a�@3W��PG-e������̍�4R��|������K�͗Mz�J�WL����k��yIdI�6�%8��yLG���㇎�N���t����VT��`����A h�:����dzG�H�Ʈ���o�O�ctT���E��������c�$ ����ٕ��9�����Oδ��CQ����!�3c�)ᦔ?�4,��l�_����1N�;�Wa���*����G9��
� �K�Z�� +���a�Ff�PR,�{����b�V��Z�N;G���Y�C�k���J�W�������2qy�1��n2e��N�s:��:w�S� �ipFR�LAV.��<6W.����[�?&��\��`������HMF5�|��U�3�6צ�VzF�6*lny��������ݲ�����mf-� Ǟ3|&��(!�4��b�����19���Z/��%V�l�f�S��J<��ox&l�&�������@�h�I��m���z��3������~D��ʇZs�ն�,$:.Ȟ2�Fؗ ~�Q���EϣL�%
?|�c�IY�*�
t�c:+��pL�֛=5��Y+�2��m̹⣴5�����I�َi;����i�YN���t�ˣ�w��0E5�|�4�l�}����/�f��ۉ��^k@��e���W=�0!)���a3\�q�K��m*��)P����G����?����)>n=�l�ړ>#��|�Z@:\�5��<zQo�[[o���������3�n��>߶1�8C�P1W��{��'�)�꧗u���n*[��t��ɒ^l�Pͤ9�T���v��HF���hdq�"���Hŝ���Ǆ�X�Y�zLT��X$w{���P������vzW��|��5Z�k�p�����̷y��޷^��|����T����`���q	�M�ـ���ө����~����i�<�k[�-o�[�%)U����0Q�8/���D�iúT��4C��[�S���=D*Bb���4ǙJE!8XF;O���}o$��3=������~�$ 0�j�Ѻg��`l0����H�\�	6�5~(���mQ���b9������Իp���v��2���?�2+���D�P�������ׇڍ�����<e�Nk�FMѕ����W�9mY�#4�7��JID��$���G$�@�<|��ςXHi�ñ�W �+�=�r�S�$V/y-��O@b ˘��]]�|||ö�ey�Xi�V﷪�8�-Ȕ�?���'��A��qz�ܞ� m� ��H�g9~3��C0|�;?︑���6_o#t^ǥ���װ�JB'��kYw|ng�Ӱ����q�b2��+�D9��W�/��ĵ����j2Ϗ����5��u��b}����b8�^|�õ�Yҏ��!���`�L�%�d^�7h�;R��u�*�J�3�`� 0�KTH<�I3]Jސ��p~y�Q"s��/|���uN3�9���R�1��3�󖂄QV�A�gAf��9���r��4l� �m���u���1Q�4�*��,{vv��ef�dEk�&d�>)*h��/���2r$��oN�d<jN߻׍|$���>�	���R���<�nH95����`|��#�z�vɠ��49&��c"Ȋ
Yk#r�9�yx�|�uHXd��Ig|]y)��i����s3�y�4���YK�͍�E��t���������t�3O���Yn��N�@`�"���Y�U<��\�
_�#�
�	k^��]�#�	��>�X���U��pI��>���G�4�� èl;UT�)�u���́ܐ[aL������ˀ~�e�'fN"���s~��Z����kЌ~�V�����n����!k����0y��b���)?^y��y/aւ*�*_��u���~�Ǐ�¶iPU4>�Q-�Ӳ�|$F?�B�IvF��C�7B�<��Z�����y���,�Tl�yL����q�]�a4���'/|J�Pf�v��f'u�}b>V�#��c�����;�9���+�J�]�,�|�3�����nE������r�{���d3M�K=I���; DU�X4p,�H�%��p�%��]&��nH��������Y,�5Y!�� >�n��u�@�?F��������Gp�t�t|���
�H3<�g��9�����=#m.���0ki�+.�q�٭�&
%V��آ��������y�3K�)i��0 ��}�aE�)'7`,H�Y���`lBL�g<aB��Y��2 �|�G�!�D�����3:�����b7*Rf�:��G��������_}���_�`��=*P[�O����ł$8�x�v&]�fU&�5E9W��0˓r�睆���u^���*Η`�I����$� )>����OLO����n"��oɧ�$��V����_-G����6���`�r7�n��я=��?;��o�i\dX�!�J�Ci��R�ע��{�go�R􉖤��(c���ˎ����^��ї��i��N��)���[C(Dz�VΑ���:��E|�]N�e7�3�o� �j-�4�,g�,���r��%�>�!ĮEb$�BtŸ/nu��#o�Iu5;}������Ͻ�+�\�} d8$)᷏���,>'����u��DP̡٣/��0�ߝli�M%�qE���|y���^����E�t%<Yy��k���j��à��*�a(<�Z�PY�i�k�k6Ǥl*a��5�45b����c���8z�I释E�v���#�\���A�4Y���(���9�U�P��H�L��5�z����M`<��!.n�Y��*Z�6�1FX��<��>�8ī�����}o6�/�xG�@�<���la--Ͼ#��aE�[�w��u2��~���$�i:�_�������d��2GB�B�����Ga��5r�::sx<�<-� ��2!`=��0�
�����fJi���$UY�C�W�!�_;'d�%Ƭk�v�����>�.
u=�7@�)�w��e,�����_WW��K"��2ZSup���&��q�����u㶂.���5��Q5���+~T]]���#֚bG��7C"xa<���������w5�P����3��w�F����-i�������QǙ�\�l-��pI�=3tQ�Ym��{#AB��/^C�<�]Y�h.�)���Na�5H,+*�(/9s|��{0ę�~�9����X�N�n��Q)2��(�9��HܣL����i�n�K)����v�n��
O����wʛ(�Ȩ� e&�:�}I�b��o���I�y�����ǧ������k!�j�	�����m��zzFԙ�e��ތe�
�#���ϐKb�"�Y����?s��Xi��)lT`��c�L����>����F��߽5�D~��V�M6 �9}�8@U@��~4t�ˣ�6����k~�m��"��]̟�~��dd�tY|Ox��a�j\��Hc��p��aaq_�VV4y�W����}L�8��NM��u��_=��M>�F}�j�#Qŷ���e5�U��� ����c�Rw��"������n;6Dk�54��ǧ��h�.a�����j��qp��BS (v��$"����r�Ϛ�Z	i����@�c�My���HJ5��E�\�:?�s�Ւ��Q�����k
�#g�H޶$�r�B�J�E�{�<� =B��	G0T�#7J��V�~��k\�;7�q�/s5ʪo)mxYRѝf�~��z�C~',�D��=��C\�����/]�u|P Ui�&�B<O��E_eXׯ\X�#���GTB���_ǟ��E�����>~ �;	��]'@ 8�)��م$�����QR!�3,|�����ȴ��-�i��1�}�A.�Z��7:�f����}$�/�(~��%"&&'��V�����S� �$��q�J�,t�MWT�@�0\��LA�츃��pB�^!T=�Ri��ƣ��Ov0�Y"V�g>QVD�$y��n.�dJ$N�� eE�Id����JRT���V���������m��������Pס��[!0$؏hw���,՜w�g<����Fx{n���5��<��na���}V��g��FM�����q<$���I0�7\�eIf/���4�M�����6:){�eF̵{j��araw}�
���[�C�4%ae,n�b����U\U��S��lj�ʹƮBO#P��(�׷�p��_C��҆��~X�H>$>�w0UR+����7ײ��fB�A��#8��LM�p=G�Ɏ�˹�v�tęcE*n��-\�D�v�M\�'�f��E�"NKX0[�׶��W���A�
�����8{s�s'����=d���u�Y5T�ɼ����_�>�$$�uE{J�'4��*�L���R��
w;Z$��Ti��k�����"���������J�S�4qù���I�%>��<Y>=��秉~Sf29�jb��W���3������PV���Y�V��e&.�9�Αly��w���q��S��	�R����8v�e6Ggg%�ܨ�����7���j��)H���gy�!p73�7,�מKO�7)���p���Q-�g��h��f��heJ>�;G�8�e<(
�.Y8���q�ԣ-Kt@-�f^D��=b���yGC�nH�p�(���+�i?�Kౢ���xv1K|�u��Ǫ�G&dmQb���buY)?d�۰�J $yD���k�����L 1�aD'b���7%@���j�S�IGʗ鼽8d���zs�^�ʦ�XM��!���`D�G��p���?�"���������I0�M�\q°ޚ�H��|zMBL�rw˿j��M��j���I2�m'W��%W�5S�āc�Ń��b�˭d�wAA]�1�D����Յ���$�2V�~�����>�+l򁴧�`�-�83b�}�:E:��b�o�jBr2�KjNJ�I�fk�0�����k��$q��7WЮ�a���<)�b;̓떂W?�h�:�k;n��� �څ6�.,���ꡡ�i�O�OS�ƀM�t�H�(e�E�!�e�0�� ��؞(�c�u��_?F�W���~} ����U
(U���t<h���!}�o�]L>��mΛʫeSl��o�Jy������=���~�����0�|�s���W����\��x@�-.p�!S�&�o�?��u"W�q$��:5X>=징�ܱ����9\�Gy1�KdW$����*�+y���H����Q}��A�mc�zan5iX�_�.��*Q��I,�yr�sEg`�PI��LEi-d�:"��!>�G��a��Yu�vӬ�@6�$ğ�LCPo�ƚ�,�b�%�A<��6���Ϫ�_�ڽ���+�f���F~������^���$9/7�cb�p��w0��$^|��o�ʯ��U�U)��������*|M���԰R`:��@�������p�r�|+/
d��W[N(��-8�->U��̓����=MU�Zm���`6��h3"���ߴ�(���;��2���m�����n�Ғ�_7�6^��G�R�ɯI�X*� �(����'�D���i�9*Gu�"7�U�_R��)�LL�TAky8�zLF��<��DO�MekH�ݥ�r�N���c���޷��� [��v��"����4���D󐞓�}����ͩ��%�}P}���@<+��h�oi~�1��O>�����n`�����츥�����A�҉�y�����������!K�4Zs��J��u�K��9(M����߂��r=�`d��rX$1���A���0L*kq��Wi��I��?.�ݾ�$O�����Q^S�-�w��a��|\���~��O�ܢD�[�51E�<����t�O>�6�K�/�|ő����A�_oD�?��;	:��@�
�_fp��f�"β"@������*��@�2Pl��	�n\�F�RW�@A����@u���s����@�a$ڗ���+�S,�������!9�8�L��]��Ui�֘,!煛`�^A���f��j�sޅ�8$7)At쮕�1�g�L|��D����(��er��,[Pǽ���:�z��i_Qy�*6�Ւ��U�A������Õ��	8���y������ݽ�-b�v�A�᳃0�fd��0^FR���T�� I�,Kxo���WSGW�N5�a����ӫ�7��<7�w�&��v�c��/:��)buþ^y]����[�uY�Se�l�AQ��d[���+u���*}/ep.ф���#��u��Q���~t?䉡b��"����ص$�@LL������_�[���}u�ĝ���Zo�*(r輋-~���c`r�Α� �*}.y��`��cu
�Wy�QQ�c6Y�Q΃[�� ��B�����y2�h���=������K�7ڗ���.�A��2W�9!�8��؜��Y�UaR�y�xG����K�f�����C���6x�
X6�N���𗎟3�$�!r�ڹ��ٰ0+Z8�@YFo������Yq�э]���N�)7��;>��=�ᰭ�S?���U{���&� �v(��3:P�Z����y�B�dDܷ{w����h�<cγ�i�gP�;��z�/�=��&�L���N�IM.n�}�9$�����I:�kK���^�2{27[3 ��[a@Xϳ�'%q�)f{ЫG��t��H������(d������+dk��$��M�PV;K�|-�&�+��=�eRX����9(/s�I(��-�M���(5�b�$�����gm��J��y���Y�	���{�[1�묞|�zw����7��t`��d�D'z���nT���sP����(䣷����O���9-�V@�v��1��?��J��o��'�P�5W��[�%<rn=Ix�\�j�yPhR�ʸ���p�j��U�T)
�~8���V�;��p��N���8��/M����Y����|J�b8���E��}�/���<�J5i�r`ܺ��Ìn�w�����ٙ�����o�:jTX5���ʺU?�
�b~�ӛ�����$}��2K�P���o�Hʤ�/\�`&��V���^�V�	���#�ln.Oi����0���y��i��AQ]��s��O��>>�nKL��:S82� >>@599;�Ґ�ŦE��DH��/�r�^���U=��rZ����tduW��y�\�_xu��I�
 ��^7sw��γHyQ��iWC)�y��C6���Xo��U���)��4��4��i9��F[��7��gJP}0  �lFLK@���K���Ŧ�{�'�|�0�����/���K��Z��� ����k�S�Cڋ@�y�=���Y�)a�GJh�>��YW�Tt8Ւ~����2��"�d�̾��}�T�(>�[W)�Q��z���@h�ʳl|ʒ5�m?���W��i;+�+L���'�#���;��ѱ�w�k��<��eK�J�~�#D��U������`��jEz�ԉ7=F���`�a�5-��m����z)�"�e$7I?�b�#^�DQ�����W=m�����twS�)?����p)�\��W��.W!n���m��F&��Q��Pi�z��2vȜI���M�.�^E���y�;k�2;�-�5T�>� ޾X�u�t}�%����r�KUm�h�"�� �~�߽��.�@O��2Q,e��f��dtuu'7�=$t^��U�Ewne��,:���T����y����=�qyy��珬~p�PK��������n6�1�j�����,y&ae�����n����'�E�<q�,}��+=C��}�E�5�Ae7��dV��(�"�w��3�ԓ�I�}-��B���$́w0sM ���ť�I�-��Y`��1����mY@R]���1F*
�/!C�tSW��)���&;1b�A75�p�/aw�XD+��Sw����r1M�����}�л��]��������2���fg%VE�2��Č�u6��P2��ľ�Y�3�6�ȿ�.���--�R�ӳ���r�I�E	����J^����5��֜Ɋ��7bo����i-��c��$�/�S{�e�����e�F� 2eu�0����UL�wQ(p�U�x߇8ڮ���� �����=Q$����Y�&>�4����Ѥ��1��W��2�|k���2P*�ϜxW��o�����&��l׃F��Fy!<�U�x���<�A��[�ݢa(#/�=���m�hR�su
��ܺ���	�wy�
\��������������ؿR[:��W����pS����u~�I�EcP}w}�W�CTy��w��̥���;�g����ę׃�c����7m#g	:��>3��q���qp�{ú~|Q�g`�x��aSN^Y����Z��D�=3O5tƗ�1p�l����A4>2N��I� _��.4�L(Ɉ�x��(� ���?~����Pc'����
���4&�)>����ө�W�D��T�ި�XX\��F�d�?�PYɭ\��o;Z	J���$�p��� ޟ/�v��ۗ����7�V�se�_k��e�q��O2a��-Z�IB.�*�h��W�Sj�F���깈k�:�e�YM�|?K��Ǚ6�!��m�X�����:���
٨�Z_�����䮌��W��?b�����uE �=����������>dqwi$��ӏ���0�S\MMMk�?=rtq��)?��I[��<�#���bJG�ݯ:����:����'�s]g�E4Ka�����İj���0ʲn挶٫{~�	�L���-�x?�C~�
��dWȪ{����ۮwS&�����?n
tߵ�ܜ��3�����-�j�TE,�R�b/;ht\�����ቍ�ɯU��̺�����h����=��u�y��U&=��X�l��<#�"�XysA����⢠϶��RK�����Q��'*��I����|��1gG�'μ����\2JQz%dX}X������9Ba��d��Ӊ?2A�b��π���w�Y��5������ίts�b�*�,�C�5�&7y����9��0^\���8$��r�H��Y��p�}w����������C��0��I72i7}]����m����;�/�Q�V@<���s�|�(A5�Y�EJU��n�U� W.q�꿰r6r!��GL��ӒD/F����=֮�Jz%P�9�w�<��{|kz�CQY|���R��ԌA0�(��דp@nI�=��#�Y4�z��[\X��j߾���P_5�X��@1g��*������V�:�1��{���{`���R�եT"�%��[g"{�p�X:;� ��ʑ�}y�X��f�ig���Y�R�,�Q:_l-"�q���2�0�QPw3�kx�DP��pE�j=$�c�A�����V�M
��~6�lk�"�?���ૄ��z5�X�4�bè��x��&~ E�b9��t��>j8��q��x[Tx4���e&���N���(,����ř���z�w�����_Jz�%�[k�D���0�@"J�¶�۫@3����G�_C���ok��;R�<Uv��0����"�������o�;��K�b˔���Ge6�r��	]�Ɵ�T�V�<)�U���ys�������I'�>~�'?U�"*q,d1�Q��;��襶&��-`�'�2��S��*���˓�cYb�������6(�}�u�/w�3���{�
�q<��:����փ���3��'����u|���+��q�C�h��C+��^��aF�5��1��o��b�7 90��*,E��4H����s��L�K�����ɚ���WW��4�X���I6r.4c���%�GJT��H�"�!��.�d2�GOG�������h!�i��.�Q+�5ߦ����_�V���\���a�K�C]J,�M�B@��8H���*6���ai�0w���O7�Y�Y����3a�ڿ�c�$������Q��-�{GاG��;�J�Z��У)��]�XJ�e��9��1�"=7I���O���6�N�u �~��FH_6հ�ca6A��NLSaNLX�wX�����ᙊ��[p�1�J��t?��`�۳�n�r�@��bec��xQ_6��b�=$��ޗ�W�:ݱ,��hS���Ĝ=�煔�#UG�F�|��+���*˔S�r�s�	������C�u>�ACV���s42G�]!�@������bXQI�ո�G�p��sT{wY�붿�i�i��F����M3G�^�k(���>dt Ը�k�7�/��yB��@�*�AA"�d����TJP,��Ex/���5�4T�"�?��9��/�Eܒ�����t@�l
�vU��drׂ��9���C �q���S�D^���t��^�'��ys��s��x��)�Ƞ)�Xn���}q��p�D�B�t�RXFcSq�j	s$ff��g��5��L�N��i'H+j^�X�'a�s�X�=k�|P��V���.P˷?l�-%��*E���t��}h\\}�W�$}2��{�I	���c&�c�JaZ(/8��I��J��V�8��5g�N��=S����R+T��Ѧ	K��W��s@��h?&��s8I�]RR�β��i���5��Ȭ�^@"bo��G��d~&A��:ļ�*fT*������/�����i��w|��ʦJo�Ƕ���A?@G��F?�g�����F)�A͂�����w0C�H�ȟ��s&����
���A�$
�������������D��r�))鎡�!�D���n���aȗDbh�g�������b�<g��q�>�!b���<�.�
j�+xà�X4�z��|���Ց��񔡢\�Nzq���%t�>��lq�'f�x�f ��0O�� �i�6�o�wC�/���[;�lY�(�	96qk��h�w�V�ԚQjkk��D��w����]��a�/5�2�*��eI-6g܉�C��޴�&�T 9y��oz@�`l����,��;�Ux �*�#�4���",��f��:�1��┸[}�gрO ��P��<�ׯ_oNN�B�a-�"&�2dF����U�a�i��v���9��^LQ[��mc�R{�ʎ|N�&R�t�����莼c;8>�73��N��!ȇ2D���6ǧi�뽐��@��vM��i�3���O@U��ªnJ]2W.����1�G┈Z��ʧ]4�^f�q�A�qs��c�z��|�{��F�����~Ə�\����#�e��Z��ӛ�+*,S�o��D�h�{�G6���T_+k!�>�%���u"�o_��5��^w��G�ﯙ��ft0��ᬷu5�U�y~QY�]sä@8K�WϾ��SS۝��-Ɂ�u�;#t��):��?'�9���A$�z?k|tk��:8D,�!%Oâ�#q=�7���{,?ś��5d;���W_0[º/�����Tʺb�s�OaД*�ڹ�Vj-܎8n�o%���l�G:'K#�n��R�8�7qKȥ������b|#�hʮb���E��C�{�����D�(F�J��w�=I�-�V�g��5z{�d=���@���p�C�$�:�kM*��ӳy�U�3;��X��V�[Ikˇg�,��V�~|��hRw�N%���U���t�X(��d)qz�]����ﯶ6�ä�e�[�V�"7����������K�,�uM��/������3/����y�N�j�u�<�;�;�~��2T��<b�Oi>x�\ܷ���ЩT.��9�ևa���]��c�NFr5��yFR����Я��s���� �]ԡ�G�/��e����|��l�5�e�о�C[��x��3�#q5yz��H)��P������m���__*�� G���bQk���"��ۦ���ۮ�W�6��� �w�Q4����˄���D@�8�l�:A�( �����d5I��׎��y�R>�_\�ֆ��v ���G�S��G�N����1N�V;�+�x ��CO��N*2��-�/Z�<��!~�#���� d���N�=Y�k')�T4���ʨ)�yv�-ڜ��~S��\>;z�[Oc��>��{Q�VVi�hY]��.?x��	����c/�����bzp��Y���қ�Gp
��2�p=������̺�J������y@p	���=�.�M=+b >3fl��v�x�iS��˳C��S�rU ,��ryM��h�0����6QpL����.�p�g�B�܀����l��8��D�t
����uVwx��ąQz�W�&Z��e�V�MHݎw+��0#��QɎYU8\�_rC���5�N�v�������XY�Z����:���Y�4g��bU��t�Ϻ���V���뎔�%|eԖȐ����S2��bl̄�&�Ƨ��`w0�B��*(pY��>��6�y�<���D�@45g��~7v�w,K�4�I�o�4ug��l�8SI������Ò+��ۓ^ݗ���ʰ����y�~�yҚ yU�DT�<����+���'w>�θ2�E1���Dҷb$���!�qi dЅ�j؂�]������ @0��2�]4��4����i2����������<��x��#��Mq��¯��S� �<Ku�+��2�O|z0c�R�aݍA��pق\@�G_�w�E�"��(��#�9���ˈ�f�vߋ�������\0��i�� $3��>� 4�8w;N�<M�p��!��56��U8��' ���A��=�>��}�n!ө�����!y~�̗��>-,���L��b#���S�J&�ׯZ�%C�O����Qvoo/�/�f��}rH��Tzϊ���ZE+++A 
f�νƥ�|���3��ee��]�����>�5����dkqO���q4"�� m��Ԗ��N��,�;�Lǐ�gc����ž�-iLO�n��;��.�x�Ϟ�J)䉶��h�D.��|*��
ق�Ml��w�x1���4]�+h���P��
��e��g|��8�b�V@K��c��BJFƏ/νP�p��;4Wk/��\�zP�<$I`�.�~��Z(,��T.ڕK�����m�qHw�J�f�}J�������zI��v�h�`,�ϵŁ�����鯶���P��Dp/l��jBa��x����K}�󠎺�X��̔��Ψ>0�h�����Ȇ⧃���J�� �|�x�/B����y���i�o�2�e%��n\~����+��7b�Ý��S�b�"�AT�[x��z��l3_�]��U�c,EL9��含�+�!FB�^2� !R�u��h��R���GUx�^�s-�����z���`k�� 5�ݻc�Ť�eim���������<��;���� ��u��n��8�+�p|�Ǡ�G�)z�#w(�x��Qu��T0
K�cF�)�%��6�Uj.�½O
��m����Fh�ܤ3��(S�e��_��J�?����S�R�?���o��(�v���q�pѸټ�aP�^'��j(Gܦ��5׹yz��f���(�������^)_1f�&��-�8}��� ���(�d���j����;I�A�B��"A���C�=��q]�O� b���<��� �L��b��6�]��+�[~5 hFL�����0ДtVL��h]��t�L�ƾT�q�fb�zP_Ą���dk�|a&|b���lX�2jr���kc�WlD&�'嚚I �g@�Z�Y�2{67Rc����b�BԻ��kW��_���y��n�Q-��7=+���<|��c�&O�]��nc���/�W�f�m�ߘ�#�� |�[����6;f=��ͨ���^�ڽ�%��>�Uӏ}�����kF\�4�j��$�0H��bvB��O�Y��<`�r�z�\��o��Q����boH�q�&����z����][S,(ݻv��WQ,
,��V�`�c�� j)������(�-�KL`�)������+da�ɟ��^ʌ��j
�*0�X�����؞�	���t�j�����}����^~�u0`A���?�x�)?!����,2���L-n�s��~����ʠ�������M!u���p��4�!>��']�ܡC�~�����<kM����x��V���⺫�p5'�Pg�n�Gך������o�5w-0w�Ub	�y�' }	�d�f^  �޶&Y�.���Zrp��m'��4ߎ�{�VJ�)���aӟ�َ;�����k(<��@S��s�A�����eiq������/�L��S0��$���Q����+�����~`���h�����j�r�CY��Z<�I����M�A|s�ر'wD<�����	�B��-.}��� �k}\��Eײ�3r�1��9A
�i%Pr�Cvk��_*+�����1jM��S,� ��]�����&�*���0�3I���'+ʞ]FGSaf$�m���O��!
�� уK�)�՚;I�L[*-��Z���������>��>��\A:� ���<�ӱ�����_̙���+D uh�lPӇ�X+؀�$/U%
$�/x`�)Q�Y{a�B�Xr�����Z0�����Cd��m( �?1���X�3�*��n$|�G_G�n�3p�f�[������+���Y�F�%)$�z|8H�vz������ڱm��R��M(�?U���Zd�r6��M��H�{86c�u�3n�S �J.��~�i�tԱ4�\��~�M�=\dR�e���4sb`n��.�q�eVX��8Ľ"I�T��E�|�-��Y$@�9�.^�svR�o��b��Ӄ�n����wyء�/nұ�q�Ҿ�/,�<l������?k��pM�}Ou�'��،O���_�$��	�ĄT���L��>�w�j���B|����7�m���w�fN��ABޢ	)�g��p�UB�@蟎�/�懂�ޫO,���N'2ڡ����uĳ��"�G=����UR[��c\i�
�M��ɷLX	p��BESC�k�gxjQ���x4�
4��rm���֠��)twrF�ouځҒo�ڶ�˹=pw�$$\����X�g��~a��ݶ�{~ɳ@�zu���xx�d%J����_T+/'��t���q(}n�^hF�ߚ菐��AEW�N����C���A �S�\�촗A��M�,���.P�v�~����a�`= }>On�UG)Z,F��������颫�j�:N�UkNV���Vދ�-�jLȖl����y��W�,�M,*_��(�V�Q��˹�|� �)|z�L����39A��,��8�5浰.�{f������b��°��Gf�t������� � ��!��}B[��9��Y�}�ю�Fj�}� T&J<�>���eF��Hvn���қ�n>H�񤤭���,,<xz�����css'#�n:^��j������/YK�΅�7�r�$�8�+��	�sǑ�i�Sk={7��I�Å�����݃��T�	dr�� �|����� G�)��j�9���=�A���I�2�p���S��l���
H
߬����������!%%�tr���<?�^"�&���UJ�]t�Ӵ���o%�'�>nP!�{��5;�)e�d沾��Zd���,'J/�<�����H��f��p,�e���D���?�9��3LD�4/@ii{��{��=���NS�Ү���ni+:�CP�+3B�aJ���GW��5k����}*��>�>n�f�&� �@ؙ�7�&��7�.;s3���(���-��)��K��{�ʏ�Jl6g?M�$G(������.6B�������޽�Z�˨9�!	uC�����?=D�4�!�P1�,I��+�"������o�!��7Y6����Hpk���f�]����Y�1����%q���7�<�������a��Ǎ�Y'�ih�w��PmR��x����ڇ�"޲����/OV>�v��ۄ���W]3~����k�>�,��a��Tv�х"�_���V}-�L��o��-��Ϯ6�k�64��i���IV{'�S�H��X�,1[|����q�ę
�>_]�����ؠ�Mb؁$]���y���p��H���Z�N�D��!����ٶ�|�t�,*[Z����i�\������[�����Bi���4�H����Rfߐ���{�xwkPU��(Kx�33=�i?�-EE���+7��>�������ŕG܊�/K3�ﵓ�!�l\�K��S8A��H�1E�2`k�N����P7�')O��~�2��M9y��5kF>3www�4�u`zF�m�I��nrX��<��b��u��˴&p���l�kKQ£�b�����ǈ]</.N'��By�<~ǱX���.�D�.Az�ajP�e^E�u]X*�ǻ�k�p�m���ƕ��T�4�3����̨o��D�����f��\����!&ޟD�b��=e�+��m��.q��H>�˶�.9�C��X��������~P�\��ee��H���[���q,�"}A���X�T���aD_)yJ��2�򄠙$˔G&]����:���,�~u+���Ec(��6��Z\C��-����]��h��mw�g &���u_��?�-�h�N����i&���$�&�c�z�趁�v	z	���IA�CzN̪���#�hŴ�\���5m��c��?�������y�"��l��?�M��iQ=���
�ҭmG������ψ6]�.��5�m�� y��Wʆ�f�0�щ�����Q�"�V��̑� ������M�)��#8�9���x��X,����o���=��m߽=��D��o�G�<����`G�o�4:���z5��z�ˠb�7�q���?��4�P�\>��2�M���:Hi���u���~���mR�4l�'u��}L�!3��^u��5��_0KLC�)GSX��?��J�X����3=�F�&4���0D����>��̋·��>4�bjj�_���~W���C;k�$�V�fX�h,Ͼ�U���	��T�g������\���Bk{�*k�|�|�)��>�c���*u^ (W��b6�����*���,��7�|9m�q��p�wng�,}Ee���Vs�G��Ssf�]�¯����.£-��*+V
��l͙�V�pק�R�o��9_p�:8V]k��i`�_�t�h�����Z��6�6��r�'q�i��9�f�m�yͮ!''G,�J�5�´�Պzr�bG�b�,�;�f��Md�`Ɛ����{�o���	�B�d��Ԗo������� �����J"kب�4�j�>n�B�m�)Y�T�"AP,��pf�-�׎s2����6���̊L�=���P�,-~(Sj��b�{���6����6Yg=8ֱNX�~�&z՚���H�>���%]"1�2/�ǩ|���l��J"M�����2�ՍO>�*�@2}574~�J����?e��M9��L��'�OQCN�}?��{�Q��c��S@/1��sSw���U�hG���� ���j"��'�;R٢�<5��Q$���bV���6�l�V�k˒,�LԂW�w<O���f-�?�4�ާ�7��U���d�%�����'��K�3Z����p���Y�.{�z��d��Z�U�9�|�		yi>���}�f�u3��i���[��_L�0�g��4�}��.5xC�/n�Pvc�wz�0�� 
?\9>33c$�qC����s��r2&���&���^*GM�`���=(Ȟ�Nx�~�I"��uϏ;�O�t-��k0�)�o��lUIe�cqj�P{���
�Z�^�N@���]�#"{��J��^���II��<�/+w�U2џ{@	�Z�=����ry86�[@��r�o˥����>?}>��7�Dz{]u�>�}"�}E��}1�-^���G]PF�aO�0bڇ[m�w�S��@�3~��$�����=��KZ+,/��ơ1��k�K��%�QΈ��O�H��W��V>�ZIB -,�Q*����&�(X���O�gʭ��qOJRikk(=��� @mb!�%�5x
T˶�s��~<�1�� �ONQ5���/�����4��_�O�Ԥ�/c�>K!`4��K�����I�;���*� 	�[�06�P��2>T���~������%J�x�p�,{U?�9�˹�0T�'̬Z��Ɲ}݇-�PE���Ibo�L٣$흣���|Ez�*�ӈd����lr�K�8=��z����*�9+W��Ǿ���tJ0��J��97�
�?yVa�J��>��~���J�@<�'���@o[�9���/5�ڙ�d�)�����ٜ*���;MW��d�ɖ�f8��`V����~���&d� P:�}P�EW�oIg^JW��Tm紷ȝ��jw��J���P9��h�G� ;ڶ�R����3$��KrM�q��rw���o���]CR�ܲ}�q��Hgڇ��0�����Q���|�6��V�m�#i�&�Д_�� �������ֈ��y.*�x��W ,:��x������4��?�Q�v��L-H �;4S���13��^�r
]����m�XQ?���zZ�I��+Jy'c�
Lz����RcE�g5�J��`�K��B��1#����r��ܝ�Y:Ӌ?�:���w`΅�a8$]}��x�S���#�;�@�_�������� U=���eH�h�ˁ����UޢѴ`�'8�UԸs�	�h����x���r]�~Ⳇ�h����?�o�_T��*�J��?��w�&T~�4��3o���v(-�����F�w"��`E�׿3��Ux�g ���.���Sx#�d����������?UAu󻺠P�G��p���>��bg�ub�ay�A�n��q&�9�֤$#99��q)̟��v� �>j���I�P0ƛ�C�֪�4��h�$�Ѳ'冄?����Rw*�	/3/�Aġ���.�a�pRo6{7�4ٻ2�Ӝ�3v�4n���lW�DJ6�8T���um���ܚ�p������T�7f �E�T�%��m�� 쵱�s6���y<�r�/�S^O���$�yz���l��8��'6�N�����X��X+��
��3��9�UKU=��C���(d[��?�:�lI�"`%FBDJ������M[��]�����G�/�:�ū: I_YY��,̔�"����钿�J�X-��6桶���h����u%ahk�]PR,D�w�E���D�3��
#�Яa�O[��? �uYy܄-2~,��K!�&�̀���Tc?f���� �@�f~��X 8�P+W�ţ�E ��%�"�y�g�t�Re�`���B8�8��/���l���'��]�+�!|c8��q�N�����qE��x�ͺ�熕~�m���/ݖ�Þ?�8v���Ƶ�?_^�)l�-�Ɍr�i:.�灦|�
%�b��Y���i�P:�[ީ��SOce �\j{��~�ww�)J���f�j���֩��H�<�JP�M
��S����/5�����4�Շ�Wh%���̘�˿�譔2�J��P�퇅������������dw�f��v�4 ����0
�׼[��=`bKt�h���^K!.�nZ�<��ΑZ������G�8�>�k��:hW�z�L�X��lj���}�IL�i^Z.P���x�
k&f���w��ѐ22n���|?����F����y� �5j��"����FJT0�G�o����vH��%o�4�V����5���mv�(,��*D~~��l��R��?J�;3,[aI���W`8�C�G_.�/���99���랛��@;�`�ޓ��g�Oe���Wp��Hk���\*�R����`�s�/�|Z���,E��������t��&�5��ҌU��eZY�X���y�-�����~8v�ˎL��1�I�<�O�vx�b����
�������9Ҟ�mc�����$�@e�	NY}b2�j�'x��%�c�B�7	!͖g��C��k?��SF��~5��r��dQ�1̤ώn�G6��5��	��α�-���}������=�f���L<�dDwQH�g;�| Y� gE��FȀ�랒�����A�E����	JȜ��H��gsZ�v�u5o��W*�BQQ�@iC��~�h�;M��L��j��'�(ʱ�L�m3�PM��y��)Hdi(��|��ݖ�9�^|�5��h:\�l<�#�Fy�f�	n����A`��r�4�m"���[��Չ̦ ��ڟ�դr�\&�d�q��߆�d�J�:d+|�����D}ef�m�nF߉�4Sx�e�k?юK	f��.�p�^/�o�f��{�O�+��>�d0�������S���,���p��>�{=�}�d�.p�G��ǈ�d�j�`��;�RC�ZoY��Ⱦ}~id���9S�$��gÆ3�X��S֭�)J�M���j�!D sX��
���e?ra%֚�rC�j��$�ܨ(TE]]��M�,EL��O}�`��~(��͘j�&�C��G�?;��FFFJ�n^���&�`~�M�������m��.���m&�pl
�ϙ�!��q����<�y4����N<D���*p�k}�&�`,_(��O�����e ��3�9kaf��}��!5�le��;�O����{��g���GL����2���{�n�L"�X�'������SF6)���������F?"� �'�H��g����9���T#,m>��W�s��}��
�/��~��H|���o��3�^�r�������!4�0���!����~ȉ�Y�k��Yx~K'K<@92B�r-�.��Q��F&%�v4��!�GeoD��g��%@�z6�Q��I�p�8t�s�p�]��oN��֕��@@k�vZeR��7l��z �bس���!dT{�����$z!�;G�Ja��,��\Nґ��ȓ�9ʹ��.M�T&�.b�"PG��|e��j�2�4����g>���B>��)�\�O��DE`R��hq��B=A��_���Bx�Y=����d6�%�a��l�1���9[�ϛ?+7nm�Pw/�)�6�V!�}z.�p.T3Bdb�(����wf%F��'�|� צwe��i��!��Ԡ�O~3���T�����D�lދ������9����5,�-<ۘ�z�J`{(�j����V-~����r���h�т�t-r���$nn�������?��d���-����KH#M�wdt���-?���ƣ�J���F�B����������n�7z���`PD���ݖ�m7T�<�D��H�@c5Z#��Yn�[q�{c�u�<�h�Q��S+c�*Y�٥9��l;��y+W�q���;Ψ�W����4p�yzlj���4Ox�f������`n�H��v���l��ݼ��Va�~����7#!��WTW�=�g哸�w�0E����f�սGCUS���D�0٭�DV`�Q(��޿cfR~b^����$!ޏ�ݐ���ZE��Z��çT��_�{V�g��y))|ŝy	B �؀.�[n�H����0�&Ί��Ag�&[<����I��_����p�X;�ҷ�i��޹*���X�ER��x[�ww�êZ�U���/�S�Qs�=�}�e'�;�����`d�)��'k�;2|���
{;= '�ܐ��� ��|_��/n�	;��!�v�S�m�۵L��T�|V�AOO�y�5�Ao�]����yR����is��x)X.�;����Iݖ��m[�Iژy�%�ox�iA,��O$6s_=���?PⵃD��)��-f�9֧V<�������Ϛ���{\��vya���s��+ֆ��B��t����G;cHʋ�8�0P���L�澬�?.L@<��i-I�ψg8�Ho4;�<��"��>!l^,��kԆ����V"֧�r%���M^e%��l�s��@�P�*ە�(��p�/^���5e<��P8��¨	�-y���g�rh":����ù`�)���n�t����>;����	��
�Lx��C�-8v@6�X0��Fs�c���h���E��o�)� �˭�bh���ód�&�{/�m[ܑ�VΤ<�
��[#�缁J` ����w[��9�A��%�Z��)������\U|�l=5�uXE�م���. L��#יej��2�-��@�{���X?���=���lY�����[v�yr�]�dER����F�����������A�1��KYB�vvn�5�BRA ��ն��r8tߚ;T�wt�U��֝��ﵬ�H�Y�Z:�- l�>�V���	� ��o�rH�2�a*���6�A1�nB���w�Q 4	���q"���M��!�H��GI�q��<�����dF���0���>�	����o�;>ǣ`�ڙ^�
�՘�Dz8���؞2�����ل]�[��s����(�q�a2��0�͛(?۟	�4�JͰw(y��9#���l��|�H��@K�'�C6���3_�B�=:�j/�� l�6��Ī��8L�墹�Bn<�'Mp����Z�����@W�Jңy���`2,�雫�_�fun0[��Zb���M�Ok�^�a�&���˃봭{�l<b�Ŵu�!S���5C%�-.@A�dز����;���wU�5�t��]D�O��%h��n���|���ŷ��6�t_��s�gy�'�}!��O��Z[����e�m���v���T�{�X�YWzqDw�dCH� rRH�2:�&�k�OoK�i�?%#G���ZR ΁���^T�_w�X >�՟�]m�B'����A�1���m�s.�ؖ��߮�}WإdEH*��8�1��G�)�k�Z����b���f���K H�_&d�6���jB�ңp�Gz�^� �^q`�$g�'�Mk��� �r���\�=���[M��0~L�T|���߾��?�y���g_&����������_ݰ��ł�J��s��bo���E4���l�.�f�xJH���߿�"0 ]uJsVۖ5+7�Q��� ��o~��pH49����9{�1l�	'�\0�����ˇ�c��u+E���m�N�ި���9����#�F�����}A������k!K\���܋,�m��_�ҮP�4����׉��p��N��3��Û	Iw���Q�1hP�#��7@�q�!�58{�[d0�V��m��l��7ӗ$&��E���,Oo1�8��G��G�퇀��Bi�4d����U�����-�S
�4n�h�r�,�>�j�j+?.���3�5�_���Q� U׫���7�a���㶿��X]��纄�qb� ���V(��v!�����0NuNq��y��[Vsmk���]��fK-���Ai�!y��c\Kw��	��q(�)C27�vUD#&A��䎴&A��Ci�c|��7/#Ղ5S?�T-�#P	0t�z�����Z��b'����wó��[��=�}�����Ba�E�����l[���k8A�=_�<����U�z�oX��%��\ί����8c���T���M�<}�����F^��9���2��Ţ �7)ӂ��" ��1܋�q#���� T&%Q	1e���`"����AV�B��rIs �1�"�?��G�����^�bď<8�6�1�7�{5<���@��3�pl��S�wi��~���`�UCT��<�-�7<�O#P#��Av;x��mh��HN-�#N�߉i3�;�Q��.�M��^y�U�H>�w�x��R��=%C��F�n�GM�]�@LČ���i������T	��kS]�e�m��˰�x��̼�I9��k�Y��w��Inܤ۠��<�ÏSv������)E�G�����8�U�O�Y4R�=�0��h1��I�gD���*ӓ�~7���NNe�"�ŢG�����ai�i>d�cO�f��F�
����k��?dw��)��wҙ��^�lYg�FJ�<�)�Q�\��3{�7v��]���D"���N���mDp�DK�v���oɥ=>�l�V��cR}cm�i{���T��;@�A@���}�`�[���γ�n�)���m�����xvd�1cc���=\�X�GS$��N$��L`�-����ꞕP1e����@��9�҉�w�lM�u#2���"@�Y�ړ����6L�w"�jd�wGqo!Uߴ�'�!�1�S�E;d>tH��KT(�ò�w��2-e�Hc*����ӱ�K]\��R��\j3��?!=0���蔍 PYUf����!eO����ѳj&5s^�	>�䚵i�����|9_����w"����A�9/�����W�Xf��rk�Ȑ��P�-t���,+-������\w�b���ᆤ>R_��;�TY��;&^��g��V aA_n4���F��^͆�<ݑ�C�xN/�j"�ZO�����a�7�d �{���X�W��v�ݗ�
��2�����_"/<�X��I���Zy��G֬���I܁[��%�u��1�'�}��:o��;�u�8/}�B����2�����ǶXζ-H�,!�(֋N2 Ȑ�Y�QO}�c[�'��'<�A����; �y��Է�q>t}��[_m?O�?�/D��'y������g��\}� ]������[�;;������R$�$����M��PN^^_$#̴	O���4CĪRu�3���!�n�������,-��F�}�|5G}d�h*����ы�,S1L�M���=9A?l��Zr�@:@ԅ6�Ӂ	�X7U���Ȣ��߶0���i��[1�~���S���{�l	9b��Qxs�]Y�o.��ؗN��E�HU��
c�O ���`�j�D����\��op��H�\���
8�i���^JȰ��Vwx���*Wĥ��uTz���O��D��D0���
r޸���#V�e*[�z����%�#�c`�����R��"��^^���a�[��*)x�C�I�u�^n��E��r��'_��q��p8�F��(�kiz��Ť-Mlx�*���b�Y%��1P��m~V�߹XqfQ1��b��{`�f�{4�5%�4c���1�j�w��5>�?���͸JG�Kj���	+u��^�g�8)�Qp��dC�4���@
���s�H��wbh݇c,���5���Hx��e�q��e���RT)џ�Z��r�е��c�M�0���F�0�i[�l/�{.N\"���yL�����W�r�r�DvM���[Y�V^7+�V%({���`��t�;7[����Y���Gu]Xx~_-~�����BPkO�AIT�dW�H��`���{! |�FdN>�aX��[�~K��$�2�~{H�(ڹ&���1��啭���ᬇ�J:��4��5jZ�ռ|\B��(R˝S̴<�OKD�s�����C'�Y<e7[�칉���Э���#�_� �������L���p�e�����=H�q���B���81���<��טo���姅��{	��N��
����f����s�RxC�%>�c7�Cr���o9
w�d�����>�#u�����wq�q$�~��(fO�ӿ��f&|�[�L(\姼�I1SBM���^����T¡�P+R
��m瞆�$���f��mX�2�ۏ������ڭ��y�[S�v���c��<���j��ݣ	�j��%�g����V������Ϻ!��ng� 5��Wk�k��#m������m��2��_�H����@k�Jw�MU���������ar�KG�|�-g���C��3�W��Z�\_�.ӻ�8�p+�˄bvݗ(sh,��'��2��u7��}Qa����Ǻs'*"c�C���{d����iݷFYs�+wtFϪ��cSH�.�5�Ard��H8oՏ��-�����P&3��Ƴ�:�f���Y�Zw$�
���ʯ��7���yQ�:�Y��u|�U1�X]M�:333^��P��Y��b�������� ��r���@��O	Z�=�������gsV��̻���wLQ�!�l�[4�w������Պ���rG�k�
�9�wZ W��?�}2Z`7���m������G��A;9i�sy�� �<Cvٲi�E<�S�z>���������r�b)�{�v���M���\�zw��ث������w�)ģgfLl�q�~r��s������$����u�l��l�F��3F@�P��	����xj(���1�(��8���scL��ذ�Kӻ����o����[AV��rԤ�G�B"x�ݬn*˽�l=؀��˙�۟�F`#b���Đ\aGr��`-����m�j]�7���*�!�#���,�a$^Oޓe��{��#�>�|�֟<X-�&l�[&d�C�)Q=���������<��[�#�G5l/�%��u_��$��b��u�	_E�>��0NG�@y���T^�	 ��G�����_�8�(h�|AU�;�`P�pe��� ��c����WTVW[�c�!'k}ʞ���R�bB�����l �=����0k����?-����T��#��{�(\V�BO�L�rDmv���Vj'���j8��x�V
e甴��մ�ikk����X�2o�@��'&--�Ը�k�����f��|�i3Q�kQ:>9I0T�o��Mqͤ6��M�]��`t�:���'`D��{�ݺۖ�dc����f)��D��w������:�ķM2%<1Y"K�i�xu%�W�q�_��(r�ް7.�[%n�O����%����.�n�.)--�ا��tww/
�-!G�ُm#¹"_�P���@�o�M�B2ҰD�e�V~YT�<l������8	�	�lH��ɣRL�k>�#��Q"H8x55R�m���� < �
v���F.+~�F|mhh��@I�ώ.M�X^JQ�P�����!��[�ˏ�C���ߞB�=�(���@Sj����N�����e��e�ϗL��"]A��KjۄuU���O���M9l[�g��T�����Ӯ� '������N���l�Ŕgx���k�o�S�!c��%��}[�KD��vR�]��?��c�kM^�9����6�y$Wr=�s� r��"���f��(���ֳ���q���O� d��Bz�_�N�Pؘ)��3{���!p9�fe�~���y�HnU�w|1#`��64H�(�0�y��#�T?mr�c�/<r�V�����^S������4����G��V�76v�%T<#C�3���`bڇKn�2Qa ����A���ڠ������_�?C�@z�fEI�T��{G^�l��g��ð�c�y2n��h���^#��Pł�PR��jS�r<O< ��2b#w��x�H�\K��'s�.Ù�A;�u�A�7�C�bj��,Eb�;&�9㋡!oҡ5������P��ie%�6=�%;k���6�V��}��K%�=����F�{K���2����4oE=5 ��bU�b�J������|5�J.,�g��iZn�*��E�8�6�'E��Kw���񺯊�y�1 n��	Ӂ�o�Y�[��m������@ӿG,�j���H(�d���	�����'�t.n�(̏�� �Ni CF�佫cp���^��{�\Y�����?E|`��'���5 ���{NC����2#����a5�_��X��>�Е��\L
�Y���䁟���0��3 �����#�����E�^�$*Y��dG"#�!�^�5�e�-3���ŽQTv��u��݋�%����|?y�{����}�紶�����L)��@��}���)_}G	!1V�]��aT}�*��B�o�h�f%U�	��[�{�n�z�}���� hX����b�#no����/N3�x��ت�yf���Y�ѡ8	���C�Pc����$Dx������M��o�c��|���]�=�|#:� ��k��gX@Uz�^���K{:-j&C�]l�����2���Wz�uv��;ǖ��F��GM�w�3�a�V��IО�<jr��U�� ��Q�&�H����ʉ�;�����:Y�I}:4��.�&V��v]�>Oއ�|�kM)CQv�����0�LQ�����;�L{�Ho'E�1�}v�Q'��R="o6�o���@���965�����X1�)w�s������4�X)y~>���H#M� �a#Z�{T���ݱ��������\ej��o�d2�`k,W�o�S2�nS ؈�\&^�x��0zr�mv- =�������>�G��o���$,�ʗ�W�R�UÓ6I;���3��?��(����8�z�%Tr�������/.� g�0���z�!z�Q{�b����߶B�
�a0��$R��<R�?���^��rfM@�</9Y"��upk�r{?�u��'lx l}*��h��������l��ͿZ��� й������U*�J�\VB>��>=:jA�uZc�������VH��rU*�)T]uv��m���d���e��$ V�:�A��L_N��E��t����g�)Ũ��1{+�W����Lp���@=�<�ӧ5N�����M>�,���Gr5�5|,N�����)�ѣCؠxr4ؼrK��k�s����Y���b(4�9Z�&��$=R��/ �����$5SI���`�H����z�p�|l��|�C����ad��MLw��/��Y4�t�a��n{ƭ���l�\YYyj���!�S��uiD���~�E�+rFð��Ŧ�vC�x�O�n&�^ك�k�<F��!ە�ŧ���2�8�W��ʱ�([	�o���Q K��_���������o��E7dF2f{�_��j/D���K��k�����H����������#_{{���3m7R�����]*E�Jn���N%�|봢�����1Ye��\�����j����ż��\ΜNQ�T�z�:��HZ���"��|8`ux���xkn!�B������T~\�f��R���u�X˝�^��ca���F��r�E��'ޔ��t}q�����n��Q8R��#g,VF(�^$,�<� �4Q�o�;�&UHZ�T��7w�� �ew�{�����_P@f<愬"��&�
M����nx0�ϩ�Mj��C~4Ğ���Y-�&!/����������(3������V:�?����'##�4����FS�H�Y5�|�;�����4�GZ�=��AKѬ��fq=��p��Mg���m����̂����w��S� J�f��FU��7$�T����G-��1�dH��w��Y	��?0h����M8�}Y����k�E3�}΀H�{��e�a��Zy8���/�'�ݏp�W&�5?q[���Ƅ���̏��C̈́��18�wQH�|?̆����=������mf,,���̀��߆S���o �b	�2ĭ��|�<�s�%�򺣇z�U<�N��x� S͕���9~-�(���|P�P�2���<��2�L)��e��gG�s�&���u���Á�7��zx�I��lxI�&�R�P%B�@ ��Op�@HX�6-�u�߭��T��;fo�&�d1ᵲ�����T�99��jj@��� �W����h�p�R8��3���k�A���]t4k�Y!��� �O�5~F���?:AE�:P�I�Dn�ˑ6n�,����c�6����OcKcҔ'n:�G�H(���0��{&VV�̚��9i۾��z��l0$�i�����j��e��R��%�Q �Tߒ9y��L_��l��M��khHE|�x��:���"H;�Q)�	{�	��� �K�'M�^p��
��WZ�,ʍ���{�f��U�I��ݾ~�l�Q�"�A�q��555�2��3�\,��[3qR����~�J���ת�?�썿�����c�/�oB�L9�`��tM���Ǔ'F3x���U6��߶���9�K5��	ߕ������r��M�#�.�?�~��(0�}zu��I�P27H%�����[�Z��
b��sd�j��$���]$�R�n)�����7e-Q :l_:�u)İ#��ê�%c�*O��u�tݤµ yH���@=�A�`��!9.p���9���}d�F��8̈́��r���Қ�ZK�hE�"R��6>���=��Q���IKԳX���0eÊ���<;������(��)̸�݊#�î �v���|��@#�KQк��X�&U�\ ���t́��A��'� Z�:W_ʃ��Bz�.!zΗ��D���i�
�����������-;�۲*����x;n �UF�5~�KE�o����ej5�G��#h�8���K��Ck�;Wj!������X)oJ�����|�L���Rh+ε���)A��Tĩ.����%��U�O5�:Xɜ�V0_%��<��E��2	 � ��-���.&�8�5�`u�p�����'Ǵ���O�����2X���" �Lܬ�����a-���qeZė�t�
��f�����?��]���9c4�C~�Y�&��Q�k,`�U�]���u5��������|sO(�0�̣u�dLu��o����K�T��G,'q/��L�`	8�GQ�X5��Yy3����4 �	!g՞aV���?6�x�U��W�z#��J-M�ܾ���o�����'��{�YZ��coU�K�G�=�~QE�,��9�}P��%
�����"`7ic��@�H����X��I������}��"�5<��ώp,މN�nZ�
��7�����_i/܈c'n��LH��ĉ^�.�y�}��s���,��xLՃ&n�4[(�S����t=��L�/�AR��t��_MO�g�q�@��*4h�&B�4V�u΃z��K���UL�nIT������"⚪7���,���(kǌ�T�o���Q��x�D�+�� �[���(~g��G2b����յ�N,?�]�hH���L�
�y�ߦ�!Vf�{�$I��{;"�;Q�VA-�'¶:gZ�M�e��^Ҵ���A����pJ������μD����`��Ò�<�g(>N����$�rjt��V�ɛU���D*�y<����GOl�U��w�s���RW'!�?�UPi7�02�x�͓�2��`Em��c'O�'�~#���Kb,_��$�I�G�=K-��$%HeV��#8^|�z�2qs|a!�'EB�f��r�K�3c�iO<�6�����x��f��!�S�,����wg@�!(�i|��L~~(��+ajcEyl{ށg�'��6�Ȕd&R�`�G<i.~q�I	�H��\́`�$�QiR�������lȓ_�Y
�0L��Lv;J��^��,�iETZ�|T�L�DRU7�(���eZ
;�2����`��hV�����=�vy�X�{2�_�g�3�s,��g3��=8�1�̳h}b�̷�o��q�	��Injx�-��l��u���ý\�������23�5G m7�m��"n�CI���zY�-�L��l=�|���L�3���X�I M��|���_�K_��?�u<�u7���Pc��jB��z���Ǭm�^\4�6z�4챸���(����<a����5��~��,����X��$qw�	�8�}{P��t���r��ﻧd�"Ԃ����\Z��$�Y�M��K+,\s����UN���GQ����t̖�k�R4�{���q>��Nۺ��o.w�����/g�J�}�"�`�l��5��"��XR`�M@>
G�ZȔ�2|Zu��2�~�x�qOnE����H� ������ �n���n�K�S\e�}8��йo;g����/����Q�iė���B�bW������_h�<Xu0��a��>�͎1�)'w�U�?9k/J��uo 1m�9!�>k�T�ҥ#/,�=�*@ﮪ���YT��#|����d,2�4�ć�㻯�tJ�4Q�6d}�j��ɚ#�f���J���_
��}����Ļ8�y=�<�N��s�{���]U 4BG���5�%B����¥���N�Ъ_sM!U�.�-�<�-��惖��/��f�<�����B`��0�������$�\ ?�����`���^
�$#V�� �nҮ__���c�0�9h��O`�G�A�Ծ���x7��8�F��K3鍀�WX�!�3����Q��t��$gQ�X��՛.kj?��N?q �>�`��|R�n�!�	q'�i�$�E/��������InB�<����t����P�^?��͜�gΦ��Zz�4g�\:������T%��=�ׯ_w��~VŜ�}�3d$P0�_	�?�
O6�D�"B�ܺ�r�9�'�� ��eQ��2�IP��jKљf�;�����B@O�RF@��t$GKzմh^��ĠtSI4K÷�R!uW�lG:t��Qb�,�H�����E�jɎ�ߜ>ֽ�#�k1���0������}z/)H���	֣t�#���4�ʪԳ5���+V��[�[��Y]�n�{�ynՁ�(f��
���������
~������9�/�����������Ik��Y�Vn#�	�NG;�B�j��:kj�{8KFeg_4*R�Z�O�R+֫�P\�Ou�z_'5��MS߾����|����*`G/�<�dH��*�f����0�c
��(D�PM,x�� ��?�Eů��q�"b.���/?�/��L_.��-�a]�Kn���x�3�0�uE�;����UǤzAcu��P�<NJ�����x�����uȈE��5���@ӣ�&߶��)/�_m�B/�L�Ou���h�G�w'�� cF\#�w���%7=�h��s�,�V��᷇���x��� ު�>}]S� �L-�dm��oB�YQ��6�+Ϩ���=;ɜ��DznxAr���Tn�����Q|�~�0%�L$�i"�����5<6ܿ䢒A����Q�sx�G@������&�	?��.�ܬ�rZ)��?c>]LM`�TH)?��x�(OOO{���۹����]��N`�/P�P��L����z��t�xZ���Nr�������ѭ�ӏt=�WF�
����������i���l�����Χ^���݄ѭƶP�,�m���}�_�Vt5� C$sEggg��B�ѝc��t�lo,�;n&�j;!�Q.y��.�����x�Ŧ���˿�\������~��Le��\�fl�Ie���
���L35�oxo�C@ ޟ1,THS���X
:44�	��C{L\��*�A?�A;T�$�UO�S."r��9�X�_DD�G���g�J�,jb��I �����@-�I�柿3'%$���9o��ق.G�"k�UzB������,�1HI4/�\ #EG�����t��.�
w`v]��<Z��(���Q� ����3�d�!ӋO�L,��L�)7�ZCw��N�'�d�+j����E,�IԤ�hڸ���ߩ-�2Oی�����5Q��� i	���wn��w��}	�iqO����9��YGl��2&�R/(
-�%F6K+��Ow��pi�zh���i�1jo#0���J�����,���~�Լ�5 ZJ���b^�j^�5�.p��FłQ$oLy�$�m�3��(��J������V$�O�q�/^��E��-�:�q�� �Uø��)9��e��H���mU��,4U��s��6�)�t�mq�j�&ɣ>*^��u�����۽T�V�(�A�����,s��t]���#���HǄ�����5[�����)�QU�55貦~f�����䥉�~z4R�����56ˇ@eG
�&�4�`��*�����|?vω�.�Iï�b|l�b�VX��o����SJY������&�m��o��~6�O�~jGͰ6l�1�#�<5�Fޛ�@����d�r����d�F+]�aE�#����(�Ex���{�Y�i�����S�T����}�@
��g�Q��<�Q0%������Mu�9i�ң��8�	�����{T���t>�$�369>[��u�·s7�ڢҪv�J�n�6�F��L&��t��*����L8>���̲�J���q%������E�xhg�j�TU�8�jJ��n�p���ǜ�O[�8u�F�Lh8!q<J|�oh������3�	�c�P`J�W�r���߂ʩ��\�$T#y��I���g�*^)�UG�9::
���Rc�pû������N<�V�X�����.�Жz3������ls����2L��s�L�ۙo��ie������3S]�v�g�~�ネ�h��i~�La.���P�X
4�>��Jr��^B��l���V�����KR2�R�e�"�k�4|��֓������?]Y{��,�խ��p�C�$d/� 4Ie�Q�&�_k@�F��y�f��[Ԁ_�F�d��O�]��;� =��Z���J�Ye�?�AFq���'�J�����ᶚ�+I|�����������9Z�|$�)��2�p{��{��4.��+{A�U�(`�=�TA#zZ�k��S<��81s�C;��@'�o���p����唻��9�f�A2hl��)Lt�,�$�G���E��9b�_N��^S��b� ���3�"��7��,���hԈIO3_29��ie��x�x�V��_�3Po����x9��Ih��z�� Qt���+J�,g �F������^A���|��QQ-��Oh.�5uq�oƟ�l��f�sρ��"��{�YU�'%ț�$���"��W�{�w���|#[���W��g������֒w��^ک
)T�м���m��n�D(EEE���a�6�eS���`�[)?Y�ڑ��΋~���Z�.����
��]�q;��'���R3�w��[e«{K�/����̎�k'������=��nX�Y'��)
Ҵ�4��𑸲ݖh�����"B�N��>	� `鴋��vOV��
��t:��r��wQ.6���XR�nV�ۀ��tu,�6��-T��,E�o~��ݤ�3"�-H��INk@�ۤ#㶆�,�ptl=�\)�K��~��]L�Iw�8i�Ф)��ߣ#A%7��/��/y�%��'#�H"������c�x�R(h�G��rF��c^�
�v��}�rh����^��s9\3��E�����ǧ}��Xix(	��Z�{_��Y*p�YnC\_l�5���r�}�{bO@O��xv,�@�f&14��%�`�휑�xf�̋4<�q��f�%_sFǆ��+�@��\r:kr�����@9u�"hb�o-F[��82�y�$,�eO������'������Kz^O
���b�A�j���m��j��Q����)���~#a���j���	�aW�i^�C~��[v��:)]�����g_м؀=S�s:��v��sm=|v��:˰�1���$Y.T/�ʚ�$�L���1���P�ܟ��%,���:��弈#S͈�%K*�N� m�z��ƅ���*ynj�=���a���	7 l+(�_M�
r��a
��쭦f�ow��]6D��?~�!4%�+z�tW��7��(|>�`��DٳXPyx��5��/b�<��TM�R)"��6�,4��s��ˢyem9W]��y(�xj��ڙN�b�0�J���?4Uݛ����ʉ��; ���e�?-x�(��uwV
�;�"���V?
w_��0� ǻX�9�D� ��;�gl��G9�a�]��9��}���T�Q��؈����U8��ԮI �j�Fz�֞�ә�B���ŏ�M�	�[����]<z�5U�.���g�$\Z�6�r�N���#�g|}w��G��=�{��8����vfm�j�y�M�������?;�~螰��6u���M�}����7�Y2�55�_�)��y)�>܈;�1��9���H�ӛ&��~���ڇ�;��/�;�+[�V�a��)����Mm^��.�y�i1�8S��zы/�31�#�Q{�z(u�G�Xz�SW�;p>���j��V�k�:3���w~�����6%V�<L뜎�PE�����W]��g\w����ڕ�4�_���Qt��4�~K.���^n��
�M��֜��>�j�S!��n��/��66�+��0�6�~��ͨЊ�gN�?�
�>Ɲ��V�Y����^�ӤK��{F��5~�Thz[� �ޚ���5��?�dʄ�E~@	~	/̱Bs�0س�Cg"L8 ��0��D��_�������>�s�O�R�o%���Rh���.
��\O���0#�[l?(:���e��\�Po�^��a�s��'+Fؙ���t�&M�j5)֎���4��Qdd�O��5��@������Af�!�<w��{�E�Ab@�����N�����2��OA�'xL#B7�:��/���DU%&U��'�ʓ���R3�a�rm��ySn�M�TVTG0�cFz4���X���3��]�L���l-�l��ч'ːxY�뗽��K-񗩱�&�8��2H
�S1����܍ח�"g�k�(��jO$�ñb���0K��2��[2��w#�'s�v�~jj��dH/&��oUψ��]AAΆ��v_&>ϡ���F��E�F8�T�N�+	4���K�o��,j�w���A���ڽo�l*�]g�CRW����`��lPZF��DjI�`8:�O���=���Nqx�}|V��Ē�T=����s�O�"��C����T�����!O��������{2=f0����5�AL�PXe�4h���䌡i��qk���@�~v��(����¿p�9�D*�Ni����>����vR�j��ŧ��#πF.� M ���ﰓ4�A8q�YM�[=fN`04����j7�b�u��+st%w��Ή��a�,�O� ��-�[6|DY�+3�Q�5q�,%7%h+Z�Z$)��VF+�E'J����ܜm�=��\�;n��n9�"~��d�Pa0�W�3��G/J���4,}܉�m�3v)E��@:�9\5������+���=�ý~��)WTR����y�X�P��p�	ف��͈⟫��Y����6L��PQ���A�3(_�����|��z�JoGG�Fq����ؾ���>�@h���r�f����p��񈯷N?'o]�S�k�o"��㋾��=q� �5���o�@C�ߔ"Q?�߼�L+��}6z_s�7���]Ç�=?�c���$�ۗ쟡���Ѹ�P^�	L������v���G.%�^C[��������с���)rN��;U̖7��1�I@�M������O��l�e ��@��WAg�Qiy�6w��l���[�����S,��/�t���p�?������vG�5�r=jL+�7E��PX�hi�z�7��?��#̊=���� ]��<��g�^�_E
@�;��ڜ��Y�J�j{����?��3��0�9��Q�����XaFr��8�!���i�9y�<脦.J�&�j��I���A<t������B*��9�0�׭�\�.�$�����@�E��jOa�1��a���F�8��2�n��u���Cr�
�h|��"�����4Qo��b��鴷|��-�I��3�
	��9�:�S%E�"먽
D���Py�V�/*��4[2Ʌ�IZ���Ɵ�B�]��7�@�(VD0��JO�:��èW@e��2=��B��:�;Pi��zieUU����ݔ�kT5_çdR��݀��cbq��'��w�A���90��v�R�2z滑��i���K"V*��*�L6�������aᅲ�B�=�Ow���o����_���`�o��@v_ͻ��pW�,�g���o��|^L�@	� ���M�@�q:G�as�t�$�k�Qb�n$������1�Q�KjA�]a�k�w�n�U�$�6����@^ʓ�3�+�(��c���e��8�h���0k�Wu@��)��G�)����⃣�� Og����O`�2;I�����B-a�@�;����~y�)pyf�*4�����R�ՅH��,�K#��۵Z��{ӛ���z艆3�'LI��{_2G���\vn�K��b�>���@6�Lu3u�d�=he��#F�F���a��b���>��v�/�Ɓ�(����J���z���A�"4ͳ����#9����}T�v.����->G���w2�\�&�{t�uL�YI[����.6��ߦ	y���p j Ѱ�C���I��-�"\燓�^
{�(	��6�(�	��d�9$����o�)��#\�V�:vrh��R�x���tY�.)���.��1:� �RO۷��Q���go��X�	���.�&���iXM�i���*H����>y������V��`�?�IZ�}��	(<#��r��1��蠎�f:4��/X��7!����8���#�= h��ڂt �³�K �O���p�SP��WU��N\�g��S;�Q�V�+Z6��c��1�ѭ��m�vI�?k�����SJ��U�"d�C��+9�}��?�O|ٵ�Zc�|U!����RtB@L30$��J҃���_�%��9C�;� �G�l��V�M6�p �U~	֩� �Ӱ��O!������x���Xu#@<e5�0dXY#�9/�`{�`mS��ѱ1���\+��VX�6i_�n���Zu���l�02���X|�C�{η5.x�|�!cQ�*}S��w�6����
~��^��華ޞ᩸zś��4�G]�'���|N�<��b-�¨{ZA+��Ǥ���ۈy���w�5�ބ��#�a��к�h��2F'����!|}�g*ᄬ��S�]a ��߻!�&�l�	I{*���Y��j|?M��wE6C� 3"�������o\=���o`�n�>X�?%�+m�$��`mo���u�m�+\��s�
���eS#��ݰL�0��7 %m�j�(��UeH{���qr�:�r�,�b;�'t9�y���|b�St��'T7b�t_����|�G�h�����FՄ�D���{��-���� �8�����^��R{�z�9�#n�2��S+����m 
�b��昚U�/6!!$yoӾ���AM��|��������5U�uE_�����ݿ��7�$�3
1�A�F��"���l�s���G�*��(�K آ��M~���L�3PnAm���i���U���x���3�j��p��E�2��5��4� �*,h����D��A�,��L\�o����Q丈0�\�D�������G������%I9R��<����B>�_B� }����ʊ���g;��f��u!�����z�"j��7!�1X��^D�A˞ݻ,�}����������%�J�g�9īH��?Z<�ᤕ���ٻo���9� 3N/�h��M�#�P��� `�k��e��`�5�pERZ�������cF����Q>h�3�fq��6>>���}A�OK��

�K�>��*�A���4�7����z����Q�^'���dJB̠�A�4@�%Kѽ�q� �1���C��8�f=�w[�n��H�YvB^K����-r?��D@��O
�vU�V5t�|���D�k�M�2���� ��@5��9X� �w����8��jG7_��ϟ�Ƞ�L�/����
�v?�Uυ���7�>:�L�'�A��oZ��}A��9��1�~Sn���w��I8�8�?��I��!x}R�}�g��R����p��%�F��c�̗��9�yz������$빴i�뼻��?;Ȣ9�+,������8�z�������S�ف����Н���;�Z-�'U����.�L�O������:�]��H���=���nS!�� ϡ.%�}�¸K�36�k\����������f���݋��U�QG��^=8���.�WLjiu�r��������e:��jr#��m��x	E/�e��I?�1o��j{�\��]�x^* t����l(��
�g�gB�}�Ł��0��P��8ƭEa��Y_cJ�3��X��K�;A�R��R�2�>q� ���JZ����bVB]�2y�����TfEC7�2&>�\T��F�|{� ��`jq��ķ�٣ƿ}�v�5��#j*�(�#��b�-�+��R9P��l���`i��Reg:l����� ���23��{l���;s��ޠ��׽�vo<����@h�)��L䊓��IMS��Ͷ����{���߂��L�S�[��1$a�U�1@O/��ܥ*`�T|�V_��p7�i�D�)Y�x�,�l<y%l�b�R�]��CÃ�a#}�5tY��$�����o{���i:Aq_`�]8�=<=����Q6���_8y%9<��ʘN��J�'�7��B�?9�Ry\�f٘E�|^��BR�r�0F��]��z&�EC�)������I��>��z�(@Y�ZQ���զ�i�~�af"��`� ����G��"�z2����b,mii���ѕX�NA�/�ɣ���5���j�{����G�������;���&�����(Kq{��e�i�v��*OGդ $Ԑ2(F�mE�-,�L��J�s ��l��NIO�A��:��O'F��;v.{��$�@X7����N�T��d}�;p����{��� #�Y��~ۈ�Y�����W��򄽽=���ċʥe�*uU��aӚm�&Q�G��c�y)+,�����X��4���çt}�N���ko1�J�4Yo�w%���,^�$#a&{[��(���A��f�����\lԪ�1��Xh��n��b}@��U�f3mV|�_Ϙ� L��v�W�!�O|=(�9����T8��M�����d-7���A,c�M�(�'���G����V���i�	���zYa�4�XON%���tZmW�7RƬٮS���Db�155)�>�o �$�1�~��_��4>�-����Y�0�1��y�v�����T2.clz*âf�}�"/��D$-�צ��Β,&����B �k2�٧��u�5��(��CD�V�nu�P�匵$s��^3�}��l Ib����H<�Pw��9�ˤ��#++{ڇk!���#�����3m�˓�J������t,gj,�P(��"�"ot��dѲ�4~�Ī�S]�#}�8����6Ǩ��P{��7�e/i7#�ȭ���r���"̾p7g�!��������[КU����W^�ݐ���_bMT�Fݤ�s�Q�5�^����&	�rs8��I���~�s: u_C0]zoml�(M,�7���Ή�@��R&ۖ�A���3����6iw�_s��H���8�7G	%�	GA�m�!7���}�k��g��?�F_<7�T��5(�`�ױ�� �r!��-jb�P�-����b�5k�q�� ��{�@���#ص������v����Ol�VF"�z�R�\�zr��v�>S��m� n�bQ���H�QVR�����_aA���a���p�F��^��k����6{�u�fl���Oy��@ ��I� ��J�vM����z�2�ˎ���f��O�o�%�h�|�-
��<���� �W*"fl䇡��v��-�����o:8�L�^�x�kEP���a`~%���w�X|����n�] YYeV,)�`dW�e��d�G�}T��&&�:x�:o���ζ�Z�VF��X����ւ�`\C��{V{�#�
W��a����|s2��o�?�͜e�ǞZ�֎E���?:�!�K|_:���3���Ѐ8���+��r@*<Ԉ��\�g����qJd�����̈́�e�|�i��]���E�C?@0������.�W�E�5�p�59�g�����;O`�2 ����HZ�	�&���޹��#NV���L��53�����{�0c�M@_��&��2
?1�|��>�9BZ����Q��(	��_�|F��~h�����qv���]R`�Md�6���tu�9���a�Cg<x0>=����˜�@'!�!�q����">��'/����վp"y{��[-v��|vV��V:�x~v�Vz���ᶵ���I��x�!���|���Id �j�(��1,��`��	�̕���'�G�C3�s��&UgJx�d�9�v
��n���r_ٝl�]���`�&�A�E/�YY�T�� =�x�=�P����{�W�x)3����]�F��DUz�gD1�}Q��� �A�q��$��e�T5���`�n�����G�_������4N#`��p�l���FW4�y�H���ʕ��r�Rt�vo�I����^��[3t:ᙖ ��H��s��r��;w�߀ܓ�V�B*Ѯ����/n-���_$R����r�߇Ѻ(��P������:�ٟ�?�9��׾�u���eC-g!��,CAˋ�d��$ߨ��_9��������ҟ�yeX�����S�R��`s8�C�d���@�X�}Q�J<td�4~lv���w�vDD�KA�<Ţ��f�{������8�׎�O��&bV [�rE�x�����t��]�|��T��R�ّS���ۍ��g̑ņ����w�~��n�U�������␗^ק���
����!!}�_L���:��7�Rы^T6��4������Z��Ul�H��3��:����L��1�I�[\m�i#���Wؙd�+�lY[A�"�\����;(r�S��m�um��0Dk��P��B*k��0�>�2��4���i����rY�.�w�<[<?q�����O$M�Γ�y,Rx0O�r�li�Ǣfҭ�L3R���������2�l�*���.�ͦy�sK�@�^��;=>f��Lt:#W��gO��O/h��H\�Ǉ"#�a����K~;��Y�A���π���4����qu�Wƌ��8�#��ҳ�L�.��򰞰��;������	o��a�������L������y�G�/��:������)w������C�X��_��#����S�H#!t�K�De�X���ۖË}�g�#�
)�0�O��'�����sg�`Z�N-�b���^@��qF�FV�i���TA�E�)�;��]&��:8d������2���:=|�P�a�����<%�k� ů;qO6���RW�䱅~C��87�d���tz�����E��N㤃�rb-ڀ�ݾ[ħ0ź(�'&i�b+ٷ��~�c��������6�����"���aS�FiY�r��L�Qu�ޅ8�(�~���F�(��_�摟=���D+�ع�N�@�� �Do�2��q�s����eh���*dv@��4E�T��M�����HSG$�!����#B
����`��^�E�G�,�4�<����W�2����5�U�+�EX���1��on�p�+k�'p�:@7(�����a 3�q�&X�
�����#�o�V�mJw���9�%RL{��m�I.1��_��"_[8uX�ފ���X/-���!�qG?�w.�Y�]y�,����y�߲�ܢ�E��]~MG"�\���f^��/-<ͭ�d��������/�~9�K�{
���t�G����^�B�+�ʺ��$��3�V
{�����sp9�
*=�iYρ�mH;Z���C���b��V��K7��A��p���unh�KŲ~_b5۴@�_����x����2�L�i�hdL4)����.�Ҡy�`�~R$��#�x�Ъ0�޸ދ%�|I�mP�97��+��2U����*oU�O��+IG��W�(��.�I:��ڠ�-���m2�xw���K�k�T�PK�%��
�	����T����߫�q��o\�ɽ�f.����	AD+8���}�f�p�������`�;I��a�(�#f�LIyc���)"�P��U�HS����|��ye�L�G"Ie�r_��ϵ˱���]∬��{���6�ٌ>(T�E����5���l��)��P��h���.W��c��1��%���T)�;��o��d��a��'AVVB��פ�՗F**=�8������V���T��.�f+U�d.׫
ٮ1t9
7�j�)���Vʖ�<*��z�[�����O��}~�1�xl�C?_�Y�}#�W��M�8�ڠ,z_��2�r�����]�6�h7�ͳ���O��/��l�t55�Q)���R���'Of�D�<��=O��H}�6;�Q@�+�WR[�	Qe<�_m;��:!݇a��2�Nvg{w�-Y��?�v��M����
�H�di�y�!�=�+�4�a�|���� ���l�m$T��G>��! �qI7�(�=~[@B�B�i�H��Yc�Ļ�߸1�"}�������<�!@�Ȅ

\l�Vw��`@mg��z&��$%κ�@D�ypv�����k�wZ�ʠb�zA���<���_�7���>�{mG;��_.w�_� ����"�)l��.l�X��Ue�� �4%�)�v����;�=��0Rtk5�=UI7Ҿ�`N�����C���߈����B���}7-����<&�^������ưGZ�bC7�L#ֺi��G�t�rE�R]�m,�	Rc�QjX�Mqq%-�B�A��*(P�C&�F�jy��P�Օ�Kyvē���qp:<2kӾ�uWSݷuc)��}l�ʡ������L��WS��T/S*��t
~�#-|���Bgn��7� �鎬?Eȏ	>hv��Y�.���/,�\@�4�=���VNrWٛ��}�Z06^��"?=�J�ES�j"_��v�;�J󬒯M���=�$_�?��2.�����H*)�  "�4(!"��tww#!
�]�!�"�tIC�0t�мg�����?q����k���y,�/��}H����(׻�F_�	�(���[%��j��i�w���6�K ��9�l�5��
Vl}7O�	��M#١�բG�.��B�7�Z��&�ܔ�P�M\NO�^�y세��cb >(����a�iKr���c�&�|R��<>u��h-z/?�0�ƥ��H��mh���N4i��0�C%����fA�7�F s�7�~�	���{{ ^���I;����� s�ϕ�٣y���_��(�\�Xk�rP,$��F����E��XZ?9_+�t��=�wh7!k�V�\*��ƻ4����2yy!.����v��J����� �k�~yz7���
���W��W���"&9�	84l�Wо�Sw�RahO=:hyT=��>�\�PP����ۓqk���#�N$��,z;�����2-8(.� :SG�/�3g�V�=%�89��V��۫�\�'G$툔��5e�������Xqp�͌Z�y�����#.�����__�^�U�w��<�´n"/eJ�y	.��WT�.y���TÃA��[�Y�������w��l�Op��t�1���D�#��\�X����×р�+P�/����N'�j(b��,�Գ՚|Q���Jn��*��o�)�I^\6K�)�z?c�d������UҢb�Y�ݩO<��)ݟfo�%�Ū�chw;��.
E��*TƇBH�0�`��[(,|Dh��)Ƌ s[�~�gwI����MS�K��u�q�0�$jw�ƿ�+�Dq<��o�b� �b��}����M���+Coۓ-�[�o�,^ʮ!ŏ:�� �c���eg�H��+}vnSvyhb��3 �?��U%J���1~�.T� \���E%�3.!��c)�|��/�Hlkk��I��S�+����?��(��V��]��'��S�T�P����A��XH7Vd��8��-۬T��7�w�/��HO���F�սf��q1A���#rl�ww��#�J��r��WY�)8��Av�&���'�nxm'��f���Yoc2׺Z|�E2��c��&>�d2뵶I@�B���zMx�u���b^���a;�a��=/��|qg�?[��л�?�}<�U�b�v���xR�O��c4�.�!�5��Z���*s~�H�[�it�!v�2rw��=�s����w�w�A"�)ɞW���>�`�I>�R�
u�_���BŨ��G Ǥ���k�쯂��A�ё#��-�4 ��4�8\i���sMZV��fSA�!�BI�N������3q�)�!�2���	��9���G �>4���ٴ0�cZ�o�y2�)"��$���7w�j.��͌gaf�1�jE6혍�����97����}-�����J��ە�|�I2�J,��2�_TU;��ln��X-I��ig�>�nO���l̮9������7!��:����_��%�z�Mv/Mh/P�Гm����gS>v<�\0��G`T4P4�I�����]�U�c=��'���>ĭ�0Kg_�)���XiM����0c�IN�&��M8R�"ᩛMi]��ք��:P�4cu�yM�A
�\�v� w���Լ������l�ݛMk��w�I��;*�������H������̵&����A_d&_f7K���7p������J��)$�T�^���~�cM	��}�B���$�41@��*�������XiݿD�SK�M��0�D#aVeZi�w�΁���E�&��"��0������,�/
|u6zA�ue� w������+�P�;"|�ڿR�4��a;�q��tj��렼���-�w3__��0Xκc���c��~H�.���:ǵ���n���]]n�Z[]�n���~��K�{���Q+�_z��1�q���M9����Sa����8"n[�Sz�6��P��J���0�u�(Q�;!�	4nݪ�x��J�&�s�b�o�c�G�QU �a���I�ӟ��EU0�'�������ڠ�Cv"'_ĥ^d~0��p���?K%7\�����m��N���Tk�ݜ��i+�d�^��]'��@FLճ�3Nԏjq�-��6m����RT��z�-SO�@^p�,���ߤ�?��͌pY���5U�Bo<�ь�$2�[b��-?�B��1Ԛ�_���I?,�W�ǜf�&ă㸺���g.�`�춸��1�m�kW�����M����O�<�]��5��@ѤL��*�h�I���$g��ۡ��|h
�DG�ڒ��f��w��h��Z�b��x�k��S��	`م�`�]t���#�w*�?��/v-�Kdo���a��š;p��*g(����]�;C��K�-Jc�6���07�:}�����l�~���6�w��Y+Ռj���qU��t5>�e���q_X���h�����	ƌ���EEɺ���Q[Ҭ�`fz�	���w}�AN��b3l���X�uI�φ"7fZ�����R!�P���泫�Ĉ��4�K��+Ֆ:-����W��8-Yl�?�dϽ���D��g	��;���Ѝ{�gG`��2�mx�j��6�~�@QE�?/���&�ⱒ���t����
X��}(2�+��'�w�^�w�
����T��q�r�g��N�������J�T��a��9v��#�������P��g�=�ls=��2�K��d2�кm��O逆�\oj��v�����N�]����b�YL��H�a��]ɡ9�fC��ji}<��-�}��n���<��� ���[�~p��y?�c�qDw�2��Y�9d�/���I�����Af��&��i�;�b��o�n2��F���8w�.�uz<�ă�s�Dc���VPIT�(���v��'?C��V�{C0���pǯ���e��n+��jF�T;F�y4�X�خ��꽁X�T{�������i�/w�N2���@�,�K 8Ӧ�PG!���|z�)f�|.\w�k���5���:�q �-�R�{��o�c��I���������l�r%���Μ��~��!���{=��d��߳k>����:7��BI�f4ޓ�,VCP �����^�}�	/�� ��'��q9���j����G�@I����{W��������A�����~�O�wA���;<
ȱXKn�"�b���3��H,�W�1��Aι\��:e������G�v#�WC��u2��xs�N>Eo��ѐ�7A{-���;�"���Fyǝ�n)��6"3����#eNP۟����/��r�4���&:{B��*S�־�V%]�.��VG��	�8�(d'�ⱹ�xY�@I�p'���ł����w���%E}ݣ�i_D8_�k�31�,��{H3Vf
�.q����@�so�Pg�?ͅP����;~��Nm�%�V�Q&%��C��~;t��T����`�SX��=8X��X\܆�H��N�[W��[*�O��С�K5�S�!�o��_8cH�w�a�G����ةy�n��zS�@Y�.!�ev�����'��%���O���`�ѴiEĖ��9+��ׁB�5A�z���Mv<��?f��aU\�E��cmy4��{�؏w�%.�h����#��ė.����f���M�!�M�F=�o�;�t�9ų��o�om�j��E)"�o*3�oXb�)�A{��MP@I� ��Ր��6~�n+��\sF����0�-"�������e��-7����N]��j)�i�j�Ð�*��P����K�cw]o=�{P	��g�B��ա��w�0�6JsH#�[�+):�XR�QZ�P��`��snNJ�{E4n�O��%l��M}hR����NB���ǉu�ƿ�;�Ny?Rk6a2��E�pDJS�l�]_����c��O�����Pf�^۶\2}[��1W�*�l��i������z��4^�Ȝ}��겓��q��>��yi�����@�}?%0�۷o�Dh�8��M}u�Y?��5��#E��..�]��H�XXDD&�牄ᅬ,�T�������J�`�|v\�;kp��ڜ[���m2�?�0�4������Z������Bɚ�5���h�����Dt�S��C�B�*E�O��#�����ɛ�q���k� Do��q��)�(C/mB$��	i�JeC���;d�*jt��Q�1N����t��nbM��Ij�����r�DA�辻|w��0<���aə1{�J�q��@�| ����̙�c����0m���:I��2��`GH�>�|�S~4�PG K؆=%���<�{�ԡ�������5Bb��z���d�\
,���*�c�7�h���8�E�ߓnj��m��Ą���N0^�ȅIܴ�u����'��{!�2|wli��Կ��v��cH����g�9�(������f�5S��V�!�ʱƈ����N_�ҋ&M��= 3��ʦ���%����c�!|�����������8���js�����{��-X=����NM(w]�&�]��t�%:�.��[�9�7�Vn�P������x��?�����r��Ǧ��wV�^���U�@�+�.W4[��(��3�j�,0<"<vi��#o;��tn����FAv���2��7�@�78^o�Ra����\��(t��D�Ol�mJ4�ҵ���b�?�QV�L��;��[ئaji0�)M�
�tjK���f?8s4Й�5�G&�>�6{dkk����K�ݬ���7�r�@!�9�O�+��b �8y�����X@�&˴�C8}0���l�P��߽����	��r��I4�PL�Up�#d�c%W�9��o=x��Q��H���.�A�|�ҏ��7�;�9Z�Nٓ>$���;�$��i���*�s�
F�0/�St�I��xJ�P��T.�Դ��UR�tǃQ�gv5�dC��	t=�k@|�V9D�_�=��Ǔ�w^��Ԑ�e`U.�!\<emCK)b���ם-@�ɐ�C@�1�b4}�^g1�R��g��,�h���9�Rov����9��7��[�ϕ�S�D��ѓ�@3EM�	1��=];���qp�Y�ej?�to��ZƂ�,s���{��^�}��
���-q�{�Uo��}�'&��qG�v��U�Q�OY�xȻ�ʱ�p�����	�J\u�w��n�r,|��z����Ь�a�D/�|��	!5[�\YS6�`���gZ��63�������A����7�_Ϧ9;�]��&��ѷˊqv�U5�xg���6���l�A��3EzH��Y�,Yr�^���Y���d���c�ۡ����E�v(���E�7f�nM����7����ϻS/R�_�od���N<�(�����D�}S�0t�4���)	��uz�S�.�D������	��u3�'/�W�FJbv��8Δ���w�����cZ���-����D)��7���������������Ώ��&\- ��e��,�F&ڿ���3�9�m-d6,q?5�#x+���Ƶ?�3������H�K����5�4�/�9������7������"��'��절�^�zt�/�����[� � �G���L�y�e^����/����S�Raoja�g��>��Rl	�l	��Y����;M��\J���߂��ǽy8���6�y��i_��wMV��r�������1���t�Jn�xF*#�oO�A�q%c�Z'q+"'�֖]4�Δ�"n�o��sdny���(*}Ө��oF!z���g��E�F1o�o�MT�V�=�wg"��zM<"�,�&�RX�*$�3�����W�Ċ6|g�R��8�<�'��=��ۧflȕŎI��Izև���1_8�ؽ/��M~�����	�+2�r�5M1�,�{�U���/�W|n�:(�>C>�8��q��dJ`�O�^L[Ĭ����&HB�6�E�=`~��\鷊�2�k�-e����Tyf�
&ibyh��g�_��b�9��(q$]|���cgչ�9�줿Y�Ϫl����; �����bd8�2�6Ta�@�+)��>��H
Ξ."	���9.��+#J��\ŷRq�&�M�O�����.�G������R��Yq���V��n���݀�p������r�P�_7f^��5
N�z|\��/?ue-^ݼ�s�o����x�n���/����a�p4�+����Nۓ֜�S\S}�#���^KП4T�^���F0�~s�ۓ�)�j���O휭�VeK�.�[oH���|�0=*J�v�*��ԟ������O�{�!�X0�ܽ�	��r�;3�nZ���8�xq�:]�w5n�wonav�\w2���y.���?)�����:Sp#�[��Gs���&�9{l��t���f(VB�wM7"�Hϕ�F�Bb��;�f���ҤB`���9���f.QWZ2���N�4������]-4��ڧ�Y#EfxsD�S�;G:��F�����*�7����i�����=����֦>8��/�bI����v�<��_m����M�$y|D�?�~�g��w�w��!"mAN�8�@bAS�I���[��%�^r�x�lR��\_�?����Y�YK%|���{g��?��Q��J�����ݵ�]���(6f�mR�5l�lyhak+Ö l��~s��LW?N�n�4&����g�t�_�``���9��3���j]v��!8�M22�{�)�+DS���t���G9R�[� }�s�����������f�L�J��_��I�;�~��Ip�7!\wbu�yx�yع��"ƒ���q�נs�f������)�ܳ�9��ǝF����[(70�5S����-��ډ��i
�V��ۅ��>����}�J'��iO?JF��<���Tk~���`���o-�!45����uHm�B���9����ߞVO��%�Î�p��2��ڪ�
<9,Ǣ��L��^'��Mg���&W-�e�`���ht�6.}��"�'3��	ȵ�����ۈ�nCJ�1֔��9ڕ.�ѥ��Vzo`D� ��	h~��W���?�֐�W����)ɹ0�>I/��:��4@�T�U�{�[R�ٮ�Bi�������V·cb2�/��]`��Z�s��~���'1����=J.�Y��W�����/;H$��GDU�> �TS�e��|�Ge�5,b�����~}�_j�\d(Ů�ږ�1�[שj�9��vh<�G��p��{���i:�w�W�M5ώ�K�%��݃�o�n�E���[�����|�U_��C?���l�׈�A����^��"[7!!7Ds��"����ɢo��^ͧ��)S�fX�nM���-���A ��V�3�����n/��v� 1giE��.���v�d0�.oz��_��+��.O8���m�`I��u=$��uu�]���]]�EcN�ې�1�&9��gn={W����#QH=UҼqK��#����,�틽c��t�*mO����U<u�+|}ͪ+ͻ����u��-ɣ��Q�����3K����x�u���k�Ǐآǿ�}�Ju���v6ؕ�zH�8���JU�9O؄�H�Yfxu��;�QW�Ԃ���@��v��[U3P@��V�o��p{;A�������]3�����o�H��Rr�-�%+��:i*��|��}����֗!���ud2��-��$��)cq�3(Ѷ��Y�>q�~N�<$�
X�̿������h���yl�N9��P<$��]A�ݟ�nhl�n����b�'oѴ���� �>8sNO 8�[no	�bq�*����8(⥷���կ��N����u��bLٚ���Zo����q�z.�Pp�ϋ6wi����F;�O�+��#邷{=8���5��a_�v���r����!�����hXx�E�J��jZ׀B��L矊K0���<��y�~�=�������M0Yq� 2�m>�	�*�]��o��3�	t0O_�����E���9'?��*Nכ�;F����ط���J���y�i㯔�R�����ʪ���l��� v��a�q�&P���Mo�Z&~�Z�{Z�CQ \em��X6~o.G��5�}�[�^a�c�ê����]��1�/����T�P4f�N�:P%U�sͰ�Qh<[*�����ѣy��\�6p~k<���M���;1����>����E��N����!�f���m�����)}Z~~��U�v!�*Z���UN�>@�����^e��̛K$+��(hi �ӣUoO���ݑ�>�B��9�Oq<."��v�C.�k�ouwo�{�I�������,{v���:3aDN����d'_�g$��1s|Ֆ��u�P5{���m���u����x!3�IK��v����S�jDU]��:�����X &VL�^2��
�;!ل�AX/OiA0�Q�y�!1�NsWãϠdO.�R����Ͽ��1��-,Di˅�Ө�pq�E�ut[�O�����ٺ��yw��ޙ�ߢP����r|/���~6h_��Fn��mhU����B{�8/S��xB�3n8���;=�Z���:z\l׏���'�do
�{����\�+p-iWM���2��b�;	���M���K����ӣ��qG���)����q%�v��d=Y�9�/W*d��
͘4�Q ����>.x����Vގf|Ѣ] ���-�*�c"�~��{`�K�+�X�kA:�#Ց�?���6�	���I#)^���#17�O,E�:��6;��T��:�lO����Z�'��Aٵ1QR��43��yۙ��ds�Lrc� �Ŏ��N��)� ��-Eo.O�~��+�v�R�b�@���>?��F��[Bh���_��$I�����#�b��o=i�A���jW��d�wX4h�լA{,7f��$���	�G-P�,���t�t����-X�R÷�b!.��n�&��\u%D J��<ȞJ���!Ѡ��͎yN��5�;}_~��r�t��m�7������(D,����3��b;���ů �;8v*>H�����-·jVVV�ȥ�4;IWW�Դ4���9��(.�k2w�?x�V\lG�eH0c�T�{4�H��V'b�3������7�S�@U54V��<~F�k0�!6��\� �(f��0)u��"D�buGUYo�0����������Q�zWx���~7E�%�U��p5�>^��fğ�qp�V�`Lںۣ�e�,R�������0�oU��$�DvE}�~� j�����i���zJT�6 ��D:a<�N_J�v���fд���A?'}�vsWk(}On�xD(����.��7�z���Y���ti�&�ި*"��vH�T�gW�Qiz�����]��_�,��YX�}y�YkEV޼#�%)�2��y�}����J�
�JR�C>53��y���pM�_����21wC$5[<��ٽ�ot��` C��J���̮P�샎Ѷ��a�k��4i���A$�sBP!S�ݘ��5Q�[3ࡹS(�e��[�[Q��C�j�;~'5�K�7g����a/���~��h5[q$Q%Mҏ>)Y�zI.�RèmL���G����i���5m��mX=�,]�Gj��j���e�H�~�;d�tE�!07d̄r)��f)x�R�JDt*$�z�r�BYr
��VW7���	O`��?��!����Y⎸I�o�|�[Y�nk���;��^R�;?�����g"\�QϮw}�>�[[[��3x*���jא�C3q%�	����eT�剃�A#jQ�C�C]��8�K�$���Ws�������/��;:s�HH�?*}Μ��L9Qb�|h�:;��L
|'p�sk3��Kp���Kuuu��#$�F?���uS#X�a�T�{EEE�l� =)U��q*R�c�a��Q8-�B��r{|8{Sݧ�SO.n��ͭ��tzu+sX`��A�|'�p(%jE��V�}�Vĝ����Q�b
;%�2��~�Uc&� ��Ht'M�M�n�Ô�Q|H,V`>�T�EIE[j��skicc�Yl��[�%4UR��,���w�/*��-~���h���pҬ尓�'ήP@��#���'�UJ��3�rce �]7��/R��紑
�������v%1��-T�$}��V�K���q~�H�+�B��4��͘��ULBh���%q�L&�g�a��h�y�7� �2my��=��3ܽ�m�|�޾	�[8忲P���}ˢ�³��rM�ùݬ����E��2�a�r�h4Bd���5fQP�Hs��]��Uc����eN[��,������[�~�8̼�j���מOS�h]S�ц�Mp�����,�+�x�͂$��ܒE��K>��c�z;H������!z=�-�2�V[ ����)���L�6O/���ȥ?�lT���Mx�1�D��H����a&��F����K\%�4��~�ڙ�N/<;����5���C��>��z����|�4ֶr`B[0s����PT�N�F"68�NqqNU	��uG:1������\�خ26�;X�m��w�]����9]�R��I���{h�q�r��J�_��|p}��љ��7�#���M�M��)0���y��p��@��:�_��5�<�+e����k��f�P���j�P�#x���[Wu�y��(噡?��qKq<�x�Q���JĞ^�A"_3�(Z�a1�����.���1)٬��*-���!X a`�u

��r֤�:�la�vpa��z]8^=�k�<�&�;W���*�o�^�Iok��`4nc���I�Y�Y��o�&`�;�]��<z��f���tٷ�5�E���!&����Y�W�%.��#5�B��z�Q6a7��j�?Gd���%��B1UI�J���j`g\�*����(�q��l�h�6VD4k�)]jﻩ�Yg�r?;�% �w[�Q���7�Wk��5��=�:�~%(��}�4 f��<S3� ��}�_Cn�y��hz��?�7*����R�~i�����dV�u�m-A�!�`)�Q�LЩ���q��>/@��{�?�G���˩����)��I�7�0"����X�ƙs�4��~}Y�	�!n�
+��^#�\���𓈃8������/�py|&Ԍ����=Bj0wi;���F-�� ۤ�VS9�5��亹������xrW'*�t�3��N%Z*C�@��r}{���������6G���/~�������	�]���f<�W�:���H>_Z�k�5Ke,�9\�!�+xil��"�����y�s�M_�PL�ޙ�L�چ�n+���i��$6�3#��k&�Rq�<���[IrqGl��a� �E�:0���i�K����G����B�Nw�:�c�t�5�����_ˍ]އ�˺��w"����am�471C��s-��6�ZC�䅯�7��% J���р|	������V���4Yb76:�<�S�P蜾Ò�cu�ID{�� ӯ<��t��Bɷ�����))��acc��wgM-xQb�(Q(�4�	�-�?�[Q)@�۹&��.9�������|jx��n�N������J�i� Į��-
���f\ V!]@uK��"�-����w�Tw�2�X�_���\�N/x�8���vSdK8W�?��@����>��?�ă:&O��vG�r���=/���X{�����ı��]{K�DRJG��N���������r�ƱZ#�����;7Fi���]��]Ԃ���A|���M={�}& �LY�I@d�GU�@���0��Ե=�`y�6H>1PzoW<sx�9��q	�s� v�˳E�}ew���.u�7/�Y�-fC������Y��Zm��LTp�����F;�0@� ,��Ģ���r��{
5�
��.�àp�Z�h��4��0�JsK���Omu\'���n�zb��ۺTIo��T��Y,�{0���ϴ��pHVie����aIxs��%.[���U�g�fh��y�)�����iV)��LȊ��CQ:"q�K�vk��}��!t/�+?���z���;��M�/Ƿ.��ƴlf�q���1!pG�rC��pp{}=���u�(�3�(a�W���)A����o�����(	Ra<��B����m��^���:諲H��QL"Z1"�zw����;��3���4�&�usR�צ��� �F��L���Q�0�>(���p\�Eu��ۗ'��ؐ���~36�cZ[JFQ/��}�5bL"����W<��9�M 0�;$�������3L?E!BM�n5,����=F�|��o�a}U��b�w�s��>�����E��]�	���
�L���C��d��������\R!���E�zgל��+���Cs'�y|�e8�����$>xwH�9�D��+�H&��*L_�y���7���E��z�O����1��c�#�ʀ���9>>�8]
-�q�%�-!�p�m�j�w:	�ʲ\��5�{?��J)�����Q����H)b�����VZ�b�5@��#�RW7~=߼.���PD��s��Skn���ۄ[����A��6}�*q*��B�%�åyl�i�hP�&<gR��3���O�[",<�u�L�r$P̆.6 �<�(S�b�'�8�D�7Jh�w4��N �D�؎R�;�����^�$�&�	�[��o��I�g
%D���	�>��Ap8��s����59)L������@�|�nw��ݓU�6��h��MW�Q+VRI@�5�3���!MG�Se���j����w���iP����7��N��}1~��YG���x[��p&�����[d��@���뗱�h�5�],�H��9_���a��WQ�3��۰�2YlW��/��a
>���I֧��ciѝ(��^���{I��T�d *�b�U�����$����}@����R�/�'��ĸ[��z�2�7�"g�L�G��q� �����y���ad�\9G����o��'6�qWVg��K��'�=����b���W��͇ �E[EE�5���6#l�>Ϡ��?q���߅Z@c,�쐆�e����ȅ�!GQ�����*��tf���{�7�@6��_Fn��ԝ���2�?3/L�]><#��~�6h�x{mk�ۑNϴ�Wu�����U����c�Q�2�J�,�]�v	t�� J'���W�����h��-��I�ܶ���;U��z)yֱ@j������P�O�+��K����,Mٛ��(���˓v5u���Z~��G����_b�DP#s/�"5��Eq`�9w�U�v��(Ӄ��Y�vcHZ�
n+�b��*�#Y������x�W�߱&��n?`!���Eu!�;6���\=Y�^7��f��𰾰q�QF?��ԑ�Uo7���D����ӘwE�>tl�{[�����f��{���7/�aFJ��H����r�Jo��GkUm��}>ŷ#�'T��=�C{nۋz�o�Sa�0���Ra����+���s7��ļnp��N�Ճ���)��@"�C�.F}'�5�[�W1��p)0ӆ'l�Fy��#�F�+�D�6��M��(���c��޾��{ή�@�j�y��&��L	�^p7*��5+i*��҈b(��gn��m�q�����)��Ή%���R��yq�& r,R�<.����c&���u ̓���Xڶ�G��� ;:&|m��]`9)~_��|��r,C� k�P7��9��dQ�S��M�Ҕm�TLݕ�#&�a����1����g�X�v�%�8��]L�rՓ.������!)�D�cq�h]�;���ų'LRL�:Y2}�Kb��T�,��^Sv�v���8S��,H�~>Q8B;o��j�1� k-
.���\l�53�D�4�⨂yo�|`8��h����k"tL=RNq<w�[0�~���|��ֈjy��p�j#$RU�Ȯ+*R�c!L&{��1�Otj0�:h�D����3��>pOJ����x�qL"L=F��̄��oP(�ֺ��U%���S�3�Χp3�FTwoɫ�z��˗�hRv������e��?����q���t��(����B�ej�A��o��T��+�M01Vp�RNSd����yR���c8�ࡾ��s����L=��<���{nvQ��PZDD�ka�<�A ���^ #V��g���P���Y�5��!�}��8�2,�5��ST#�!�4�d�"n�~j�
uO;A.�n�oe�>�������Л�`pm��@=���W@=S<x��FD�6ς���Lqov2����������&I*�ȵH�Jz��~�Ë�R6��m��)W*ь�\�g�?F��������%d�.�7���\آ�G͟L�u�	7�������n��:��|5*U�z��Ǔ��C���_�x�r���+#X�`]r8m���zS8����G�<!˔�����=Z�@}7�?�ʲ� (�3����W�ݑ���߅m�ХZ-k��ӈ1�����S��2�i��΍�M[<��d��V!~G���T�������`����wQ��w�
��BT44>���<�`������P�I�:�3jq���xϗvmS,}
�3�KL���Ug���o�N/0�8{�`����̵��q#�)E,���)�� dY#$b=�A]\�`��䜚Ph��e$Ы\|jj��2�C�W"ፖ3��}m���@"�j�Y�a�9�Ź�9�s`�wo���j��ٙ��D��r��ؤF�#ҏ>X�E �j*��wS�3d�.��;�UQ��fu�$��1 �r��Z��c�{�1�'!�kk[5����=�
�jG�J*�Q����^q|� �$�Y�>�j�s�Ṣ9 tl���঒���Y����0�۷�����P��I����_~��������Zy!�-��4�61�=�x�D͌M�NR��;
�%?бҏ{2$�#� )������Ӡ�31YUR�x9�{w�zf���U�8�s��$��@;���R�4�5rt���,���/h�
�3ݸ�z~ɚ�1��q}Z���ꡉ��;��������R!o ��(�Q�<�~�L�Xd��Xَ�'Ύ=qOƞ��T�m<9�̝��~E��Q]ǩ8��5�D�;0��=Q�Aʒȝ��	��}�3�MJ㨷�+2��}�l��iaWoѥpY�g������h`�j�y�НUU�v-U��v�����)	a��'BL(�:��7vK֞�BLr�;���g+7;��/�"kf�(/T�㩎;��=�}6=�(@I��
/0@K��f��s�mУ_PUCi�Ĭ�k3<aQ[nB�;E%��f����H�鮳���;s�������iq�"T�H��QR��ڣ�*�F��0䕲���w��E��ۀ�R��
�dt7֝�m�1��@>������T��֮�=x�ұ�.��o;H���N��d�X��.
��"�摁�2!�y�V�|@o��n
���q�g�6@���8}�!ڞrU#��+���~x����n�e\���37�7(* K��d��%d��Q;�W��7K������G�6�CÃ߽�ݮj����f�� �>���GΖU�pS���ig�2�^:�N��'��<˷�}��`�?S��gJ>d�
�a���-��6�����-�m�����3�z�O����rAi�������p��W����C�M�k&�=��h@N����/�+���;a,ӑƫ�v�Äb�W�[�OC�+����`t&�	�7��c����ݾ��S�}�d���������c���/C�?�D9�~�C��T�h¥�x�+�k�f�F�kvF�K�z��9 8����&)�`!�Y3�?|u)��r�uD���yyn-�o�`y@�2w��1B^����,�-uy�#[t�����X<�"˹E�SXX�Ҵ?1Љ�:qpYD�����\"�jo9>������2�����p�+T{��f��[A���J�����+c�R֖$�*�X�1�ڛJkM9	]��ޓ�߰�UWx1�k���d���.pj�6��g[�iH��>bWh(�;5
�i;l�s�{����v{��|�J(�� �����M�juՌ]�n ����]��8;�@}���~�T�H��
<Js>����-Q|b�����Β�t� I��'�]���c�|��b��={vjc�{B��ux9�e$�'Q�=Z���!�&��ݏ�L���7�G�r�_����"����M��Kxy{�>�Ô�~��A�U�8˙O��'))�D��#TA���C�iG����w0 � 1��&�_>f{zW�'m��n��3m���*�M�;<"djS���Ҧ3�,v�A�ا�8#���0Ë����a��پ3-����9Ay�/ہ� .8r  m'�����q�L<)
/��ݺ��T�Y�`Ns3u(!�$;��*5UR��ԌO%��<�b��������8��4I����I�s���`Kfk5���^��gx2g�TW��i�*��0�;u��;=����ƶ��x&TA���_����\ɹOMK���=_�uc�y�����	��Q䯴��;������S�E��5�����1h6:5�n��.��	J����.��+17�����5��\Fu������!�cg�p���--�]��2(}I�����,�ZI].}kƦ.�׉� $ùT�9h~^�5"P�U�ڝ#v��Ñ:�Ju0�� #�r�63<s���SD����^�̺zf�����5U���i�_�n���O���;:�o��.�S_��E�ETP>::�gF���(��ӜE㺪_���T�����jA�֟8�5B�Lf����i�T<кp;>k����[XY���Ĩ��� �sf�%�e�yMM���� ��l�G�����*k`ԲD��p���j��-�����>�36@pA��V�ٷ<�����}96[IځV*^de�~�a}t/<����gF�o�<Q�}�6��N���V��_ �bQ��4Y��V�
x�@�/lF39٤M����r� I��U0n�o�E	��'�țb�P�I���[NO�5�U�7�[���!-�]���5.e����*+���<)�ܹ�Vp6L��-W�`���ƻw��d�D�r\��31A�a��uo? աQ�g{~�\�uX����=��4CR�ݡ4J)�1tw�R�%� 5��t7HKw	C�t�Ϝ�OϹ^/����{�u�Ͻ�z�,��Ckm��v�Q���9Q6H��A' qTTk�/���~���J�v���e���	�(�m�؍�п� ���b�+Y@���Q�'�2������W�Bm�IC��1�E#O��քC��&F�H7�"�� Y��BO�q����V77T�ty���ǥu��2aTUU�:�ك]2T;��΋>���#��(OI��V��+�V�'W�B��Q�NA�%���b����577ӇD�wo8��ك����ww�s~�q9�6�z��J��9m�)�`����l}�!i	<瓻����~3�?־[���TU�!��?�q�hU6�K(��'qO��$��Y�8q��au(������+,��7��2~`5�.�^CpE¶���@m�7,������?繬�Fb��?O�Hlk�p�b�v��my�E|���i�&�B�[�Q�WD �~V�Y��B����v-&��Y�;;�dڀŃY��QF����D�> �ұ�G:����(���M�I��ޚ|��`
h�U�;~��,c�����A�.�Zv���@�7�$~�E�w�r�ޓMVl%L��s�L;��I3.YTk�?�y��X"�C�M�,|c?j#���:B��^�3`l����m�W����]%� ����%�^����/5�^t.5J�u<���Ѣ�5)��K������,$� `��W��m|1˳�/�{?�}K��jG���0��+��^��v5�������ĸ"FMJ �2a��XB�;��u�����h�Q���F����ׇt���	������py���!�gO:�ƸS䐀Z#`��4hne%����pׁ�Q�8=>������c�؃�)|&�c�[m����0÷��{Ҿ{��3�;�d�O��y7m�� �f�Ͱ0)D"��).��,�3����K����7m����#�?{��ka$*��ׯ�)G��W�����zOC���b�y���P�ܠ�ݣ��$�-9�Gw����Hg[iv���=���}x�?���.GJs{������GmmcFo|�#X����5ӈ�{c�%�ۥ�c�q�m�e�k�����s�̷�A�X�)�����,�;�y�㉦��be�Ȑ	��9L�_��"��)�����g��T1�Rat
	t,��( ~6��*��套�6l
��ॏ����'�N2��G��"���M��U�� {�nFl�n�|�ɕ5Z������ ����*��"��i9�������l��---�9ocU�9v�.�#��=Q��=�3B�.W��%p t
�L��;���0��I.߶���q��Z�>��s�E�����n@���Tbt$+0�$A���ó>g���d������ż�dއɩ)�Ƃ�j�������h%�@ �s��`<�i����/â��	���a<'dq�GE�ڰU��u��-18�q�̞��bs�ك�η-��>~�%9��J��@�x�<Y��PG[3ɽ/�f[lH~ȉ�|~�s�q�u�׼�@)�y|	P�֒Lk�Y��%�?���|HY5担Oy���ECٷv�P��A��#S��N��J��}4VCz��9>Z�/zI�����ZH�����=��2��9d�������	��[�G2quf=�%��I77^���W�R�]�'��~�)tݴb�B��e��O��'6���e�Қ�|���h�Viα'���Fa��[���E;�`�#-*j�����_��ɾ1|�,����C�*~~���i��<5n�f�v���bDT�Ć;����~��Ȱ�G������k�߭j���*��^�#y�B��9
\]�IR�U�!��G�-|��Qn<�*��N���t�ș�|ݺ6��E��G���M�eD�}��͞��g���4&�_�w�ߞ~j')�2,�N��3_(|�B�^PN��<��V�+.&>?�Mw��J�A}{eE���Ѱ����Y*�׮�����B	F��F�R���P����B^�W �_RXm��%--���o2wjh善P3�(�z�����lkx�ֆp}{jh����Y3{�܌��4E@r�G],���D��<��j�x�ݯ! �M�:e����m�
�$_(	�S^e(���D�	�_w���|��b��O���׆c֍Ώ+y�"��	�y��̴Iqs;�U��� T+���:C�0�5�w����IZY�x.�a���[Z�@*l(�e��q���C����T'l��fC�kb�t��:sX8�d�|'*�����{�T��=�s�d����aj0ޤ�$����RjANnng�����J�771
���n]����go������WO:H���h�	H�V�2X����I�)r��;������D��.��o�%�r�4|����_�<��4�Ɓ�;a��%\	T/�8�'~� ϙ�l�\�ʕ�
�$�Z=!Ս3��c~a�F����� �|d�j�Ը�>�S�d�M�x���
A���s����	����6�Rֳ�s�u]�~s��8���iY `*�-,ު���al^KS�4��E���Fs(m��E�"�Վ�85�K�B511��Q"�^�m?z���Ո�׬�8�;*��Ҁ��t��$Ё��hpE���#ӈ�I�FV	����5���1Qor�e��,2&��� 0i)�$�a�����X�b�s0���*_�-��B~� ���5�xE����d���P�����'�o.�V�kkk��iNl��\T��_��o��ag9H �I��ļ�ω)NMJ�,��Qm�����:������*w�|��&A���es0���%C!͓�<5 �8��5g���^����G�6P�e9����l8|�}g;����5��l;X���[�w�J�1G(	n8�+#�B��6�74��G�-�����%a���O�8rcV��4�o �$N�R����L뺎a֗�\�4�ʇ�f����{ ���^�L8�ԏջ?�U-�s��
8s�mJ}�f�p���Q"j�uK���j&5bR�ݓ�k��Kf{�\ ���$�䬍׶���Hç�X6E+Q�)Z񉴝` �������O�M��+5���n��B�|��+����{g��E����h�`�,"��h�\,����̔��;J3�b	�}q&�ġ�G�]�����
�ft�X�?�t� �QQU���yr~~^@lӵ��{+�,Iϳxm��Oj,j<=���L���ו���O��=ɜ����yw�\.��P2����y��bAM��^����h��� `��rbr�L4Y�U�jky��_]]�Z��@�ܴqqxd�j��e/%��ڝ�/'����Oє��|iޮ4��,�<�	����B"A
�:ۚMFٸ��O...@���*f�h���X��"�����֋���7+��g��|���,!!!��SY�$���0czz�����X�G�����?~%���\�Wk�WJ
�![�w��ή��D�X�\Ss��o�*�������h�w�r��j��Nl)K��N������4�� G����!�U3\�*k���L��\+,?S�#�K8�]E.�惾"(��X��u���t!����W|P�R���;�_���4�fVdށ��1�/x/M3ѲP���܂KG�y��@�u$�C^��G.)�C�6[�S &�n�nğD��@�*]���>�$�;N(������?$��=4��j��Fm:Ra���0����%�08�'̚6&q�䒶Y%������8w#�H-0���I̲J<��w�|��� ס�뗂���y]���R��?X�ht큹�|I�ጻ����v&���ٳw�[U�M��6:R�ݝӨM��uO�d%����B�c��π2~anii��NZ�b� {XM���ޛ�b��ֶ�	��럌|8�����o��u�Xw��p��:ی�\Sʡn�R�j��S��t+��iֵn3��F!�g.wW'�BL{�L�D�}?uh
.�1�*�2�`�(`�W}1O� ���I�V/�� �o}ը�`���"�݈�IV��1�9��V#��}ɍ��_�h�b�UTx�p�[���\@I[;ͭN��mG�xȻ���.��N����3C�����X���j�L�?܃=�gWѪ�]�&,6ULH�w~��j�|�#*��' ]M�43� ������������Oo�����޾��_�~N�	�U�[�6�[�1�$R���������w@-�)-�)U2M}C�;�J�ٓTW'�[���7��;���� �"����=��0	���
_h��V����a�ɣ��
�=�$��A�ŗ�K��x�)Kw�~$z��3`�kR,Ҩ ʰ~�X��w�c����zk���:s��m�noi��v�s�U�+��wx�Br����,P�~6g]��X	"��i+)y>��	9��:U�q���#����G!@��9��67g+{n���wL�+T�-~z�VE]=(�q�)ZF�j)����Ca�$�!����|T���oK����a�a�?�=���y|��l��\�7���WUU�6=d����xt
\�d{�Ё9	�$3�z}tj|l*��zq�����*5X��fbȝo����{�X��� ����kV������bH�gw� 0��m,|�����)3Ł�K7^��Ր��q�$���Q���l�Ȉ�B��7m_[[TKqqx�����vc���2 @��#C�Tl�uA�\�p�Q���yr��z �-k�7v����V��ϡ�r�K�E��Ώ5
=UUVFn1x�!��{�b�nH-MJ���
�"�ei�(�7�tI�n��Cˉ��&�#a#��`�)-����o�����Aț�z�F�:~~��_L�Y5Wz�������~� �Cև~�QK�M�9k����ѐ��3A} 7hk����F ����B�d2�,92���'j\���M)*��w��VԐ.w����
��.>o��>�R�#;]AG; }w��������B�R� ���a�F+�
�sr)��������v�e���:~�0�v��&������L��<ޑ$d�^��=�Gmvnɰ���{����qr�G��$�Y���[�;#�T`���Hs����x}wUO�t^��- M}ί}E�	Y���&`�IL��6�mlz�oC�Df�[(�`��'}i���	�ެR�-��`��z'�Y�d��O즻�uX�����c$���8�!�KS�\�*��s�x;VN�V�H'p��PSE�wux-RM�eY C�FKbBw�]�vj\�҂�r����J�m�a��Q�vc�w���L�יL��������r�J�f�00�):11������,ǸZ���9(�666�]��[�1�F�4Z<kv�����C���(���rп��c�2�2����5?�#·�-,�ʌ��d?�&��w���j�� L�F���,;��b4E��oe�|Q�6�Ѱ��Q+�:�jEw�cD�ְj�Ƹ��!�Z�)K>�Qr��v��$�"ɚ���H춋|�� �&**R�6���������ԔI����0gM8����k�Lk�Ј����M�{%�a5��� *�h9�D�=\�f��(���{����C>��tm���fj^�~W��T�3��vBQ��8P��D��V�]w����1|Ksr��
�s8FjW����<�$R�A��\
��������t_�Z�/�I��.X�b���gC�dc��Ș�\��;���4�%Xr�9��>C��&�*��Sԧ�M#w����S䐤�H; ���?�9Q��g_����c��"�@%'�젪�m0���J�������6�S��y_j_��$�6Ӯ`��q��_ԠW�m��?d>\�}w�����ccc���7�ϴ�2�k]!�~}��=1�A�vu^}H'ةtn��F�>�����Q�Nïɧ㤜N�!^;�Q���p��$`�]G�����\�����?�oE}�c_]�X��5��2�ΐ]����@]��������'�{�
{�F=�{��������,��*�qk5��o�ֶ� ��|15<B�6�z#���Ԃ�� ���~�ʋby{pp���s{����?���y�5��<F��'��R�b�[C�`���|MA7'y�j�	�3X�,��Ȉr��(@�8��E�o�[��)�FE���I�?#ߔÕ)|��G�"���
+����q@�x�62ly�z6�Em��]t����r��E(�e�9��:V@�z➳vC���4jKE�_)�!𢦦�u��B�6~{���RxW�OCgh֧O�����
휽�U7Jt	;����$tO��x�[�\>-)�&��Q�w� �^��@
?'���i^yï��G�{�/��ܨ��CR��>���Ғ�Z�>�	��n��'=�>��?"����_E-<^�jYs7�Mlk��YYG��
�Sƍ)�/��L��t�����{I��&�)�PQŢ�4�F��q�#��?��Hn/������'_���1���
�CE�4��!K׮��6`sg��J��`Sg���mJE�ۻ�!m�@��u�0Ax ɍ�]�3�)x�o�N�D��P��~6�c�-1&kA�@agZX׊��62���#�V�<a1	���u*@������'6�Y��/$�[����a�)�X��RĶ2P�NZ���/��`�;"����(g�����]�\�-��K��t��á_�6�=��[g?��&����%q��@ڽƎ31����/�	��4�z�.I���BXm+�Jr�Ǘ��ʴ��GPw=2�t&~�0b���_D|{E�؏�CG�����M3�uf��ࡣe*�f"�@E���ڹ'3���a���&��a��w��|���.���"�BlQҍU�d���2��|#�$�3{��0[���ەG��dfg��@՝M=r���}wն���N:���pTV]�b�L3���^04=!,��X�	�}���jȑ�O�[ޔ��H�"���4���"G���3��t���7z�L�����4vU&VG>%��~�j�e�%7j.��g�Bow.ߵЧ{�JΡ�V��S##�6���zF˝�0�K��>��,Ri\LP���}R��!��g[���I�+$��I�%߲�%���RSS�Q��T���2�����w���	]K�R���Ė-;�@w�~s{�55��L����PD���u��n�$�Q`��ի5��U�����2�-�"V�:F�z�?�K�D)�����@jT	^?�
�x�n໋�h��U�~��G�G
�&��H�Ũ�(���7��QC�6��N�yzz�7h����l���n7��sG���ϻ�U��z	�`R�x=`?Od�Y?��.3,����jS~a��s����P�kty艏�ws�	�{{�j�Џ������{� �F �\��Z���M%���6Bٷ�=^,�6a���]���dեst�����Z^^ޘ�^!y��b� J�����B )����Qc��܈wO��bm.�91d����w)�z����7������x�\�������� ?L�jY0�w�����3mX˳�l�q��]�f�A�6��Z-��O�D�w���^ZZ�~�s�U���j<�(r�hHp0ҏ?^�b6M�u����%z���m��"{�ɶ�Iǀ/�K�1���d�e�V>����_`�SP�FK.=�e��gt���^T��r'H�T���~�(�`T�u�X����3>0-�p 3�G�J���p*�s@*5ЋU~�7�<�"���z�δ�@�=a��{2B.L���("7�Ù$Z�mB�m�o/@H�t�:�P�������I�����.0��'Eyf�xL�;�r{���P^�1���1MZZ������,m�p�l�H|+Ǭ^X�4����~f�a�oab�ݧ�E<E�(yO^t��Ur��U�LQQq����y�� 
	''N�t>J�-m�CV���q�
��ko'"�(���ǫh1��9��O3�l��?>��������ե���r�n�JY�07��BvS��ϫV�f�=�f�G���6_�c����CE��'���]Q���"*�&v�ԑ��m��&*#,���}s?�l{�;��}`S��{cy�������-�p�2�e8��r�v&�Zt'B�7/��P���н��~����i�6���ic!j����0��If�0�����?w�ؘ�!g ��}���E��Z��0��t�s��*���F݄�	~V鋢�Ph��=��+��	z	0`���@�vڱW��I�A�<b=�kor��V�KX<�@:P�Z&X>�q�"7YN�&w�c{�hӊ*�W	��=���6��� ��0-+�������ᥥH�R�3|||U�(݅�K��Dw ���BeS�jY��d��e�t7o����2qd�@E�0�\9x����MŘ�tq�S���[�rĿ����Q -��f8��6x�;�N��w����St�<v�``l,Fy��њ�Y��C�5���%�3�R��K�=��D"�;CA�<.Z*OỲp���%��f��Sn՘�vlPH�?��h�B�II��k'Q���<�e�~6PJ;f���5�z��T�"�I]^^�~=�1��K~"a�j�=R �{��0:~��
��Ŗ2C�I�kݡx��< �?L�H�]{����;>#�����0�X.�����S��z�I�����G�e���׎�g�-E���*��	�5=��e�o!R�_�r$���s��[�Ş��	om��珁�9Jc���ll,Π��9>yt�FZ�/��-�T��e�|"5NY�i0 rPu
խN������G��Ps{T�֚�Nx�͏T�<`�k
zi�P8�X���ϯ_�� n���N1�a���>E�J���!>�~4`E͈��6�Q��H$�"`	�0J������b%��1b�����bޝ$-��=MM%�n"�0K����T7T"�[A�תּ�aJ�nmM�������G�~_l��Y��Řtꕌ��߼<~�$C_�l�m髛�=eX�u&՚�������`R���n�l_����������8붺�Q�S�_�ճ��H����(�{m�\:tfk��hat��2�Y-d�"A�p� ���i�Ã�6Y��9]����F����4���]�2��&�Xe�!��i��>��1̒�@�����;.[�i!�,��;&\��!���T�j}��U�����i��E�A+w��c�Z���3���+ v�B	���bV=g���O�T�2��7l�|�=�������SIhU��P��y_�a��������D��i�+�������-� ��}���m�5���`����o�^���B���i|��Kll�Q�a�'ǀ������g��L�e�>�&�E$0��E��2/)t�K�$�5"��!R�_��3{�i.B��f=V��:�؄ȱN��~�]~�������h�.�ܛ71��V�bƪW�:�������,k���˫J�s\U�ԭ��.�D�����n��j���e���YkZ �՜k��H?����@�R@��d��PB�hD3ّF��p���[.@������x8Հ�OX�j��	@�������nH��I��>bOJ-���V:�%n� XP�oK_w���vlp��l�gC7� �6b7OE���CbO9��㥥�U=�|ڟh9��`��浳�d4�;�������������{iK����V���u�2ݐ_�i��B�_M!�����B������'�\������Rpc��=!"���6s�oD;\HHHc++���;��f��A��f�������]j��B��*{�剱fm��
��:�����F]�T�\�N�2��w5/��Z���3�`�%R\�/�������c�4���)H{u�pq��qz ����h�N��J��k��Wn�[M��b�K;�jn���T��J/�ڈ�1F��C�,�U�_ȇpA��F��jV!���@!�k.ʐ��%0���8���F������Uȷ�+پ�G�iSa��㧞�N��L�$�12rt�}��)ɯrZ]�M9��^iԃ�|��+������~e9w��S �i�q�c����e[��i��Z���(p�WY�YW�!AL�<���:U31��q�:�U�˄%�{)L�R����|G���w�W�v�t���Դ�W��.�9�� �n�i9�<�va��m�@��M*���!�.�;�:�|�w|�'�]��)���%߮����C!�B��&�qe�O%�8Â�VTVV�b�X���^-z�����@H�{��������Y�r�<UUw����x���p�w��Djc�$Ys���Γы�%��ҷ�c\SWG�l�OE���t����`򎊑����(��~eՆ\�Ӄ����;E3nF䵙�����+I#� ����m�=�4]H���66��~�e�.n5�_ga����8���Ҿ�'H��AyF*�^T���:��a�߱!%
Wr�ԫ�i���p�KBnS()W�wsX�k�~���~Cj�r�1rF��~����x�X���t���y���P*���JC�8>NY��,H~�g������"*�c3�Y���m�4	99��f�[OA~L��KUIqq��Ѭ�j3��G/� �'��m�����ʷ�g�ڹ4=� }7�Lڬ�dz�:?��m%߷{�#����^��l,�h0�M��ޔ���Ȋ>�~h��Uۦ������<���}�X��t����X��V�nT/�_���9��.�r�W���ʬ�,��
6DQ��n�T`Q����Phӗѷq����G-���>fpm���2�		E(��*ז�DPf�*j�gR��Еt�$&!��|�rղ0�Y ���-::�����p�q���%$n~��K0o2��H�2����䤆��g����Q2q�cZ���}��՜8{2���qr��~�.�߿(76�ҋ>[�M�u�o�0g2��G~�7I���;�_K���{��ݨͭV�Q�n]'/����'����l�N<[���L":�ΩpC#�TF�7^�] c3�sn ly���"���u3�r�����25h!]�{��O��}0����w`�bc``Ԗϸ,9�}*.�5!,8��Ʀ��x���p� ~�`�1����]�<*�ް^=38�U�R��u�����#��nW`�.���W�c�#*�Xtw	�@q}��"�/�AQ-^D����8�O�0m�vba�ӶX��#/�������Oty��dΚ �Q@�p ��X�K�f|b��^TRз�6G)پ߲���h=�a'@�3��N4�3+���z�ќ5�#d�iݴq�.���#;��q�(L��G~� Z��M@��&W P��M�T9r��qɶ����)�;n��Xce^GZ�D�]^>��0�i�v~\�v6�S�aʆ�s���:�Ⱦ,�`��!Zr�m�6�	J��|@t�N.C~=Q��lG ��H�d��F'�ѥ]�*�Ƌ����� d��1��?<i�@��H�5��靲��ώz��Sm�E�F���/��}�G!Do�-�4J�L]��+v�f��-��(eqs����yf�{�B݅����^�s�,�,������w��b��Ə�������i�
%+�\A�+��!�{!D������h[�П�P������������̿�U�Ag���J�U���&���ņ�@|t�e{��0�������_�6����ƋOPKK�އ~�bO� �D������ަ�څ�V�yD6�"�[
,X�G�@����)�)����,��M��?ƬF�K�~�ս��X��RI�� ��������o�=��~�w��]|P����T}����3��sXx���k�~q�d[��0���I+�aם�x�B��ͷ�)`8�b�}�w$��է�q�7Pz�S�9��~����?5�dyq�As�Ʃ�4[I]"#A
�o�s�s��5Q-������2&�P"��`��u@=P��F�|��AR�
����,�98���MB�i���.��s_����T��u�u}|Z6��W�_e(@���.������]
{�G�4�Jʥ���D�`#5\�_��23ɵGg�E�F?by��xQ㾶�-8	~����/YROF3Մ�AՉ�@��5g���w�L3�N;��a���_bd�_+ǟWߗH����U��������0�`{�����ʅڛ3����Z]l?b�@��7���6Ϯ�Am.V-�����R&�{`rrx#G��V�� �O�(�\z����r����Q�˨���f���ko�����>�H͙�ku]]2�?9X�h���(m�4S_���OTU{\fta�q� 0R^���=�\'�B|{�Ntw�]�ϓfb�^ڹ��鶶�^���؟�np`U�F���%����nxy	�oWn\qɣ�U�N,8RУ����F��L�f��^�<�0�}����	�ɋ�w�_���
��ul9�&�z�S(�ĕ����Zӌ���ـ�����Ŀo�dL���5��y���qy	9�rXs!y���C��@�в�t�l����+:����wg���36���X	+2Ք��#����l�B����O�P��Q��<�,t$6�T�[:��-GJ����#*)ًZ���ҽ۹�;RfI�3֊�� @��>�����0>7?��g�O �NEhd��G�u�ᇡ�����d^"�H�ΰED?����z�����Gܛ\FhGc���V�!X������_�|���S
�8�,S����i�g��ƔA6N��q�#�׮֥,c1���3o�h<:�-u`08�K�{�
3{$}�i��@�kҊ���j��Fɮ��F�̌h%}}x[>`, ����[R$��B����ʆ�ƌ�+�X-����3��=ᄂ݁�*�7�v�"I]O���V$�c��Z� %��b\�3�-�f��`,ѻ�eV�'�*ܫ�T�
'�i)X�J�c�=��{�+È9�#����7�\�� �G�p���`�ղ�J�b�8�r�ڱ��[�
�H.�jn3�8�{�k�EL�	���Tm��!���`�l�{��th�0Wn)S��;rs�T��Ȇ��۬����|�,{{���v�ݙ�U[��P<�������,a5ʧ���������W�8���l˦ '�������R�ej0�j�m��h
�ך�o�ܿ�tOM,��\5編q�t)����e�
`ǊZ��s;V���_�[u����P���G
�xO1,\����V�?yR�}!��p�NRZ[K��Mv�*@�$MnϣK��53��֪]ݸWkj��e`	t�Y�h�蝭XIm����l\=����=�7SQ�rE�����IG�K:¼9���x(�V���B#�.ڴ�ԇWwI}��f��9K�����^�wO��JUh��y籮����Q7T��J�
���lTJY~+��\�<`T{(�QNbq�Yt�j��h&���7jZu;��k�`�we�����>rq;��ͽH*�j�?��s��
�����e�ֈ;E.󂻋����3 W��j�� l}����Fw4��5m��b,	�be�����x
���~��d�irA����X�L{�U�G/�$*���.�XQ�4�H���r�������I�k�tf��K�q���l�q�a�|�4T ���v�������ڈ��|�!�M����I�=�<��x�e#NI6�� ���H�Æ���|�vj���9 �  ���ݿ��t����\Cx粎�9�� ;-HB�.�@��
�F2qj>����vN��D�y�0��m���w����@`��Q�g:mRD������qs�����'�P	�
OŞ��Cr7W/�]b���Z��?���W�999�Z�>���򸺳'�c��{A+�0aw<k��FCccJq��u�U&�e<4���t^�(!XRT�����r����[�e.�w|JNof�V/o��[�΀���޼e�-k�z#���~Ն��((�*rG������K�Ɲ��֭�c���B�]�~.]B.��E�D �EF|�;�*x���aI�_�%8��z���C�����m�Y���,]L��P	Dx�w��P���JDl���ӗw�#tq2��+ӀL�a���MSv�]97��>^��M]���#�2�Omo���7��(ę�=��X�T���Pw_���;Lw��=|���� "�� \�ߜ�G�{p�:����e{wW�ʪ�ώ�`�zW��]��!�N�ZH���|>��T�͍7�B4J�v}�,TB��~q�#���Q|� ����V��AĐ5���_v~�|� �=�SD���F��[:;�j�F�^t�jT b�,Jtc�Ԋ!}Hy�`q��t)Mwo��#�588�y���y_�ZM�21��p.�s�&j��Y�M�[䕤�F���777U���'HU�_����z�qp�Ɍ�~�l����	&�@�xfK�;�F/�Y�]!`	��� ����Q	��Ӊ��Q�7i[� 
�|}so�V�DӵQ֪�EY�t�si���
�Ղ����e�
�PbbⱩ� x�3�IKK�l�;hA ���_p����ԫ3�٦n��Hw&�ή{M���kIa��|�۶)��8���s�A��\��噧����Q����Ij#��/.,I]�xtcKK��>=*�<Զ��-l��d䀱c��t
C»{���G:C:���q�/��K<�ۉA��H�saxW!���5-V8�ჟB������O�5�M������ ���D>Hi�� �g��iz��X��n���c�uZ[ʅ�k��ah��Q�P{5~5%n���b�~��[2R����K.��g]k�7u�J�(����� �ξ�?��y��vT[�������qfWXu����\�-z#���ԲQ5��fW��.��'��m�&⃫k�4e1&Dզ�b��ZZZLn��l��>���/�,�eժ6��+�ڐ�S�V=LxWϘ~Ƙ��;�=#w��"#�5�[��m���?EȠ�)���S�)�.�H��rqC�''5b*5��|z�>�T���~S��6o��3�\�6����6��3m�%j٪��k�r�#�B�X��V�����KJ�c``Da�e�?8/iil�&�����Ȱ�%������p�ߞ�g�_���ޚ���r��<Q�?�U�_��0��3��e���4�Ӗ.^��M2��}����'�X"W�e�kZm��:�ѿ"+��»��Tֹ���E�?��z�F2��lN�/��Cir\����T��������Q/�âj⯛�n��(������ye�oUƸ�;�[`>{���[�k٩�y*���gx3�5�oZ�_�ʠ��T�RfӇ�)4��_R�N�7�84�h�#�o��F�?��;���C�龎:8��k�����������ڊ��W��48�Ђ�At�.1`��� 1��>���7"n�JX�娺��K��鏣#{-���1Ԩ�CSOWZ�Z������'�v�.�[�>z�mrU�׺�\��_�4µ�>��y�(Y?�>�;�8���i�1X<Ё���U���:C!� �p�$<��#��9[y�AGɛ$A��߁�jB:�<^WWW�S��\�������� ���r��-v�k�;I��������\@�t,o��2��`��W�<��ʼ=u��/�o�}�1��Y�pBq�5���w��*_�M���VOܭ��J��������S��ª>������l��Ve��1��ņ�F���o
k5=�i���Bp[C)�J���#�\\�M���]i,:_TK�H�@/��~� �K^����
�]ljv�e]���k�ۃ��Mo��>�m��ll�UT�S�l���M�D�D�u��͋~[ޅO�Kfb}nl� ��z��^�JXg��]��V�G��e����?^~�|���5��4�j|�j�A��	D���&���K~�
xgF��F�_�><<���*,���^_jy��Ͷ~�yr܅��G�r���E��E�����È��"�n��2܄"�:/8��ƫ�t����I@@�׶�"Y�$�{[�j���j�^����W�ԭ��>NN�{�^`���o�V��H6+��g��4�рC`X���&����Bg�V�k�lݔ�	FO�~�M��0]?�qQ#kke���=hC���Q�v�kv?�C7X��\��Aw�P��d���GV�B� H4�o��z.O7ȁ���7�Z�ߘ���C�m"� ["o�� 8��I��i��|��fLr6�H�{����,?�lK++���
ڍ�P�|+Y{0�L�G���ct{qP;��yh�c����ٝ�f�
��{iVcʰ)�߃7�^��iM����S���sOXM���5��&&&Va.~����٨��)N鴈�E��E�������'|Y,]�oПt�?���c��eYP=ܼP��F}���S7��+���w�Ga�8s�_�e��w�D�q��n��(�V�V��)����f�Eٻ �'n+>u.��!x�eE����q>��/�kH�S�3^߶{|2HiimS�lܦ��V0�d+��� *���H?��H�΢}�fk��$�+t>�����X��)d_8wc�����VF)�0���O5�=ϲ����	nZY�A��Dfqy���Z�{�\(�Le��ѓ�/�d*OW���;|.����_ws�Ƀ���[��TU��xwD� �f��B]c$�
]w�0��l/<�p��>	
-*)��9Ul�_��׀��;�}I��|Qu�K?�)�9������������/�E�vZo(ӠF����C؀U��OU�/6�M�?��$����������:���~�ftReB��?�{�wQY%�?]�ow;����`�_0-�f(!�޳Y����i��]62iH=\o]��F���-�'����MԲfrU-۽$vL{�����k�­P/�f�o��-:��U��=��NXҢM��'��V`T�~r�)C�q@��cU
D���G��t�+�>������W����c�������� ��=�W�����l��pc6y������3������n���~.y�[7��Y��?�ޏOM�*|a�<���͊��8.�̠����$m?}P}`��yu�����U�5�~o�iA��)�F鮑�D	��)a���RJD5F�0�$ƀ1�'����\/^�\��<�9���$8�/H���{���sCC�0�rd�>U��,O�f�Sh��/��
E�[�\-嘻Ǔ�����7�I�;�w�b{���	��ߚ�va6�� 氣���t ��g���HLۤsGFEE,�x�;C
��Ox:�ض���U��l�n�L��m�A��󑶗����
���m�l�?�(�|��V���c�'�3�&nU����&�G��e��T��3�$�1e�k�,�un�`�����fx��H�'�-�5ж�m�*�ҎR�7T� :�B�}�$>g��Y�6U�UHlN�S7���O��<�Ql�o�@ŋ����F牊G��S��͜mesӼ�߶�
��-�8*��}������]>#�u�Y?qk��c$p���X�"&���p#�6��X�<��9�b=��O�/$3������ܳ2Y\�$[����:����6�a�i�x4o\z���'jǶ����P(�i�N�uq���=_�H�߷���qj�5EV� �#^�|��T�;�P3�x��9�6oM�x�A�H���A�[�KL��E��[@ڦ�w�7*F�����u��S�Uu��t�)��O�=�(��F4s��/V����SKT�F����Q��‬����.m���̓\m���oz/���* R���J~k�TRW��
"@N��^B(�d%X:�Pk�fz�\�y�9��p��\���o/��P��Gdj/{� ����	 �x}�=�e�a�׷a����B

t?��"���O=��s.����\x<���f����$�:I��ٛ@�$D����٨��{�Aqǋ
��޻F~Dx=n�4K����(_���[��asN�^��QM���|.����7�3
�u��y������BG�ϟO'�۟����ƙ�4㪊qJ���o!��*k���ɓ�����9�!��X�R��G�7�w�Xf	=��J�l0��9���w�k�}��MLh����8���v���
\�o��?4��c>�(T�{�2�%�r�\�C �[��Z���ɿ�{������e��J���cz�{M6�_�/qo?�T�� ���M�Z��'O�C^��0,�^�m�m#J����b�2���P�a�srr��.~�y�Ͷ.UF�;�dFV�}�[o�����r4����1
� �_fq���8T��o�~�ܒq�F�~C�_��f�b*��:>��=��{LϦ	t��%g�a�Փ���)���U̑χ~�Y�к\7xM���W�J�^N�.�[��W��<�/''��JJ��/7Ӳ�ˡ�kXl6��r�}2��4U�����gx��Vɛ#�z��8�G=���9�U�2�,V� �3�2�|,�6;���ދKO�o�̑���)�ѓ������#�Fr��1�y�Rl�����R�Csτ%)��rҺ+���E�dU����{N�������f����A�����'��ty5L�f��:&�o6껊�	Y��{�n��D���w�D8 g�"�<z���VG�6��mp-kd��llB��|���L'�<T�]I�g�e�h�M�WóL�%�8���/G�d4+�@���!�H:��[f�����'+��M{��'�)�j_2��(�yr|���:����>�E����
91"�o]~u��&�[������yK�k筢��[�oSR�B�����r���p�����)U��>�2���
��^B�k��=�|y#Y�f����\�J����(�/p�2�g;����܋��*��z#n��MɈyX|�r#3l�Ѕ�J��Ǝo�x������F-�%�2����?b����'��M'i��tD��5�{&�Ο)Rd1�����I�R�	,�V��y�Mo�s�"����Zz���]&S���r.KD���>�?��|�,��cc�M��Ql&/�
+t��y)4��K ɟ	������G�zm�+���^2EZ;_���sn ��2\I���6LI��;���B��zv��rP}

���a<��ҵ��!ڈ���Cn����<~�N"�ئ��8-�e�Ը�;9��o�/�Ge�΁Y�����X�>@Ќ�
���n ��ɡЅ>#��$O����#@a����<7;]$/�[�����1�l�w5�k�������9��̔�ͽ	0������cJ h�88�}!g��	�g�$U�nei�NCB�A��|��iw�2�^�dm�	S��ݡ�Ot��2�E�\\w�ɆO�b�~;��*G[����$ˠ>�6,�8����\��xr���y�^���+�4u���>y��ӵ����%/�G)���L�sS�1u�G�����O_U7SSw,T\㑳��������2�J
�)���F�s���>h=��89.��_k$����ǝ��/ڼ1���I�	P�Ƒn��7Q^�ۮ��?ϗ�ީr�L���{�<L�O���R��܅_9KmA�m�W�{x��K�"����c��R��o{5Xy��%�Ug}�
x��Y�בG��� ���D�V�A�������s^�����$RϦ�Xв��*�k����),�?B�С
k��ʀhY}Q&A�n�dD<_��i���L���Ǎ~��tJX_(t|R;�2|����~�ә�	���͒�t��d��=���^Y�K+���C�̤�Rj��
HS�^�؄*żG��eͮ�_]�Z�.4�,�< ���EN�D� �1"��h�߲z*F�C�G ��qP�b"׃�ר)�J�u��p��\����<�O�~�����L��;�j����'������+��m ������Ǖ뺈$����0y�c�!i><��s��AW�4������^��q���o�80�����g�e���T6طbS�Ge�w�e����6>mq�B����&nb��j�`(@��m��6�+O�[)��J�mpO�/t�/O�����d�4���K �'=��VZ�E�x���[�����@Ր?�H������yE>�'ۃFsE�����%�⏋�v��4��_���&����i��ePL�er�����s��r
8�"�� ��ӝkl(�3Ɖ��3LV%�}�t�~�:.JR١#o��Ey!�xC��iu �ee�����d��\@���,6y|�Uz�����h����� �
`���pm������WsCio�m���U��չw���\��+�^jŕ����~�]��'z�qM4-F�CÞ���2�"H�R2	�Lړ�f�����/;�����^l�0���`z�CY	�@%����}~���k�?�ݢ0�4������J��ֲV1p�>E3Dww��<���{S�+ڥ`�AП��e7ó��݊�:�k��K]����G���k$������{�7Ћ��^,�����������k&�_Ң��(�^�es_�5��{fy���wJ:�g�@�n�o ?�������D���up�R�c��:�Ӟ�D���}�8���Ğ�W/��Q�z�&⸧��;
n3wMNN>U��<3�T��D��p�3s�3Fdt���3����_�H��7кH�g���{ [��N��'W��H�{G���Ƅb�����Ţ~�=��10h�����)��:QP��9�-����
ݓ(�`5�4fB���Ѵ���AG����°�c�U�zڭ!��@q��ȃ���Z�c5/ݹ����l�{ ��e9�*��4��Y�uB��?�MPY��8S�� w����2F�����G(ߪ�~����0r�{n����I���i�zZK�C�M�*��~�*w�����Ш�=q�V29Xv�cP�|����?�<����iY�~/H1�>;�</ۏ��yG�Ѝ?��b&�ق�X([b!��i|������ou�	��x[����0*�'!\udUG���YmS���n�F�A�u(n-�
�sC��L\��*��Gk}͟��mIW!� �˓D"?��k���5��׼p��5�DPZ��G��j�Rb�f��T�8�@��0?ݹ�g���;�SK�m ��4O`2��K��!%�gc �|�oJ�
Z/jq�Q�F}���y����+]�VOk�F��>[�Cq���7x�2E��/ �Q����d
 C9�,j՟�z�_M�~	��4{�e1qp錖7�<�]W�<м�x?�J�p@��I��_����/��䛹%�����H����s�F��b�����x�2l�<��w����u*r`@S*E ��(��Z׳�ׅ Z7�WM��f��B�}�wX�1�|v�;ڿ��0hݚ1�Z��0i_z��|ݩ�(6B`�b�=�
��d��]�x[��iyWVS�>�"{ZU51\B v�A�����B>��˭\�闣������oi�i]��627?YU��w��~v�W��)O�1qp<W�s�t�S� �4�3�/�[��n�}i��ռ����s]x�E��$��c���I��E�X����e�B����n2�վ��U�(V�PURb�nOm��Ol��ybus3돈�g������J�CkC�ѳS\I��Ŭ0y����n\��偃.���Gp�ʪX�$izO*B��~_�+�\��f, �!k��kEyx�vt���qNʦ|)ƙ�@�AE# �ڈb�~/ሷwQ�-P�>5�:�G>�vG"�]�����[�y)�2���"de�E�e��Q���L��$����Jޫ(p�
���:�Fx�ڞ�<�B�����Q������>4\���������Q 5����j���ݫ�l���K�B�
����s�{*�z�*�����O��q�x)��[ϗ}xtψ�X&@���2�צ\X��_�Q�U��uUK�݋{o�˅Q<��ٕ���*{����g� �u�=�W�=9����v.`�,�P�����^`��q�¢��C�B���|cc�7����1�����+�*?��6�y� ���� J�ӏ�Y,~��8��2l;ԟ!l����U�q[լ�.B`����ǻw�1��cN�1u��n��/��$E�����=%�;����_c#�L�D��\�y*�>��������A+G+�Jw�2��=�%s�n?6&��&1/t0��|���wTY/|AL��@����5�|%�uhPf��oI�C��g�C����Lk]�9��7�R@1/��	=e������˘X���#�9`S��


�U�����w���PI;�D�gi���g�J5e9�z���5Ж�oG�x�3v�ŵWZf}\�^��/)DW~���䘻�J),�XQ���.lk����"��X�i�p�7����_��AB^���ƴ�B����j��:��x5<Ҥ�/_�������TN�퐯)o@e�W n��RT��?AB" �G
5�׊"�"s�m��L�!���ܘ�}���56�k ׳%0{�4��Ѝ]���B@5Lz����5֢����]A���t��l=��?k����?�q|��ut	O;#�4J�� ڼz���/N�Y��ブn�o��豍q}V4R~!�����iC"aL�M�9�y��{�l��2�H�'<QY~_**�\T���э&���]����q�m*f30 ^����Oύ��2����]
$�.���\����p�l�L5�̒4�t�6�RAo{��������C�P��q�7@YX�N�i���\�7��y��,�j��0��cZ5���vb_�~�I��嬐�J� �h��s��a�G��K	O�0}n=ױr���A��"Ҩq$���h!'�'ksM���i�H��`L�`�&��m_���n��jX[bv�4�������R�x��V��3�j�#����@��чJ��{ܴ�H`q�`z#اM�2��xiU�8����^F�ܳ[���J�����o�S�9�M��g����e��?� ������l�)��W�ʊв,,,�{��R���r'�c[	}w��z��E ��������FV�X�M��X�6���_X3���ap���l�c����c��@ʰ�l��_���ܵ|�S�zf��_��,R�732�L��՜�X����|���38%whf��#���3���a5��|��\J� Qf��0Q�̳������)�~�x{���u�����&7��碊�L#��l�b�L����}o<VA2������Yۣ�pV#s�������g�h�$~�w��y� ��l7����X_ش��ĸ^O�o��{M��/�X�'9<^��(�`[��!#	�1�#k��W�;��f-5�驣�g���ӌ��sӉ0�vd+ ��k]M��m ��C�1�&s�?��'F�=�۞Ɂ�e�z���z}�J���t�;�7	�*��q�N�얍�Z�n�ێ*�l~���6�)I��ڋ䥕ǇhO"�W[k�*��!��%X[�n�����0$P��p  ��1�E�͗7a~��!c��i(���r��6VF@ot	��p	}�9�t�����Y�f�������r��T���n�q4;?���^�DZ��+R����NOt�D>{~:h��|$�":aM��;������U+���Qj��~��oiIVuTAnek[��A0}צ�����+u�k�r��d�|�v7k�D�������_�^���
7�[�B��ַo��U�$�R���l<g��_JY϶3�����P@�<�Y����N��ֺ���L _"TyB� ��oy��&F:������ΓtGj���>�K([Ѵ�_x�)��5d �����K�_�s��t�e2�lE[Q�6!��_�T��u��m�830����e7�&ϦA�Hh��k�?�7�P��{�Jz���~�����w��F�W�Wk⑇s��F_�J���ݼ��}ZA�o���<�XlO�>�c��;�&�j~\� ���(�ɐ
2�%%%��G[�o����^���A"�o�����X_��P�-����:+�5���{\����*��LxR�N�E�!����L�z��lU�n3���MU�U�Ji?��fߓ���R�q��!?��v�Ӽ����H\�Q��D��T���%/���G�kZ��ɇ�O���P~n׵��|(,�kP'uA��=_���ٚ�;�[=����B�p�Z���x�_uvr���>�;�8f�RO�ۜ�#���sE)����;�����<��=���Z���܄d�p��/�R�����.�v����5�������)驌n��s��#�0zC���8ڇZ��ܝuJJ~	Tt�Rf�k���3�R�Aj�QP����7�Κ��W���0�O�v�w�����%��3�oqPh%\SM�ug�����^̚��u�M�[K�{f`|�����vs��b�;c�z����k�،9�ը���y.��J�;%��/C҄�*Q$����c�<�j~�꒶���忂r0%�q��I0Z

p�6�QX>i�������\�.�N6j�G��]�vr���N�3���
|�4���{�C*��|�I�:`���o�n���͙&ö��<�yZ~�h���{%Hg�&��{�U�����0t��i���f1OB�B'��~���6�CM-I�		��~2o�����枪�4�a:�Xo����G�QQ>�?�_(ޯ��y��\e|�`�@�ؤ�Dz��C���*����Wk�Nuf�VV�O�X880�U�p��ZkKbIȟ7�?}���ҋ w|$:���#�e��Խ�]�ݸR�޸0\6��F�	�/��*~������^N&4t�܎�%B�!��k�
`ޢ`��Z7��hj���a�Q4M}� �m����)}�������n����ڢ���!K"�r-;�X�#�����Z�q��:�����B�SS�t�;��~���#�Rw��hET�M����@�.�)�1#�b�]ۨg��Wˈ�`w�]��X�&�~m@]��ygP����z����r������6���c��2r���5��$����*���z���cT�u��L(�X�������:�H�8(��إ��Q�^bk��\��j7��sR!]jw�r+r�ߛd#Te���;ys��מF)�`B�Ut�g�����6��?�t��Z/MP���������-K�'�Y�U) \$q���  �܎���'��z(ᵤ+��|�V���� B���y�Z���ќ��+v�7��0�89cYZ3� �gw��B*JO�-�`J$Z�<�� yIElll����4 ��˩���DV����d�8���1�w�1�7bi7��˔�A�H�p��bbb��>l�
MȖ��q�ԩ���y�zHv��D`0=ܴ���IX�bN�ӎ�'k]�'��Q>h�@Y��2��r
�4�4ꍀ�����W'+��$<.�̃��ј&l��9�d5W�d���Sd�����t�&�x��:w^Q6Xʹ�m7��l������P�	j�Napa�]�g��\u���'�m���\�g��"M��T�N���񫵦{�UG�pt�qE���.��mS*�/ ��u!��	X���G�<SG@�SPpY� ��Vk�b=~�w.��@����$6�� u��3v(uXO��U��/E"H+���:d\[��ȡ׾�WKܧD���Y����X�`#�|(�ɱIz�T[cyӛ��T �=�'�����t�]#K��D{��D�7ׇ��D����[��!5��;�13��W�Nkč���-ĺ�<t�n��t8��\������y��@؁��|�,
l�6��φȥ"��rQ
bE�Md�i+���[�!�����:���J������E���1�d�;�j���F�T�����;���muI���G�-�ݕJ+Bs�K��q�Aʖ�I�7P��88��3|k�b���cDBY���>�a�����#�5ݜC��T��YŃF�ֽ�B-N<n��N��hr(�-�����j��㏚d;��Z_vDz"|�i������u�w�!zr�cƍ�ݲ��Yn�D���[�q�S�du�S�; �3uL���@ٍ��	��U<n9�����4w�}��n� �X'L��ѫ@�~�ү��Nt��ɕ+��͵�DonL��v��Z4;�/�����)}�yh�>)ː
7��$�������\�{{�xp��{��;J$����D$��G���36�����%:,#����'� �z���b�i6��!�d�W? u�� ��cw����P��D���^�w��d�L�:���F=����n�E�bzhǣ%�L(�?C��=өl��s�{hbb��m�2��	wҁ;����O��N�G%>Ñ�1� �u�e�H:��"*:i)�:_3���Ȼ^���R;<��<�^KO󝙬�;}f�����c�M�C#6g�j���J��,���OV�ݖ�N[��X��{�*�1	&w-��2�mп��^l�o|��g� ��轿�%-��{o������O�͇+����1�2����R6��*�Z�kO�O����L��p��oyl�@������S�y-�����T>C�䟌'�~��I&����PM@����L���AHwBsV�l����o[Ml8��)3=�)�o�E�����[�9����&=C�@�f�Nn���P�� n���q�Ԡ)�����n�o�A����L݂0A�0-�����5:e9���qPF �ک�;+kJ����32F���ҽ��O��9�oZH�x\+x �����r���8��N�z���K�R]i�����]�l�K%��Iw���=m���͸�X �Zqe?�c������?���)���h݃f���_�����"%$�$��\������ ���eWu���C;���"�{,qR���~�E�E6Pyd����LP�2��R�RR��Nmu^hҰ�`dc����F7�>�$�֔�i��4�>J����Jg��9�%���e�yC�?~�^YY8롆�è��@|{�7�ns�<��<�=z�9f��@�U�SnLs��N�U��$�e�HK�����?�zJ���t�o�{���'�>��ܾ�������T=�<��Ã�"##X������O=�o��t�"Λ��cZ�3A K(�X�G@�歝��H��d���< F����9�wMT�/k>g�q�8�poN����q�,k��\MF4Vq:�&�MJ+^�8x3�`���%L� h�{�b a��=�d}�����$7��O�4<��zՌ餢]h�44�r�D�� 0�#@��������ȭ<�xN,^ԇ�qg�.��&�p��'�[\'��	�E�!�[,�'.��ZB��k�4�K�j�9�!}��T�u�p�[R]
�5�r��l�Z��%�b��CX��O��SF9�u$�w���)���)7ݪ|W����V;��"	��@���g�A�?!�j��C����|#J�J^�{(a������A��L#7}[�DZR��/�pE-���¸��$݊^�IX<�f��8&�ybAg�H8�"bjz{�S�M�gI�x���\v�����x�݃���N�3��ݍ���_�+���ۻV�����;BM�S���`��o��*4���k��ji��ȫ����P�P�`�!��� 
E�m ���+�[�f�TlA]9x��������l3���1dxe��9?c,�t�~��B��3֢H���s��]б������r�c�����sۿ"�A�2C�T�|�<U�`�u����e�c<i5��%�:88<m03ܓ1Z9&`�j�U��w��LDG�����9}C���x6�/Q�!F�]��QP�m��m�Yһ�=�8�����x"$���|p+O����1���[2v��e
����<K���������=��V�;�����P��� ����kba��6����y"|/e��!���[�O��dF�q�����U4�'��<��U����}Wf�@���xZ��������5�ͧ���l-�t��,����{|���F=�k�ws��W�ԧ2�{�ω���9�
(���>k􆹺�9KH�/>�NK��q��U��P��^<�0���30�e-fl7��S�y<��ٷ�'�K�U:S�N�O����~]U�3�8t�3Q~�*��Q�}�� K�S�6k�C� ������r�{U�@�<VI'���}�������e��?�@�_mmkE;�	^�����(7G��Z97D6��n7�n!*h����Le�,�%!�"�gCTq�V\8a8a��S�"�%v'x��Z7g�Wxb�[�⨵�ع)i��� E�H��@��m����ۍC�x�8�0�;[�̬��@�Y��aq+��N}{�tU�۹ڭ0,|��	�0�/ܜ�]�j��F������(r�tJ�Oh�j��'ӎ��	Lni�������y���@k�k-�<5�4Z��%ݧ@nWGu�|��<�n��&���� �C�KYƹd�fI'���>w���M��aG�}�|�g����v�]%������+�p�O�/Ҿ�Mr��-��"��abg��5���V�q���y��g�w��)�.�f)��1�8��<�My���Z[	6�3z�]�'�'�O�{?��h;��kh���$qËxd(y�P!g�v�ݎy<����-t��^�z$	��Bj�_�/N��>8��X�`D&��ŲW�O��P����e�E=k���;�秣"#�R�|+�8BDRډɈx�6n� ��ZA��Rp���������NSq蚝*<�T�v�����t�n,�(���u�7��~]rs<xFپ�J�����>f͸��os���v�T�.�9�k�^X�WܚL���Ua��b)�����m�skE�÷<_�ku�љ��
,�|�5�����ҸBMݵzVkY�?@���u>>Y�Ct_�g�x��B�)@�V�%C	�����{�DY�>��l#*K��O�����yb��P>
jP��6\|5J\�T(_�$� �wRͶ�Q���-١�$��N�}�A���=X����/t��"==.hsĞaw<������G`�Z{�<��Ǽ[��ǲ=������Vk�/�Dh��� f�'�qY��p�# �
D��-.�!�ke#h�+��o��keuķ|��c�s\�;v�47��>l}i�Y�g�<L��&I��&�����L
»s"�8��Z�qh(�bd|��/v��uL+��&L�n2��5��Q]'5O간�	�al�y��#��멮��໰��沶�)�M��T��3;Hd�6���d�/d�]1�-GZ��k��ȴ��&���-ƈ(y��˾��\�&�"����/�h���V�mj6{z����\�Уo�=Y͹J���,�������jX]�n���������-������&e����la؎�\�)"ܒ��J"b�<��C?���O]\{��	��8�`�-{�4�s��O���9�q�O�]m�>@��>�Ѓ�l��F��[�]��F�L�f�8��n�悖�m�g�;���͈�؞��	A�n4�]�r��y�(�����Ե�I�~�mS�I�#���9?�SIK�i���4ܛ�P)����y4��kn��ܐ&tI(���4a��mo��0O�0�-��!&�0a��R�^3\��S�m	��T�dghs.�ĳ����e8���$�q�d�0�������]�J�6�<�YXF��v7#��a��~�D�5��{S"�7m"�d�E�	�%7���Ra�L�f����"�7'��:��$�i���nI�[ުL�eNH5^� ��ăg��­Q���E�aq3�)i��4k��'3��b��!�]K)���n��@DÅmm?�՝����(��˽�7��Xu46�(�-�ܸ��\�ټ��0i����M#�nj�k�f$�3�Td��������1)�2Ky\dvȱ��;j"�'kf<��"��#����(޻j%ݴO�x�I��>�k�بt耟&��))�,:���X��!����f(����������`��#�����ik]8���H~�AjEEI��� ��<����p�,򮈤|�i��:w�0<ЏZ�.�tn��u���s�r������;�)[����Dm��y�]��_��lӊ����^������4�c�:#Z��[I�T(!�xV�m��t�m<L*ݞ�#Q��Y��4�9��0"&e9qW�%6�4vf�9�9�����|�n�]�W��w�{Kg���km�>j�wʣ���W�&� }F� {h��Hj�q����������7�]�8ǖS��e� ��j���;_Ԁ}��؏�U�܅E�pw:�$|	&����M��x�8�&^�@��D�������#0X09H+�9T&�u$�s�W:.�&~=`�<L� �iΊ�#o�a;JV�gL��6�?ۡ~�g�¡�F����o��q0RÐ7�?\����w寸�d��w��'Cj�˄㎸�N�����mX������� י���;����ǆ��A;���w���R�:�g���lLrv�8��X~���Ƴ���~|��])���كl������me:"r�_�|���ä���B�����C#��c��WQ�fH�^38�2+� P�>��@��-{~�C/2���VK�%�kd��7N���A� � �t^?�q�������h�[wl2����S�N�V���zgqC��w����Ә��e��x&����q�T�:��gϗ��1r��o�M����_��,�_T
o�0��a�F���ӛU^�/ �pg��w���bXN��mcg΄���
���k=��3n)��*��=���8��.W�3l��:�E;Sa� ��(����t�\S�zr`m�'?%lB�elQ{2P�w��4 ��x�W���bLȑ��E#��R�?��	������U�l����s�ePD��g7���
KψV>�C����!�0{�C#����g��>��I~��L�N8���&��ej�Z�"��v˜t�O��X�;phi����]��p�XYU�s�i�{���T�r
-���m!�#(������B�C�g*Nh̤q���[�x8�!_��n��]<sE�~Vs\=�nX��0��&�j�<�[�莇 �_G�9o^�f��+~�.��Ehe���#�D��Y�[�����?|�yQ8[���8��z Ϸ��5�c-:�i��W?�LoWHV�<�֠Ť���?��b��܉@�&d�n��B�_��]wa����J��llt�s�i�C
�{��<�t2�:�����ͭ��������Zwq��# ��o7��CL9AM���͹��2\�t��k��q�W��Ta��/�#^������VK�{��.�����L����|��D�s^1ՓWK����_�bA�'�9��z\5��KPЀ ��C"�� ��ag���M�t��-\*h���I��(���t�$��W �q��%�a-�.���v�5����s���||��`�Y�9?v������
�2�>������U�͙w_E�����Mr���ǻ���h�/�����GUF�[���cK�1�E�>�"aFذ�����e���&����f�c֚)\���c�Μ�Ⱦ����`N�~�<��0��>�42B�7��q\|*�z!_�=�{�35��T]�s�Je}����QV����,Ԣ�	F�BQBΈML8z�f_��3vx}�HI��qo3�g�B��gB^��x	��֌o_��~TE|S��,���$"��3�3�*9�O�_ۖǝ�N�Kj��P�x ���7GW*��"b/�;H��d��4�O5�/ �o�V��P�)����	zh=��1��zm�z�=R��kI�8T�C6��.fM3
��&3����5�ew�I�@��a�9�{]u�>VIX�1�[�Z5j̚7������K�����*���x���3���n�k�B!�m�h���!r���-!\�['�ĺGi�p)�#�kZ���Ne���8հ{��/��"?��5ѽ�6vFLg�Z�q,qQ��d���ĉi��p�9����]2���:ߴ���jLu)KB덱�^( ���������Ӌ��nՅj���G,�S�޲���u��?֞�߱���8��3���.%�`Ǹ^�x��M_������@���툋	����/[�IaO.���*���?�=�
�A�m�p .q�R��kn��0����1T-;��%j
��G:���}�+ܩB�
PR��'�8,�����T0P�ĺ���]<Qs�'{;NGԀz\�=�mK��T�[}�m���0��΁;޻�.���x.�4��Iu�ZC=#*��S]�ke���7ZJ��`�ڰj�!kc@�%�ظ<,���Kb�Q�@����O����l>e��0㭑�忩vϿ:�O��^#MFl:��Y���։�2GI�i����c�k7�� �vi+�jr��Z��}5�����ظ8�,�u;c�Kz�c�)A?�������J�����S��j�6�Y�%�2��Ta�5L������e�
�*a�0�9l���V���$�J9[�mN1�.��.�ê�����f|��&����g�m����߽�~p������7�O\ێC�[.L#?,�9���m�K������y�A%w����/a^P�X_��=����F7����<z�Hn2��>j�����x�q�mw�]}�X���v�������¥��D�o�l���T7\(?��B��W??�	խ�|ޔ� 2��|J߲Ԣ�?��)н��.f���d�^���'�V<�r{���[,�,�
̆\�YhK��k�+���G��Y§ ����(�^���V��>��\��lvu�B�#�M���-G�G�2�|���j"	�˘q��R|��6?	&�����D�s�{oK���_���㙬������oU���Q�ݠ�|�o��~�F����=E�fcǜ���C�/��2������p�������q�J7D!+��RS��F�1��l$F����Z�Ȉ�!J:���9�r⢴hw��y�2�<O��2r'���0�tE��C�M�왵jt=t��b�\u��
T�w5c���	�P)��^-���F"f�Y�����2^�{�3}��c`y2��.��x�G��Q���$n�г���H:�U�_�QeIԳ\;�xc*g~�lYf��kGjr���s�l>P6� x��n�cE��Tu��9a�署E�]�
�"`9�p�Hif�!ao�p&����(�W���{G^����[y/d�_>Ϣ��}�fV����Z+k���$n��WX���a��.`E�q* [�[=!���Q��ҎM1m8Av��jis��8�cL^���j0�T8#b�Uv�#ջJ����G]$�{�]ܠ&��)A�E�y�4R��2�y
M?c4�?��R�5պ.s�o��t35 m1;�W ��VUt� |`��^qq�|37\�����S�H7[�ؕ��C���<���F'q�	�$��u�-�R%���ͽY�S\߷�(Ǔ9�A��:�պ�`(�5��A2�����@M4�'M]� �b�ESu��B��J��4?��E!*�$E�*�z��o�^��WO�AM6V�<M��ZE#���Sc���y����<Q*V�3�T�1g&��z�a���H;)@NM}�Wo�2�ʯ��W�T�s����\�Z~:}����*�p���4�HZ�#y�@
""N'����港�W}�����?I�jR��p��������g�~1����0��J;S�s��_�U ���j�!�GG��ɿ�0����&w�h	�ar!���jk-�x�+rp	� #��wG��AF"���O���Wi������֨�p�u4@?-����������@G��cW
���'�Hm3����s'����' �-��0P�_C��qo��]���J�,�� p��P�4<�j��l#�@%c+�\0"`!h\w��12�or�bז�GcU�����ŵ�T1����L,!��w��F���ḁd�Tb^V9�t�:��'�!��j-h���s3O} ���7<�M&e%���uL)T�h䗍(3���kލ��3NP�
�rc�<,	*�M��%�i�jk+��{��/:�����9�W"�c����Q=(��(ê��M��I���i�rA+z��-�vnk<OU�4�b��L]TT��A�Ai�TiIi�F)�nX:�DJB:��Y���f��^JX��"��{�9r�03��'�^��N��?
�P�����7�K�S�'C���eri�]�����al3�����/�U���U�g��tB.7-5���ͪ�r�ۭC[��s3d�#^����{2�B�6�:�*������7L_���>JJJ����?�Kg�-��������q�!���w���]�p|'] C���"�����'�Õ�S�Xv`�@X�A9U�U�K=O��KIGX.�t_��Zoa��瀖 2�z꡻��:&�#}3s�#INc$�^%fj���>��ZVA_1j�@"���iW�ދʩ�1�1�T�����rY��iR�}q;�P �U���pQ�N����M�����\�ILLL �t��J �::���`�H�:�ۂ��I�ظ��Q�1kn��ICrb��f�A�����C�'q腠�O�e�Aӳ��\h��`�� �S�7`�� lC	Q�eJ�e#��R��4�s gE���S�\)��|�<��U���IK5@�|�<	%�j�I�}��������NV[z)+򫫫��>1P�ɉ��<�w��БͶ�r�Wq�-������5/���lq&QA�
�
��/@=<#"�l�}���Jcp<��Zj��-K�  ���@rǷ�
0�D���T�r}Wk�ܠ�ޠ����h�+��:�	�N}�Ev�	k��\�{;���  5���Pj��n!���u��p��b]�y Y@-ƿ|G���h��a�ii�s^p�f9�6��[A��Vɏ%�c��mdJ@�cύ���Òз"�X*���tƁ �IKȋM �d��P b���	$F5PF�]m>:6P��:��ݹ\�+G�k�G�H�L�����"+�ʔ� ���Q{ˤ%��ʒ9gc�HD��ݩ��1��#V�/u/TY/��\�Q�]�%4e���ÓoZM
~���D�%3s�|�+�ƨ�4�+�H�$���~��5��GN�����	dr��5��o;�~k�����!�Uj2ܧ:Z�f�����ǪL_Q��	�(@��SR��������SæEO�F~##��}*iY3�e��6�g�e7��Pn����(7o2�JM����/d3/gff��,�� �6'�h����F�s����Y��p܄=I)��{Y�x2f���[�l7��x_��vb?�K^���E�<
��v�kb���N����OM}�6L`"���۰2[	(�B��-�yL�`a�3?Q�Җ���y�Y-K���)� Р��$�g��J!5k�uR��~#0�S�Kp6�J���I���/�$)�#9X�����{��E��L ڥ�#cŸKO�����a�nZ jC��2���w���2T+U!�x��b0E��kY�P���Mw�J(��I �J�	�eŖ�s�~c@� ��Obb�}bwS��zj�x-/Ή�[A!�+����h�eW��R�݄T4��0oyAr���ؾU�0��г���2��1LiT
�M7A��c�k�y�/& � Z�����	�N�XK�6j9qO�s\B�3�Z>�
1-U+T5�Zc�S5e�����LnLOo/!���O�D�g��$8P���3�BpF4��b< ���X��@` �iLoz)�~(���ݨR��.0;�Df�3��0p��[<i9_�$�ߕ�W^�],��Vc�¢>�|w���.����a��uS@�[��"��>���\7ws�L�S�T���;��
��LՓ�����^��O%g�pI��}q�es�g�7mA�$ɩG�>
ޕA����.�_�.��Ѣ�~�o�r#a�ɹ������z��zo��C��e���7qb}e*�T�j?Z�9��=�=aT�L_~��m���ʦ���谀9��tX��Xj"܃4����\�3��V@��Z�fUVV��Ϗh<#�����R�i&�� D�J�/5݈f�����ޢ��N)���]I��c4a�E�ﺗ���*��<\��������n7�K�u��Ї��@����������������We6컍����[Yt&.��ճX����7o�l��-��J�PU&HT���0S�|J{hp�  ��>�e�4E�;+ H$L����Q%������;�˙���
D$o��^B������krm�sI/��ǋ�������I�WX
�^O�E�b?�"�_>�<
�� T��]W���?��]���!�="<<��U�>��z�����Co��~F�)�NNN	 3@�[;'>7�lp��X�����u��l�� ���}s�l�*qP� yD0 �(UX�MfZs����g\[��989���n'�C�u��VF#cEJ����E��-�
Y��F22255�e!���2�c��>h���n��������^(��9F�q)���0�B���|����;W��U��Z���e���̖�%6����em]�B~��b�?��, �Az���X�����HT)2O�$\Au��"w�[�-�5�v�7|iT}�@)X��t��P�a��E�'�|�JϜ7H����ry�[P��CX�sݴ%�l��o����q�M�q���vDမU�Rl��z�U ��8]�ڟ�$��duv�=Ӻ����� Q���� �|@�\@�X���b��{�<�zR��L��ŞC~���mkP�X���D��#$x�=.y���#�������Wk�ו�Ϸ"�u2n�E�hʚ�8`ص�� ?�32
d]}|(�b���vy#�<���ch\y��gbR��θ\t5J�_|���I"rk��c��� 0u��9�w����?�w w�6�^NN�9�j]������f��R|D����۶�H�vk+����Ԫm�����+��i��ښ������ml�ja�(��M��eΜ)C�`Q:�`��{��8wX��-|];f��ٝX��#���v�+H*���4oP®��2�dF�!��x/�45ץ]3�r߯����G���h/���ޝL���bx_k�N�#�7�)�S���ڴ˥���Ԛ[��4R[���m���hP�.(X<"�r0�ytXv�Ʋ�Qրv�F�rlH�	}�������"��1�/��4��VS��?��) @�U�^��W{��{�]l=�l��,!�<��˧�N������V�b�Y;I��R���$�/.���-�|������I
[--@�ϸ��Yp�}ߌ�<�?���qƸM�����" ���:��4C!�***��T�'����u���ձ��4VK@�����;	m[d�N�R@��L^)�<�w�C��N��I�L/������t������l�b7 �W�Jwۢy9��4���T� �ˏ))6�̉���,�����j��hv�2'JI1p)�&������	fc�7V�
^ې��{*a}����I�l)Ӳ����3a	Vf&f�V������߁�O��-����TĲml���Rin�IV��/ �S��@��KH�]�?r�ײt���K�kqߋ��ݣ�:���N�&��JL�n��o�8d�	A�V���jp�T���[m���V~A}���46ńT����� i=�/J'@Ʒ�k�5��k]"�W�XHI�VD}Ғ��'�e��啽Y��/����N�:���A:I�`�nmɺ��i��L���زŨ9'A��R���e�Q8h�p�D�JL�[F��'�d�a��u�D&t̎c!eȴ@g~5jd��/>S�n�F���w���U����<gǰ��#��r�WC=U
��fo7Z�.khI�|��-�g����~�7ݣ%}땐��*��V1R��ץUF�q�������ξ�c�A�^+Nu�Y�==��o^+��u�\RX�'�0\]|��"PeE�(�}WN�풑:]�8d���b��8R<mٳ�y�j��Qd�Sˊ�Q#m3�SZL�Q�������)�Y��yt
&-+ˍ:�[������SSs&��Hp6�<F�H�L�6a�����/��*��x!I�J̹�E����s<�h�sK�k�����������q�&�۾��m9G@���v�e֚��d�d\�|���7��~��:+�6��RSh�	�����Qn�@9W�6��"���|o�d��w���H�:�n9����H��2�̧+/��������Y�CSƘ�~�j/�T��" w�g��ΐI����6nğ�7ѿVx5z��M
v����g��k��>�hF�9��`PC��G���.�M9?|
~�gsB�T¯̃Z�X��~d��1s�W���E ��>��'��I٤��x���WO�>�>���� C#}�(�掅/��"TJ!��i����"����'7��5��ٿy��U~��%Kn�x��1�c�AnU: /���r+�A�^�ٶ�9{������l�L<>��V����0��=}��_�ސ���Eϭ�^9��3�a�Pa��.��T����5�A_��[N��6vv�S��q�����z�:"ҍ����Vc�V3�i!�E�8�{�*��Ga��&��6m��$ �G�� 1�`��ˁn+ip>��������d��oji"�]w�{{��`��M&�4��%p_D��Z�|v�2B	���̻�T@�۽ݱߕ��HU 4d��N�7�[�[7֞<�c�o��T	}��r~23B$(+��פϑ�w��^���u�e>V��o�h���X�خR�q�r"Hpz���w���C��Б�'�_�C��Ku����p��\:�7�e	��vHߪ��J���P`Ss�Aeh���>V6�U�(���>}[e_�=E%G��n��*`,�8����	��欃�8�Y^��/)׷�G�pgv���C/�o�+27z𶪢��'ډ�NH����t�7f�m�ߢ�����Sn_àW^��aK��A����2����=d�2U�_�:<�Z��'!�/K�C���5��g1G'Lu�njPz��s��8�³�U2�8`�Z�81�/���}����;���H��Qx^~>�yӓ��g#/b����ǔJ�w��mW���ݯ&n�+�C�D��9��h06��X�|�ˮz���qV,�m�ɰ��;����Q�O	&V[��Sg�R�P��:prp���[�kt�Z��q�9�T�h����(�_�����>�al�,*5�
�'(a<�89W굛�9���"�~��r��.��ҝ�(�1�����Q<4���G�H�Z����e%7�ѵU�)����)겵\%_����U]W�����Tduq-��@ ��K��NQ�N���8�u��Q�	i:���_ t'e��OV�G
�u��)\nF�c�9�ӑ{!��nA&�ƅre��U{��{�L鎞GSs���A���\�� �<�i����`.<b�������Eg��?,=�acv4���4��p��)���_Z����3�$=���k���R���itb��W���,I�M����r���i.������+��	9�yz�7,I��o�B<Ԋ �,���R$��hwN���|-��(s���V�����>��w��N�Y&�������} ~��ad�"���NX��^��I�]�S�Hrv�X�Jp�dA^�:��:�#pCw̟���K��+9 9{�֯������ˋ_��'��%����^��W�[U>� ����4A�+�=G�b���B"���4�G��u�5�	R��ф%�����4B�Z�/�<�U���I[4�{�6d����T��D�GDD0����9[�+Wφ�uu�|8$7"s�	�Rw�~��Jm\�H�7�?_s�E|d��yLh�ݭ�Ot�R¦�.O��Db����dXX�����WL��Ȩ�p�#J [;��b�ʒ$�R������Yk�S��Lg>ʢw� ����[�AH9i� �ݩ�����`4ЊH)����()'��瑨=�� ��R���m�@�u����J�<���W��S7��\U:+�v�Q�����t�����[��#ٚ���vbƢIˑN��/��h̷�Q�z��x��:h�Vsݶ��#�s;�Ҫ�- lV_�_�=L�x[�NWdl�>O���ޮN�rM���iU�ͳ��v$8~�57�NgL{)H,�Õ�m��f���ː
�B_�¦�����]μ�֙{2�6�g�<{��Hi{9������
�����ܔW[RMsB�FR<��[����O���������x8�	�3�̯��TV۪���u���%w�5]��B�;� ����&�;g�{Ӕ{��<�mC=��4[��w�Y]�����C�;K�Ó+E�8uV	��m������p���E̶�$F���/b�C�c� ǘ-�H��ٵN6F�T��� ��k��E��$�����2�}���[�޹2H��4��	�I�<�N��+^�x��]@��1up�[Dˉ���:@Wmõ�K���Z�8��
p�Yd1��ؓ��Ib.�]6�n�Q�ҩ�1]*�"D��	J6_��><��w��o6lmpS�B�����w�#w�{�������&V�I@D���( ~�FT�$`9_�F�W��=��u��ಞD�"� ��X��n�&�`϶��a��E�jMf�2��$٫��J��WeA��y��0�������5���ha,̻���D���~��,�c��§�U���r�wH%���{&J��_`ZZƽ�y�]�P5f��+���I���J��!2U����Q��ZO��N��*���Ѡ9'�[�Dvp9�<���؉�*�~�6�^��� ($�I�OL3T@��X��@\�_�E�'1�)�8$Tf��n>�"3�2��������p�uU�mmecջ�_�D.����أV�?)<?������ƭ�U��])aFr\�Ե��蔍�'�� J�1�(��r6���#����m
���z��5h�RF5�i%o�7�~]n$�?(���9-䨻ʮ�U��݅f��;G�aC@��2�� �i�
�g��$�M�G��`�v�$O�^_�h*<9ym���>d��
X�Xt�ag��߳������y���/+;ƙ5�g��$~%�p$������C�����$��i������]��C���ڃ��=�rB�3��W��$��h�E���t���2�y/�ᢦ9����=�>0��r�c[��slp��^�{�����	�����ry�xJDKKK�a�(��5�h��#�]���J�{�WN|uq�q���D�N�f������E�+���)K��[6�tO*�X�>*��N�|�5>��$0(��|b�;o�G�=i»�s�o�@�EE�	��Ɔ��ߦ����W>}�S��Ǎ��<XEg��ۏ#�,*q.�+"��+>���S�e�@6��9��/_nR'���d�9�'xl��#����x��͒h�4b�?~�ye=��ڮ�������S��,�X��!w�E����M��ȍ����a:ցS����1��ID!��
�?�l�r��`�s�8����SU&�L;r��翋��_3	���=u�ޑGK�P���I�T>��
�Ve��1���h�m����Se3�tH���9�}��[e�ʩ�	S>[LoUjq&�7�r���p��VN�����%��(��p����S��T����V�<s���f�I��~Z�ܿ�����lǖ��:���K㮒eIxq���f�kW���n�-���-�F2h^��1��'��_�ׯ�F�eO,�g;��hO����ړx�~��5Cӈo�{�������4�;���qfA�3���<:,=����/�>�o��K8F
�;F�7w���~>���C�k
�G_-�7���H�}Gx
�ؓ�T@1]o��9KחYc퐵�O���B4��5�Bo�+`C���/a��O5�������E��Ł�\���,��./Uٽ�� �219�?��2FpF6��@����#n8>�5�eB�b�&(��󫩝�g��	��:}��������m�4��	L{Թ?�������_�2����F���&y��"F�Y�!�6�#���c�l������t�����|��׶��ޯ2��Uz�����&��T���(��OSN..��Y�a��I��&ڻ���5��&�c���=��%&�8J���ZJ:�7O��À��V����r2�ݜB7f>�\>���X��������*]���)+�C���\�<O����K���xh��f���� �hB�䩉�e~!�#g��AX��AH�iT��4��F>� �N�i�w�ȵ��W�y��SB��Y�:�UՆ��tǍ�G7Oh���-OϽ��	��@��s���
KBYIO��r�3=�X����h&^L?����]F?iħ��瑺��;����ȅb�)��xQ�z@�~�@e*����_�'��s�s�b�R��{_$��u�#�e���'�T��0O3�t!����`,�6��s/w����&�v����Z%�s~jll�BMJ�r�;���C��n�������1KNN>6>n�=�A�	$533��=�)��;Y!|Q�{d���H����lrP��q������
����N�r���v�B�bߢW���,��9�C�����'�>?�oq���s#���*�y>#��\;�^=�"@�h�1�6xW�����Y:��8mu�l��Q��<i����耒�mMߞ1/���S��޲�	�5���)�-�+<@uD�j�� �kk+U�tWd�#�ϔ+��iY��5���7w�ńE�o@� M�L�!}~v�#ɑ〈�A(���u�0�3�57���qZB��,��6��y -H4��E�+��))�����p�<tt|��=/�V�K�.o!�%�����&L�;�]��|�D�uyuSU���0���y�ɨ�iN�h(m��h�	C��U����n<���.iȩ؟�4]>Ѓ>���:�!''';�5�wnC��FG�4�M=��ϥ3�j�������t��I��!t�kI.�7=@&�rÞWIU5n����gIq���!M_R0i�º�x3}ʧ1�@������u�;��`$�}�v��<��z�J�<77�6��p���V<>�K�c�E���9]��ٵ>�G�?��zfne��<�@"-����3>>�(y�3��O�͍��'wǨ�"%꧰0�N�[�M�'����1�Ѭ8�:6��6U��J��v�P�>d����"�("a�	�������4�ɦ`Ҽ� �%�IKi@ ȕ��^&�4Ĭ��k������| �%a�f�A�c�p�D�����
��c1�׏x׎x�߽C�����ɀc�/�m�h�7jj��'\���i��$������N�t�2"C��*y' �z:d�|�rv�]B%!!��r�������FVv�BB�A�|�{���#<�4���Mvübo�3|V�a�G1�.ν�e�Wc��EE�hS]'҇�)Z�垒���!:�;E:�tfb"N9~ӱ�k��!3B����ߣ���t�S� �U��<T�Z��lT��Ѕ/����-���O�}r"N�����	����#�У���I,v����)On�V���1M� ��)kh$(�ze���$�����bb>��&��:��`�(�o/!"b�MUb�4齓��ܩ�1��m�౉]لP��G���@L222<�����>��q(�  �̮&B�3���G0��>b^���,����fPN��������:���`�WJ��[v`�����y&nh �4_qi�tD�ɉC4�ECi�?��&/�,�����#f��
�[,�~�l��RH��Ф�hXz��r�`�|��D���D��ӕ��_�-(�T[[>-��4=9I�߸H�a%�B�CP�܀�.�Ʒ����ݝ�H�W�Н=��1����O�w�'�y� _@��;!g���&��i�y=_���7�ڳ�hyӂ.�����
y���zΒ������%��)��Ɨ��-���e!�����I���ۭ�.���hA�?iz�v��]�
���d۶����p���*y� �U��o
Y&��?������lӵi~��d�Wn���'�,����M1 t����)q��Fz�hP�V�:^�4��4�l�4��ߘrj�y�B�aM\jڵ�,qQY��4J���=K�9j/��$�����[8^B���TQt�O�"�t�%����r?z݇�rl�~�m�ef�u����}XT�\[�< ���#<�Cs��G044@�g�٘?�\49J�ӆ/��Ƿ�̆�G�%,��G�`�8��0���6���T� {@�Um4}��_G����4O��5���v�*(@��S̗�г��� �΂-����B��'6 �mll���4�Sc�����_�Pz��K=���"�9I#RF�4p?o.{�z�ú-��O���йj�g�/��P&�(���ik�Kr�C ��:�T�|zXGEm�Z�=&ߵ��Dd?����k�|��af.���+�噗I:,���%D��&A�F�J
� �/��S؃=�9��ݯ�"��h�]n��#"��4�%G��MZL���3t��mZ��d��ZMb$\���@��q�Ј���vϞW���'�'��j4Ί@X��AA���EE��� ��M�<p�<	�5����wl��ɶ���|�=��.  �T��Z
��@Ii��G[6��ˢ+X�2�ң���܃0T���b�'P�:��r�ȭ�J#r���`�+V�C|��MlS&�P�5��4'vr^��Y���g�Hu�F��00�a��E�"Yc�Sg�W
��p6��������{ʃ����o��ma�Oڬ�LE����Tjb�c������J�w�5+驫?�hB��N�X��=��٥ތ��ƛ�+iV�iW6h��kK��ޏ�s@KL�w�"�.-��ys�b�P�Ӌ�aqˀ��]�»��L�9�&�>T O �x�o��w퉘������$�A��Q�UY��n�$"�b�v�>��|�:�O�x�%�Q٦��	�`��7�t��;剦o+I����#iɍ���+@@'�@ &�J�:� �f=V@���k(��;��&�L��brw��ٹ��� б/B'�s#'Buv���@�x	���1�iX��-��	��-���.@( ����Jh�<���
�s������W������R�@J�)�ߚ�,\L�F�v��m�|s��,\���B�	�E�:\�E�����D�'m��t��y� �Y0pE���iů�zs�C���LP��M���Q�'<tb�����P�j�p]������8��� ������u�
XX���d�$�"Ω�>A(�2����uQ�@�ުA��w��"C�3�>�WVS���VS�g���C���V�	��ͼq���;�k���4G|\���Z㉆3א����ɉPGtF>���������C:����"E����?����UPo�����ZX����H}ʄJ�3,�����v�Q�>8 ��rj����ӵ�m�m�Ǟ��=U��܆y'�J����>�K-�C,�*�hB�w�F;P��ʓJގ�O�Ş������)�0�`�{���H�l�L2�bՒEs�ȷ��\�}P��3�m=M�:si��N��~��Q�!��i�df�um+<���߾ Q���)~��AYk3
�H�����aM��֧�k�����`�?���9(��"�e�ܽ��3>V����������Swb�ȡ�_I�d	�:b�e�9�ݕ�8�ѹ�#��mm��U5�(��CXQ��Ӫ%����;�@��g�t��
*����t�n����>���h�+ɞ!���u��j;�4Ⱦ�w�m�(���H�wV6�X���#QS;����i����>v)z��>�~�h&���!�����ķ��U�ƗZ��c\
3���7�2k����&P�ͣ�r��OI[����#<jWF�,aT�±�4!�o�dF��$��� :����#F4mi{K5)�bYN�u��?�d���EW����"����^nJ;.��ȤfQ��V��\�ňm���$'~�y�nZ�IH��o��I�Ԫ����B�\�)�}x����E���|^m2��ώF��/H?a0���N������I@A�f4�uu��/����)�z9˳,O� qMU��%��nCvQr�X�<�w�8����:�%�`� E+Jֹd��țc�-�OyX�]*�!��7nH�j��)v;����ާns{(�U��
-wo��Y����J��>��E���-��V�]�e�<Kw�2�g��B��݊����^:]��osj�k�M}0�'��Jov(H}����ӆ�'s?x3�|���q<�b���	�jF��b�X��%7w#0��e�������4���*oL��ߞ����+3�C�D}�ަ,��u$Ξ�n�q�>C��dٟ���j�Ĺ����n�/*��l��>��M������Į������H�!�o?qό�d����pv{Q�X�2� ��6E?������l>�	�hM��'�xD��M�1�"d�|(P����I�\L|*���-���>▉$@X����@�C��-;n��[�A�u"��B���#(�w�4�]T���X��P��ܻw�R�#�r�%в�E�"�g��!l +��^���	m��f�7��3�X��ֆu�>�A��%N�oxÚ�:W�b�G��1���Ԡ�1~�Y�Q��E&E�ƣ�{����r7F�	,ko �e�b49�b=#(�����N/�����������8'�=����˩|��uG&]���{���<4���o����9)��o�&����A2h�R#��( �	&Ǔk}�{��tit��=��,��@V���/Y�E�T�����%*�#���>��.�P��%�zM�J�?VV�l��C�q�}��9L����U��$��w��X��YDwa���/ϒ�?�r��z�����ͼ��jj�4{,I��ׅ��+�>����r�C�jM�h�Y��Y����S\W����e�hw���������b�?��	{To�S"�\o�:O��:�bZ���V��3K��v��k��4v`�a�P��/<���I�ߗ& s���߶�3;B�M�M�	�Wi�`�,��1 ��4���������ETby��z:��%�p^J���Q�vJ$HZ��~�nw�I�-��MF��Q�����@��Y&y����&D��DP������YN�e*���{P���2Y�f���W(�:���֍~}�&p�ـ=Sa�����Koahe��ݴ��N&��z�}�����{<�J[�y~����!�5d�L�s�u�"�7Ph:�,k�dt;D���E~��5���xZ�`��a��EP�X��ɧ0{�}��ھ���
���{�U�zAm�]�1ɕ��j_ �OTXr�A=&M�N0�+�q��<����߾���VP_e���k<���� @�G�jj.f�(�zoÒT���v��m�x|"�;rYӧ�gZ�^����3���U2�����Cs�(����5�Eے�2]^O
�T��=��@U����IU�r4�]��GQף�i��S|^;��-<�$�!���
�L����EEC�,�e-�((�[7C��m����!��_k@���nh�!��8��uN��;>�����8����!XV���=���3�e�?n�J̏	ł�P��"����q�f��W�^ǅ��F����P3 kȹ��$	�(_�p'�����@�����������⺋~<
��3��*&�1�Y�gv.�%���Ag��"<��x]�l�z)\�Q!A�{\W���Rf���@A3o��e<��� £���UX��]:@(#�1�l}Q8,��Y_��gv����-��:UgtQ�i��C��К}Q4�]�t�D����|����.���߭x����".�����e~���vgۄ�d���ߟ�zگ��1<[�}��H��Pݛ�+��^>�����ұ~�&N{�����ifއl�P�<��^I��Um��>˃��}(�e���#�B��[+��W��Lޢ"X_��}�"qQ���k��!Wr�	:U�|-�`MjI=:x��� .�`�\	�W�Ǭ��)ea7�c�����w�w��x�nbD=cj�x�[��p�v� ������
gy�w�M��-� %�Y�gzra��Y�%�^����)4v�W����z���c��AR�3Ou����/6�8{`q�q�a3]������|H�Y�Z1�>i��R��������FP|>󮶒\5[������X"
X��o�Ĝ�M�0�qeAzz��Kj��@zE� N�KQ_�%-N.["�'�}��{�o�����3��c�ˁ)AV��x����,^W���
�^����ΣR;�b�n��w�C)<���d��D�n������Ļ�q2n��XI���R�[�a/�?�����O����,I�_�'�|����|�9�ԣ��`١�c- �#��̶�~~������iH���4��ɖ)��E1����h�|��=^7(�c�sK���FK-~�i��?��_�]~��1�����7�J�@�/�F�Y��~�+�c�D��#�u���reJ	>m�m��8�.�=� �$W��E�a�@�}��Ȑ׾/swZkO\h'6�&�I ^�q;%[�"	?�^�,��[>:JXP��X����,erf�ē1jy��L��z\\��A���Nj����d�N�SS������آh�W/��a���'�:��?{����i:h�c��i=�ݰ۟���.?!�I�s���&�Cl�}�w�sv�<ן�'�
hΜ
B���U�d�B�Et;�y�H�S@��JvL��wZ��~���˧�)�Q�c���˯��J�ll3V�N^�WH⥘w�qB(�]�F�...�t��:p�:��w���tY�M���g*�S��]~��}T��(��&��������dH�i�+�~_���<x�V�?p�
��/G�q�g�%�s��c�j�94Q�h��yr�TP*�B�)��<	fH�9*�	WV��|���Qv���d�n�+�]���Qp��Q���+�l�%��1!+K������(dds��3T8!����Y����V�ަ.��o� Z�Am��2����\���ɋ����_Y(����d�o��yЊ��S���e@�K����ӗ"�����O[/c)x�W�.�5G%D�Oi�3$�9��_Q�g����-���cQ�|Djjj:��3U&aj�;�z�IĪ�����[]*�	��e���w�|�!�ޟ���%�l-Mu��̇����ӕ�i��3��d��T������z���Dp�e�����\���i�ڿ�����`�9{��l��;�''O{.��V����zyv�ʲ��|ppv�+�ps e��
=�c�g�Z+m�@���M��Yw�Au~�,ּ��o��dvu�f�|�a�kW�{�jxA�D*ls�1�������d���K���ZA:Aՠ��s+�������K���u�G�t=�^�I��G�J%�C�?}�Z��Z���*�P%��C�����!���Jji]v�G��d��>���"ܜ_v�92�0���ܬ�fG{=�Q�K��*>ه�J��i�C|����d5��}A�/>���ܐ큊��)?�څ�߆(�X#�&��T%K�+*��C�߰s[��/���c=�<#���Ň%OG{�����};ߦ�bA�b�Վ��SM[�l��A9�hWp�f��! 2O@�rF���=�������	%g��
�Y"�k����������+���ap�3����c��-���ڦ�0,J��o(�z9t+vvSz4�zo��w����TNǗ~�B�HR����m^�zނ-�gd�?���$�|ڷ�{~��*1�j������ _;��/zs�>y_��HA�?7y4�[�ys��f���`\�H;��w� d�,��w5�����oEqQiMM�,s���GC��dG�gna�fq,�bQЊB���o4���`��8�jj���G-޸����7{����\��#a� ����u����T��F���P$��3�����钻�hf�����WmI:�0��톙�)p�mR��ܮ��іc�, �n�����U�1������U���p�F]�ǲ�*}��`�s���{z$u<�sgZ<y ��^�N�ܞ%�f=�浊���{5�
U����l����YY��p��U�}�a�ҟ\���h��9��
��i;;ۿ�@	kU�Y�Wo�wO�.v�{R�U��NG�3��0�Q�=E_+�q�K�z��ȥ�1{�����,uj��j�y?NO���"�h��cD�tl��|߉�E��Zb��Clҍ9S�AU�G���� &�}^��:�u�9?9Z�<X=��ｂ/��ᅳ��fe=������v%�E�y7�h9���ձy@38!Q�~��׊$�_��=�rC�ӱכIg7���2��7��=̶;���h20�9��^�g3�x_^��= ��l�5&I��8�*�8�����7���k��2~��ŕ��Q���ݻw�~��z�<a�\[�9F�8[;���[c�GM�W8��������Ő���g�����=����Yj�wX?�s21f�;���cQL��ߚ�%�ыܙ#e�'����8+�0����g8�K��qV��j	C�W���A4���p�k������{IX�(-eb�@��VzF�`Q��%(f�w���<��c�͕xY;��׎'������-�0�H�9g�����*(�?�|h�����t��ᴂ��o7�3�1�Y� ���q�'	5�{���0�V�]��>7��r�/F?�;X:j^(��?������O�k�/���;���+j�U�zA!]��jI�����X(�vc�o��uo�袵O��k���A��~�ح͚et�0Ȯ�׀��
���~}�o��z��C"�������_(~bBM�����	k���F߻V��(��XuȚ���W"�'�r�`BFڦfd �#�qd�ƳS: ���JFn���>U�5��l�h�����w�5&������V��ɹ=P�o����zȷ`�s�O�� ��>')�$eݖ�O��m�������$��������0%>�����"1����J�T¨�=â�����[@Eu�߃(%ݍ 
�14�"J�tww7�����! � ]�t�#C�мw����o�k�r�Z�=���ݟ�9��ۓo�2��� �?�ZO��?)>yD��o{�
��|�������~v�?�	�uy�̥J��FbiiI-<���O�'�h� ��k�;��`��i�'�h�|A��w#�*
��;Ģ.�]�R�_��%�6����0��_y�Mm\��@���p��WQ(;xv�����*Q�IWh�v"�*�x�9�W��{˝��BJ��u��E��ߦ��n���uOch��T��T�'C/AcL%�	Ϯ�>%'��C�kv�������d��0S����]��P�p`�j��R'������͊�����vg^#�g?מ��3� �T�{V�N ,�#	Ru�"~%�8.����V%z��Z�	j���2d|�r���,����.�'uBp!=]�v{s�*dOt����Q͒��fC���F���J��mGKʬ-�߅y�l�7������e7�?���NWWׁ$�
�z<�G���m�-N9:�)Vׅg8w4/�<��_1%�s�h�Io��sin���ؠ|?/������8�RlY���L�6�px��z���R�^����	�?+�ъ��-n.��;!`d��Q����̭VA�.���C��y���:(��V �ݳ.��1�{W�J�����-�9b �%���V�!�|�MI�dAA��;�}�jjo����k������������:k�koc���	(�w�h�\��z
E)\`�,"Ȯ�b^�0�~Ҍ���F��}���<|"͗l(7��/��]CM�|^6��N��	�+���e��&����4��4�Ϯ�\���3N6S��ch��ҷ4O�N���"S��hz�	$�����0lnMSKA��)UB�HY��`���M55yy��?���pi����U��;�xKK+�oO���.-|y��ѕ<͇ʊ%Fw"4�}�@_�T�B��c��t��A:�oa�I!�	e��į߄�=6��7�]IO&��H����V�z8���F�RSC"��	ؾʺ;'"�d�@|<|�3��|�d�U>�^"�tb�P�yĄ�DV�v# �X�����
�묡�@ͪ��C������������˷o��F����O�4!C���O��E��mųZF�a�+�8Y�/dt� #��Q8;�]�W%����R�-b|�h*+����C��m��WU�\%}���h��|]�����ͧ[4�J=h���������Ӌb���#݊[�4s��gm��粲aBi��XCi]� ���J�̷O�3M[���}��6�I�������;!7^�N�Myh�D�mmq1�S�x���Ֆ(ʹ�_�$�;8���Si鼰:�̇o�֌	E���b5LF�������Fh^i%�8��{�P��كFս T��I��|7)�%�y;��ꧦ�tˆ�c3���y>�*�e�;�9���d���ӗ�&j�F	{ss�Z�>�� H]
��_{�m$��ݱ91嗉_�F�Ol��|=�k�}b�s�9g�Q�>��N��Q�-���쉍9�b�ƣ��>�7�T�1>N� ���%���ƺ/�%\��Z��6��wاO�����rDzj�)��w;���L���Κd�=Y⃨h$��=�����S�?�8�HxǄa�g�����dvk�Ẁ�{~((k�t��m�n�����=~�A�aT�%$��ѣG�L���w����n��)A���#Yq�k7�4���� �~���@��W�#�
�}��"�����_�s�c/��	FJDz�c���G�%�?ݺܩc`X>�` �70�3��h3b��]�S�ָ�M1����v���|}�x�z,��w�W>,�'ny9�J�J/]�?���<h�@'c��+v�̒<g�t<�����bg�敌p�W=�S�/6��ohO�h/_������+��~f��~�T��5�jia}	���IǶ_J��i�RK�B��.9�FZ1��g���i$��)�ĭ(��A�{+oT�(d��~��f�A�A�����_o���r �+��U��6��Å�W��ȍ���-N�N�]y=Px{��;k�a��Dy��m�ir�J����[��0�i���m���Y�D`�Vk��>J���Ś(R������Q�NF��r�RN�Ɏ��-&G��)��SC����DLk�p��w�a�������F���np�"ʽ��W�Vҙ-�Wc������W�F�D�]=��a��]��:�l��|�� R�q莄�v��q����M}cL�.c�5��K)~�W�i�B����ы�J}���L��	���H�؊Юɼ�q�M9ݻj�)�s[ZZ̓;h�J���U���J�mT��j2�$���8\�旚�/������FM�ů\{g�Ͽ`���@���?ԭL<T�"ǻ��bD��e�x-gM�G	���D���S]�}����]~�y�6יg� K�`
vj�|�{����B����R�����'�΋i�c70u��Nzl:U��^\9�L�h2�)ש�s{�tk:�.�dz=A���$su9PZ�~R� 81��U��y�I��@�o/x�`��p�8$�l�C<d�0�svO }��{�X��ֵ�!�&��	dl�39AR�Q�A�BW��y�~�
?�e[i�Q��H�I��I����r��U��}^�r��h��˩|���M������b�_�jj�Ƽ`qNox�7�Ys�(��:����֙\��Q��ԛ�(�ֹ?<l9/�ݽEu޼��n%܈�!T�=2t�-i�n�W���y�8u���̷�/�՛���Õ6�7e���h.&�Z1��J��t`���R�9�� }��u$l�b$]�~��f��	X�2H��&���woԔ���ӽLP"N�FA����/$��]Bz�$�M.�κ�A�I7#:��d����{ZB�0�1Q��k''.j��������a�?9�,g��^'����:����bZ��G.^����������ڄO'���B��q;��-�g��C�]Lqi� nk�^1&z}��T�J�Ơ13�a�����4T��ޞ�������y���LS�U�n��i`��6���+ŜSi��{�`�:�M(��F��e�۽��WtБV�OAb�58�ݑU�m�/�F 6�T�V#��c��ᦢ�N΁����ٓ������݃nw�$F=���)?Nu=WT1�����/����bE���쵣\n�Q� ��7mf(j$~V2��wKi����pj����D"����[�:����S�^We�>͚ #�R�0i��0Cf��8�		��Qt�m'��4�Z٘0���РkR��R@嫟1�^pj%0i�����D!3=aF�����1�:ʿ-u�,�Q��_TD���3�������5�{F��}6�\.�m[���l�O�W]Όg�]n��{gb����\JG��"�;��Dרe�X�i�! cj�N���I!9�]7�%CoX[N���M���OB�����R+~@P%��Lm���#w��Z$���XC���T�Ρ�q�s��s����[-4ػQy�+���Տ���B<�R<n�����{r��[$�[�P���Ʀ��> K��y�l;���� ;����/,�|ڗ��3w$"���W�8�,��`Q���խ�awu�͎�����4��M�Ւ��{�v�'M?uF�>^�:܀��ghF/"'s�86��o�/��Zvj���K�_��Ue�'���p�U��}�aW�,�t"�[V��S��1h%�:&&�5�����U�I��N�UX�>z>��I���=l�(�h�&�f%?��"�n��RsH�Ë�����yE��DV��L1�z;
��Qz�V�!�x�Sj����%H��.�60�����V��ͬ�%T��n�j1	��]Z��$�^���3�����8h!�a H�ԎJ�h ��������<�@�lF��V�	� �\)d�xg�ڷ��s$�[�?��"m;�;[�����1w�-�����-�?�8D�`IvL��v|wC}��ȧ����w%r�5"�@�-��!����}������c>g��k��@8'٤{y�0�H'm�o_j#��^J�Dtě��F��ub�=[�׎x��������6w����m�&ÜN6��U�$�Y�T�$���0�1�fh3��m��;e��A����n)��v�����R���A�?~g+$s�����ې����%�&v�؟��F�쥶W꾽t`���ގZ��:��9�N�$�y2AE�+֚[U���x��b�tÇ''b��cB��Մܞ��Hn���]�
w�pbe�)WO�唔ba��x��=9 ��L}z�{

����}�#����|20�o���l)����@:�6v^sg���y/���k�\�b���}��鉻j��O��%<��!�� ��L֗�"��k���A˪��͇�d8a�6�����J�_I.	'2�T����h��L����N��`
��I��~�>���:��D�`����+�/�:oZ��ۦ��vZ��=�I���3"%K6c�O�����+{{���S]���͂��gG�R6�BR��l{�2�iZ\Ӷ�$ �;�¶�N}f�;W�8^A~�tYr8o�>_�Z��2a���Ş��D�[E���΍J�=9�p؇a|jJS*e�B���T_�o��v8P��2���jB'%:x#�p�χ��S+�B���+���9�Ϛ�8��{,�A��ۚ\�8-�'����S���W�gR�)��P6��Bw<�U@_�����Ӿ�&j���H�-׭s9�7L�����ԉ�oB�B'��2���b�*������w�������h�����ϗC��%S��<�p��h��s�)����(�㪡���W���M�:eXϤD�����Y}��q�
 y�D�	�PtuP��r�N) �ݡRg��A�Ϗ��L|%�:qlz:��$v�����-}������β�-���2�+���6p�n�Ѽ
����s�D6�}z�>�G� n��&�L�Pu�{y]e {?�R�J�sasʲ��D&qk�Jijv�[�`�2��z�� �T�X�@�"u�o�:��S����S(������>~�:o_��ݸ�ޟ���V���($$��ό���vս�?���߻�rt�4vtFl��v�wp�C ������A�>2� ^���v��g���"�qy0��a���q�ݸ�b9@MiΚ$Qy��삮#圼��?���E%��{�*��[oo�`�:��?֩1��U���=k'��9MQFS����l_�(�r�D�g������ak�{�uP�}�z+ 삔����0)��Fj���kh�k=~�����jK%�[%�B�a�C
qy�3?�&�f<?#g��pc»`-����y�&�[V��X�\���/���Z�n��]ϥ�j?��D2
7��V�kwZ��E���i&�EWl;{{G�<!��,	O�^��9���l^��Y�Y\�4Ѯ2r��mL��8��%���v��H=~�y"�G�>��\����q�L\�dR����=��F��L�!��;�㩆��q�ؓ�����W��P5��Dا�O��/�>y��f���x?�j���4~ʂG7�{�'�gS-�������M+����X��յ�}f��뮬�����1'�������Ed��0"��\(�& ����I�*�1�����|�!c���A��]�J+^�"So��z���oN�G���N� m�8��6uY,n�rc��� ���!������U+Ĝ����E-Y��;f`�u�p��gqi��m����qj�sJJ^#���9d���&E�����tH;["+�X+ҫg�c~�z9+�)��6s$N������UPpsi�Ȃ{�| �J.�!�ǣ]Ru��A7��ܜ�+�/ ���Q�!�K)��gP���S/�ۍn`Im4�c�̙��M��U�����*��q8rK��n�������2l-ڐ�G���m�������.�_JK�vX&�li���YpH#�sY��`��pAʰ����޾g�Dc|�n(�-@d�4��vߟ�˞��ܦT\����k{����~�\������Ж� �:���Xh����5����ǯm�8v��&'�R*�[;*6�)4��^�y߭6|�������W�$�ٴ����o�~�Ɯo=�C#g%sx�%/��B��r�E2��KA��lq�3���DB�u�2EI �L�1ēU�*k�8�Oxuw�F9���kRIF"�����[(�q���C$�y �^x���0X�(�o�$������F�q�֯�Ǔso#_�)-����ϩ����%�KN�?��7nE�Eg|\�[��(m�oOG�$ez��/pa�@���<�0B�?���t��|���7����Ʃ:I�����9�(��Ɂ�h��o�>�%�Х��9����;ͩ��l��-֧<&8w�����S}q7�C܂��G�A�h�玫���&GLNjG���,����/�#�0���ce�R���uT1�w�P��e��4H��l	z�S�|�U�Q�}PѸ��6/�m2Q��t�]��[��׫�{Ñ���*.�2᛭>��`��!�����@t�U����=���28�?��$�X�4�.��"،> ��jo�*��>��Vr�5�a��GK��`rY[2k���%C�jtP�R
�E�;���+c��'XF���2�N^N����wz
F�y�Q/R/<�����Y<7����7��Io>%�Ο;]��:@�Y:�����U��7\)N��_� �Uf"��ͣ���[��YdՈ�� N��������&�[�6	1�^��UX�j�Zf0�, ��.��,�x���-�=�e~�lY\
'��`�����y����-��QR~)�|�c��C�h�������# G�k��ע���E�����Qa-D�����wB�5�����l����]����<=ۍ�$�\za&����Ї�⡂���,���{RM>�:���6��wdO�=*Ʋ�7UK��F��I+�$����	�d���iZ��)-��$u���(e ��Ǿ|oeW'��j��T���z�^����9��d�Z��[_y9?�|�E}�V���t=�2�P�Z'���ffD�Qܤ�+�m��ܻ�.���]���<)�/[X/�yu-c��`�e%���;��P���*����O��g�<�6�[o���a~��KO��1��޾�%��i:ˉ�ݴ}�+�*c'Ǔa�!"�}�Jzp�RbK+�0��@R���g�rd}�;�nـE+S��j�>̛Qй%kRl���u��ɛ�G��ͣ��%]�����]��s�A�1�rf�
e�n��J��0�+�f�w�:ȯ2u8�.#hIs ���ae:I�Ӧ-���ѹ�kLjR�}Cn�NƑ\��k*|:9�b]S转�R��s+Ftr��M��Z {�'�o���b9+o��[yޗb9f�ㄛ>�����<\��|�F�4?�X�钘[�F���ӱ�F��V��Wp�����0w�
0�j�Q�O�hٍ#_���&�D�Y-�*ܦ'ꬤ]�t.@�[ϋ�y��56ƿ苘���3�X;���'��8R8߱K�k��,A^�J�XY7TdE�:`�N��l��n��ԉ�`LM��:��R�#E�c��������)*����
����/�m8�
�&1Jܿ?Y�� 4��Z.���DbU���.��`��p���fs�M�}��Ϸi�By?L����y�`�i���&/�oWeV#��m�M�|/��KH/)29��!�d�n�|�p�����*[�&+�q�K?׫?���L�s��������]m���;���Bi�|�sU�	�gUx�Ŭvh�E��KX� �������gl�L���g�A�Ji�#�p�}��	�
#���t$z��6���MNf���k������	5~�;��r���r�wE�~Ce��o8�)���Z&��zr��]����h��R=���(�k��:0�1�?��W,(]u�8%��T�Y��楌���A����ԥ�T��R�f�4-�����c^�4_Ж�yc�K��l-�t�e�#��b�u�t�4l�qtΕ�������B7
Ϙ_1h}�ˎ�F3�IVp	�q��q���Jm�X���4�"�D�<��1���-�I�wez�4O@�>����o�1�k�<��RMo؏ 韲�����o�8b�k#���oJM�VS���5����2S0.k|�W�l4�3>��͙r���nq�>�U{��ӊ�pi�D*���o[��r��u��<�
����Ӏ��xH?���B������5�;�p>�	p����J��s��f�a�>��>�>�
-��7_��\���.�\���<i8�^ \b|a�$�3;�f����݃���C�I�;ĭ��w�-!��Jd��S�gi������.���~f͟��9�C��G�8�-s��a��_���s��K�������WC��g&5:�#w�*�wJK�1��*�N~�1q=��#g-�l���v}����lg�6=�Aq�/���	P�m���� M͢�I�DV�R��������RWzA�*M\6����ڙ]O�kj���#���KM�L����Ѻ�r��ٱ1�0�����:\���S��c'� �U��@��3�������D����͢�r,U�/
~BT����+��{ᥥ�z<)}�]iaSk����6�!y�ܶp��[c�U�3�� � ���ɫJ__��*{���f��į%$�G�V�l�E=��$�^u��װ���zn楎X���'ykc~��s�O���c�$g�7�E�Jp�\�}����9�R����){�í�qR捚�n�G~��f���5Ry��q���.Q&f�.��q�쮥��Ͳ�]������ͺR� �@�#��
�u�J�jll�g,ee��k 9D��8 �uv���e*�>�a�����FSV�QN�>|y/G��ke���pF�'�Ȫ�.��õ��h���v>���s��^���@6�0P���״E��ۻ+�-O��+����mg��Z���CTίDVh��d^<e�|�\����2�`�DGCi�#�{�%M����~?uh��8�ч�0�~�>�B1wT��v/���]�?�"�tI4C��?E$�6w؍�d�mF,��6B���f�-α���>�b
�w���;
'Cֆ�Խ~���hB�v�T�O򏀈Veg=�z?����V�� �?T�r#�h�<��[�t�:��2�E�YN���@����B�et�]����Dp��=�}ۆr!m�t�> ����� �k�}x����(���C�5ϧ���՘M	~U~�����w;F�*<�6��S����W>�l�L���O� -�ה<�V$���I�g��>��	gx�2Ⅱ5eߋF~�A��;���7i��@�	P�W�{��B��!���])F,�0����K�?��>457����T$�"�'t�`@��j����ыV����
����I��O����`���f�U��f����<���	� ���}�7�� �D��Q�͎�e�Z��j�s�%�뼷�@]�`�4�
E4���?������a�W'B�̻�2�V҆�����[��
��#4=3�)�^B�i��S�:�y�����٬?>�Q��f��c�Q~ı\��a��k���㈕!�95�(Pp���H��ѫ (#1��,�'���J��955�H���ީ�sG���������E���g���I�
�"�%7�%���+yR0�F7�=/aG�]b_�1��}Ŝ��T\G��^�$
��,��>ۏܙN��QRR���̏�4-� �&))I�ר>�2o�cB���ɋ�1#>�3�+��� 5�����^t��o�tGϱR�P����7xi�X###GVm�\���Ѓ�tG�t�U��ʕ���5��l�?��v�엛gzV����yW��"yh���a��6)��e`<���R����1���iæ���8��z\�/�""�F�[G0��Z\�]gv�rM���{�w�o8>��TB.��������4F����?���s���n}�( �D"e�[����J@�~�,�SH��;M+.�BfC�jZaT@0(Ndj�g[�M|����ǹʤ��Fm���R����W\�q����`)ަ֛�a1�Ut��j��ι�<^*`.RO��L�k�>/Y5 �܌��&e!�x�Z*&��Ax�~�`K��q�M��)�ˤ���?`� ��Ǡ
�M�v�z�_:5��h~	��	�X��~�ؗ㓓`M��
��M��x��1��Lw�t��v=`�\=���=ٹ���38׀Gz�/y��� 6���,��B
O�v�!��R;jɟ���ʭJ�Y�[�,c�Kx�oϸ'�Ç�*<[�ӟiqQ���S��x�#�{^�Ԍĩ��K��,��E2N��^ ���~=M��W������������������AOO�}Ng%�:�hV�o8*Fm�s7��0}��d<̺�Ho�`m��S֚D|k�O�f��;����'�e"k�:���"����듣߮�I�����Y�3�IP.��:�֨��&�}��>�
H��y ��j���&���83�kHF���ο����@�~w%�s�,�{9���/���t�MH�۫�I݇B�`ZYV�g��glvd�k>=ȳ��9�����>��lM��fQ��(x�Hْ� �6�$��G���J��G��O�5n��"�%o��G�"X_�P����t�2|p�M��b���d�p?��bw��G�l�Y�%�~�(�j�WʰD�����#��y}Q�~9�!	s����)����ݗ`Z�ĺqj��@���7���w�U��fejI�|���Ȝ�ؕ����Y�%�(:�(Z�s� ,�C����s��.�%QZ
�i)��d������t����&)ŷ�P�g�l��?����_U�	���G?�	��!�z���hܠ��1I�I�+)|�Ex����9��~ş]-�r�Z��+?j�H«��k����9�?��|]�����y6�s�O�v��48B��MA���R���=+�{��b@���~�.x�U�����`��&It-���i����fm����6��eq��]k�,K�wZ�y��y��r�}^Iw��Lw�KL����1�����u��#]�𤐑*�}
߳*nw����bd��Bg�x�̹ܽO�Q}f�iU��oB���\v�î���i��	u�3��w���w�
�~��ݟ�=���J�����<�yHGI	�^��#S���X/[��q�1n�w]9�F9�{����%
z�>/��99Q���M�^k7���d�Uu�.4:�1H�w��Z|9�-���"�k��Wr~������g��X�48;�����7|2�pX�v��3U�d�MIc����ѥ(��W�����G	�@��<;zR���u� \
���@�S%�;�I�/�5֒��A�V���N;c��)f��ۓT�GR��m��+F\�9��P�>@BI�D�������nPӮ�nbc����N��D�&�ɪ4AO�g��r��ư�������ļ`�s#�?D��%uR5����KS�d��d�F���^��F����6?f�H�'��p$�P�Ko�;2������5"9�x<q��6[}���/R�	�Q���~M����ȧ\��y�1�ӓ7��q���}��ϗ��v�t�M��������¯&�]�Hjj:29ߩ'��R<�&����~SZ;���E��@}u ���G�iJQ6��| ��0�>�C�#������רe�=�M.J��W�p ��m���Fj��KJ�<� 4��i��^+w�h�KR{ָ�W�F�yD!��,���
䫲ˁ����G�q�Ձ�p�9��q1 \��jd�[�M'@����:: �����_?���z�H�8�^z�PMT�&��yi(7��8Y}����"t%�>�� ���G�hkgG��r-�0Ҁ'"_.������g�]��(�q�&$���ݳE?DE�Qv�i������9X�6����<نx�y�YBP��O�.�+�5����-D�6p../���mҗ��<�����)Ӽڱ�v'�3`'��g���nJ�/H)�% ����g^��74�A�K�8^�|Y���2��eN"q�Lשy��,Ϭ3�Ń�^!��^�75����*,�`����tQU�	��o-\S`���ؑ3����AB&H��
&�8w�`Y7��D��6)�@z�{	A�]� ��^���@Z�:;WQ��/~�� K��B`k�'k+^�@y��^>����[
���3���苢�mrͯȜ� � %F�?��6�	�ej�6l!�6��\a�4�і�܋���A��&[�<"֘_m�_��A z U�w����h���8��q�E���ӊ+c�w���v�'D��]�u.G��su�r%��b�$���TTT���H(&���>N��/n���Dnn����G?<�l(��opx�:ǉK�V͠��+��oe ���0�CH���/O�s�W��� �}���H+�w0ή���'�H�o@����]��~̖E ����5�M#��K��X��;�`.ʞl)b|,��櫒7�צ|�� B�ݚc<ĹwB�+#�۰�wبޱ���À�!�6��u�U� �m�$=�'O�]+15�8w��QN��*Ӕ�VL���W��nsS�r~�b�����	��r#�y
֮�O�;�Dq�>LSd!���7*)*~+-���p��u�,���m�3�������aV3�����~@�{�7{�a�Q|�D���G�#�:�؅w��3���;���\4��Lx���*O
�.��(ښJ2z}u�Ϩ���*[�;oC*���:��'�2�@כ��u�δ�Ԝ�������eϩ�gx�����'�ϛ��[`J�*a*�r�@@[e��sL̳k^���l$�,�p���})J��'%Î��򚠤"K��\&W���e�v�e�:�aO�n��pt���˃0��1�Pj��(����vd�Y���d�f�2�L�8UvV�'Ϥ�����[X�أR��د��Y�@tD�^eo`��%K�O��>��M\*e?S#�+:��_�a�S( S15���F�#+��9vf���Ne��n ��?,���n`��3�Q�8"|�����U���2�t���w55��� j6�L⋓H������R7h/�Q��)B�0p��%��rb���/�v��#�<g�g}FZa�p�/��sa��dp�� ���|jْ7鍰Pu����q�bY.���F�� Y���I�=���7�Q��p�&���>V�'��#v��7�%�\�Ƙ�K�)F~O:��xu �`�71}1����{�,$�G@���9���L�.k<I�������abw�d�I�,�#�����sT���'��V�W3Pr[w[��"$Cjt��1>�5�33�ɘ�<4�\h�,�.�Y�9Q�W�j)������{���#�O;��/�xsW�ՠ'q��͒�p��!:�]�S��}�}Ⱥ�r��X�0.lκ�Ps�v��t2��;��A4$8���B j��R��e5#c��>������������h3�p7�u�c��l-�%���{u�� �����?)�W��K>iomk � ?:w��*O�DP�Ҧϯ���&�+����@�Vw�O�E7l�����T�nf.�xNi�4�l�+׉����������{^ׁd�6�'5��q3!Z�fV��ĵ��/�-����UUV�J�H!}��@�5�����>�?����{������!�9��;V�xR�j�-���ޙ)�¼�?@�O0AQy| o�@I�}[��9b14+�ifVh��X߇�R����4RQ�br������%`e�ڡj�X���>���A��isHK�z�uv��O�D ������!e>�e� ~�DX 
�j]v<o��5)���\g�����y�;;�c(q��to�9�����"s�jR�����2�H׻hij����a���OK�Fb�������K�〠�V��ZH)�j]�vzͱX+s��dg�^����jvlv�2��|���9_{�b~7V|�+IJ��	����O�>�Y�fP� ;r���X�M�C�c_���K1_N܈&���h�����i��?-N�\Q���:�f�x}�3'-P��l)/e{��ϟ���P�T<�3�,�k���E��K~"xPh¢ޡ�Nn����?ѸS+� !�O�[�Q�N�"[ZC�z=�����x�B�E�u{Mc�V��=ܓ� ;;"Jn���Xg�"�W�f-Gڀ�����]�L�M�"'��٠>.�J�}�Y?c6Wk�_'1ڤ^���r�M	�ڱ�� q	�;���U��vF��\Fs�p(����~�62;R�"��d�>�,٦�2�qX����l9d��JN�f�mE.n��.�+{Oh1{��	�:n.�W��ȉ���T�`����MO#�z�P~�^M�������_�Ib���?��Р����3>�au$Dio�V���<jA_�}�APU�{O� �����+@�3)����B  ��=��:fJ�n�#��cőm���Y���.-)��<���Yկ�������O�Q���D!�*%��/������}y�3+n�>�oa�/�$~ �b2{�<��ї��an&����(��__?dO�2�>���d@&���0����u��CףsIÜ�@�����K�L��`��D��*s�J��+h�W8���h�9�hw^h��`��.c��k,ԿFG�ФJ�\q��HrE�Eڥ�P(�ŋ�_�͠Qmf���l<���'��g�#�77u8[u�Y��y���)�r�����,zQ�̶�����*yo��"ʾ��e�ƏOTS� ʰ�0��Q+�\Gi�$cNi���NZ�G���LI��~˹3�rSa���)Fv��mktz�ƈ��XXXkF靟� y�����y����T6��~un+c��$#��wL������ߙ�3U�������
.3�� ����$���$�J8��B�=� ��Z8gSJ؃R�:��܆��48�$�����|2Z��<��k�g=��6�ת�^�����w�<\�?՚���t�t��1��^�^��$FI���,o�O�9X��o�~C��疁�F�x �nT�=Cߘ'����l�V�ȷFI��6�<15u^���˔��F��A��{���ߩ/�i���jUDF��}rV��6�/��.���J��\��?�4li��^��A������&�A��g+:B��jX-�j��KJp���Fn��T#�ؖC��9Pk��P�s��ݕ��\��)mҽr��'+�y���:��K�D��7�L�s3i�;����1:�TŎ�7�Ny7 �S ��Â4�U�f��Lj�ad��(�����V�a����);�4E�9�B���[m�υ����2�A�Ѭ��dHd���%�C?���E�F�+�2�ۛt{l��^rL
b�M�%k _�#��#��~��xl;�Z��a)��Q<$;�ڛ�lY����_���y.1%����lF�� xܠ�����AH.0Ǝ��0�jۄ���V���>�+s�Y�ckS��;I��׎�s�����m�n#����� .i̓S
�#k����K�O���%�i����n^�,�� XI�|�k���2��q9���
�R���%����2Si�s}2Ӯ���1��Up�hx�-��u�n�q���f�Fӑ[w*=/�q���1"��A�@�x��9ZW��;���iUx�<@}�I���eF��R�յ+�y;]��U2����`!���T���*��_\t��
����'�!G������1+�f�1�w�DJ�����xíY�zA�n���!+����M7v<�h+�B1���;۔}n�Q�Y��Vz# �eQ��00X�pՒ}F8x�N�bP��"y�g�G�)�8P?��ʯ�P���w��3�x����Gf�!,	�̭x�-��_��e�,��R����/��O���i�c;��}��>��f���ۆ��K���<'.e���}f$�Uxjl�8��b&`J��s\���b§h+���is���6�|Ir��K@�~�ծ�u�b^��"Wt}���N ����"n�u�ү�+e?����Ƴq����
M����@a|rr����Z��OD�pѼ��d Ю�
�ŉ+����8��i��]Dc���z��5T)j��º:2 �hŢ����FŖ|6)$�|�ޚkU�262sFHHh@����?DF}L��lz�J�1
}�%�$h��{d�F����U|ҪU�WV#�N����ӆ"j�ʦJ7[�rUOa#�LV4S��g�w��5�M���a��'��,����ՙ�'�G���[��S�7�J82���c�{ݝ'�7��@���5ދ��G��fE��b�o^n�'�N�n�)��&�Cx\ۘT���e,���B޴�|V�'"#qێ)Ș���o��7� _4M/�/��o�󒓛�n�=̎M1�-���ї>���G�8�Ie��J�߭���<#��{B�gg^ 2�<��k{D��Ĉ]ڸX���X�K,l�=��o�I@�M>P��syB
o۵%�D�d�����i~�c �Vh[�g�D'm�p�q�7��U���7_����=�����P)�k�{o�`H���0��#q�M����ǡ�����ee�'��'�(�ONV���n�	.=�W�8�z>F�$YD�k�ˊs��������F�X�g��}�t�m�9�]�NjM�Jee��J.W�$��T�����bͬ�c`?�c��֖��((vܚ�8Rm�
W���?��:.ʮyDJri��.�i�n��i	I��Aji�\�\��߽���������>g��33g�}��}�������\R�d�M�䶭jl��e���ܭ�"���A�Aqq�e:�]� ��/[!��# E�� `��{�E�(t����d�t�c��{eǢ�x�8�j��'��Q�ڄm�͆�uV�j4�vIZ��w�4w�:�\�vKqI(��;[�.�!�񺻻+��ϷƷ�m[7�[6�wτgX���^ɱ�$�?�/���xD��hq�� IM�`	��z7�c�J[���[�>>��	�/���:]�����+&ƿ`��� le��~$W���g
~[lþ\�a�0A|~i���A����ĥ)&�kM!�Ա+��Ĉx�X�����à��81�#��#���������I��`|��a-däw�MKklz:������香䡷c��ѹ�O���s�;w[����/c�K����SKВ���������mQg���m��ؘ�~ք2_nm������{_͟�rD9�y�;"��n�9�����j��VGz쩾R�����!���wd�'K���w���l�#������#o��3��|s!��޹6<=�!ܽ*�0�y{O��u�R�>�B�M,���G��X��2��ư�3�VD�=sc���j2�w�#+�~2p���ϋi�M�*�(���ؔ��VY�f�`d;���>��Y�<���Z 77���h��s�H?|&�<i�6<�?�UF�T�K�}��h�e&��9�����Y:�O��6��_s�&J��Ҭl=�Z IꝎ�&��T��1d�}Ϗ��!�C�mv� w"���^3�^�P�D8{y���,j��4f6�$p�JIEճ��l�'�PٖT�0r'����
jC��@�^�����)u�}�X���a�T�)D-ܴ��B*�ekY�����<��H\�*�"{#�t�RN�@��VՁh�ӫt��a( y|O�K��=z��O�G�#��:���d�x5�Cm��t��� �r���J��06�p��7�;PDf0-A�?�96�b^/OM��c��?>�hP�	=������Fת�t֊[Pp�q��w����Gu��<��2�)���k�������G�R���y]~�����yz������R��v��S",PT����B&��8]͑���^��= �&��ݜ&.q���eF�ԏ�P�M�qB��5�3���N���e�EH����ZL�|��_�,��l���@B�A��|��R���?*s��T�xj�(������.���7�]X��/;�����x��
��iIx��|�zװB"�w�3�N�1���9
%�/k_�)�����TR_3"T)E}&=b4�-už�\�(���,e�1�c�Pm��	��r�������)|�Y���OZ�.L�A��D-�H����3k��2�Zt1]Y�|��ʆ��w�m�;���r�:���4v�,���y�:��5(�Y�w�u�� wE�ު3�R�B�{jؠ3�I_�C�����d�uF&��㟦?jF��� �p�=*���*J1�n�5@��q�'��s`�l�f��)X��(������ � �#[�$����yt>�y�~w�{V��ߒ��]�ɇ�
��-7��B >o�GW~���I�ȫ;��u-Mx�%���1T]�z;��_�ߝ�ꑑM�z�J|��I�pm���p�g�PӀ:��a�ԡW�k^�lQ_��#�\�*�(����������f�G�� ��O� �)r�\��Q	��2 �k�v9	�]]�n��r��a��-�CO��njp(�g.�$l��M�����D9,2�x�����vԸFjB��v/_����K�{�ԅ_�d���P�,c��tKq.�[��/��b���!���w�*_�x����i 1ε�4S'���j�6pJBb�/:��݂��B�|J/�\P��9Nޔj�bլ3#I������7�����o�l��J�����t���h,����ʨ��*))	LF�yy) �e��ա+ۓ������P���K����3.�����*ec�_�ֽ��_5���kX�|nL[8?2�'>�L�ˉ���հ�U�q�<��.L)�IG����1P�=��D��々����ZWC+N�v���BKX���-�u�bj�6�{C�$����C@2*sR���ae��{ey�{����HB^Pn�`���Q��=���/I:,Sc����۱�����p#Ɩ����=�w����Ae�ws#h;3I4'6j�+���.� ("� �<��r|�wxs�wts�����x���\2�5��q*Q�𳕦�-H�����5�ܼU����^�+��&���TH��Ay��O%�����+N0���:� ��\?"��}s��}��	J�;y���wM�B����us��p���P���xTD�_��)��6�?߀��z�8�����l��]GU���!���m&�O̱�&�^�]!�#�cv�܀�<%��:��h
����
����e)C�����zz�z�����o���I�w��+��VQ�R�W�
"�g�6O;S��x<;G�.�O����mZZ��ȫ�(@\�=&5�/x���:�t�����Qa<�IV�����Q�zGR�[�&K+-���_�ce�x����46��͑�:\�1�f��ron
�cܕ��@��=����c���ʤ�r����^v\��ԁ[��=�N������X�[p[_�4}��m���\�Zҹ�?T��
j��!�+d�@�c�7�8�w��C*���nٛR0��c�����ĳ d	$2��n����A��|p�e��g�\oaut��V,�W<���׷�z�є�ͦ�f+5����+6�[}J��6d�'pr
�GE�@�DF�����Y�P|�E	 �k<&x��BBQ��\�,�N�;(i��R�挢JD/ݖa�+,$o��u��9�����6)u�o��;Ә�B���9) ��ݳ{JJJ�E��LO�[�m��9�����m�����Js�>���Lcֲ:�&���/3d�r0�j�Ve#��ۗ�D����^��Œ`��ƪ��yd��W���j$�HǞ$�0u�WՑH�	i�cF�Q���t���-}v�u}Ja��D	����/����E*Z|'��I� ����ܟ�y���U;���rگ��z�8$��TWj��Qq6w�ּK����k��G�e�dy�e��Ɣ��ay!�@��,�_-�l_��:V�e]=t�9nyUu$��<���9 ����p�E�ھ߆%9��G�fnrMF�uz�a�Ċ�˦�=r"(��K&\D�%�D��|7H��$���Γ��qz�y�q�n��w�N����=�B�ÂG���y�n��.@�*]��P���b��#�g�r�#���Wy:�w�5�7V\�p"۴W?_��"��9HC���g-�W��\��8\�I|����Q4�Gw��ͼ���P��m/����c:���������' F��1P"O_�S$�������vũ.{Z� �[�̨�<(��<�5�� 󌈄�T�/9�
Ө,��wR?{g��M�	��V�Iw�Z�aF:�w�͂�%��Yʀ�IԩK.��^�p��|	w�z�����%��U��b�g/~|��ׄ��W+儮UN��x����g]��C>�Ð���'��OT$պ|���ܬ/�*,��0�}�tN��2t�7�������"�09y���>8�]��$»M�w��@5Y�]x�fl��Jò�����[����w%sQD9�G剔Yϵ���������8��AJ�Y���/�8�g!��|�I;���� O���r�6{�c��� �/o<*JW�G���9{@�021��r���e�5�Q 1ƅT#�k%�QG�	,�@a c��B�������?�-�i���5������E��122r

F�ӇH?v��|��ђ ��C4�9��s��Rmi���M9qr��ҰW�|c��/�W����+��C����/G-�}���W��lm^�������Z�3�̲��LN����tZ}J9�Lڇ���CA� ��Qa���[n2ޡ��-]Y�l�mӰ,�e�M.ȾJR#�Ng�᫟��ߚtX�T;J��v�Y̭(�Z�Q�udֲcx@@R����@E�~ć�B��)3Ya���	��"�φ�R��2�����H�W_e�������<;zq�C�;���G�
�t��ޅ�n/G��� �����j�?!��"�%����s�\fnwk���;��h��0��>,����\��� ��{+�d�Ż��S��8��0��� ʽ�D�d:F�z��Z�3���~)Gs�����臭���	G�l�/ .Y^^�h!!��_�)���j�S�gL�4��OA��c(i���2xb��?7j����Mީq\�=TT����N���?�8������#`��L@�4�Dx�ȗc&��;�D�R����W���[g�Rq��4ۇx~+�����M9��9�O�5:��3훠� �м��CcX^�U2��e����ґrqS���F���霜AnB{���S�R�VIV�R�W����g#7w7�$;���6P�$[����VD<߳��u���Rc�(SDE�Ë��%�\�޷�M�4�����f����T��v�S�k\J��sY����ӗ���-z���j�J�P;���AD�u"&�)�_l!�Hl�})�ڟ\��锃���qpa����Im�Y���2rmmb1�����(�$h�������uuu���_������￧�ʤdB�~x>�;[o���0tB�7:�NF,�w�3KII���l&&#+�R�?l���;>�b9~\��+��へl�"̹|�c�6ť�7��l��hd>qQ/e��+[�j�����Ԝ��$��#��-f�X��5�ӷ#����7��K�sSSa��k�L�S���,�üPzqR��������Pd��P;N�g�}�p�o���y{��T�z���T�p��4NǨ��}c����/oF�K��D~ ��V�f�:@W�#9������7щ���)-e��B"��od;��bm ����bN5��7�}d��Z��l��!&>�n_����+�c�S�����@�ŝ;-���m��fڥZ�tZ��Y�kA�%���l���|T" ��k��֣�Wr����Ծ|���]�5\�]!Q���ڞY�n�ۧ5p�S@s\�����|!`�X�t\P�	Ä%��#<��_����ο�К;���W�=�-�5���7
,�;����_� �DF>�p~�d0<���p>��}�!B贘�d:��)V��?�Q���ˎM^��膁�O�WH�/Ê�X@9��*�X��!ۡ h���G �-��^۽��Ѷdُ���nm:[!�hS0 ��&�S>Z��Vs���N�oA,
7mڗM�G޻����8{��{�S;"��ܻ6��N��1����z�$��� g7t]Q�qYq�V� o�
�VY���3W2�R��$�
���߹��疔+]^Q-5�%�,���[=� v��vq�g!Z�f�������yO�iR��#��ĥ��2�5�f�D���p�`k˂&�+�O�x�D|�v�q�w
��� O 4ߴn
aܩ6���{�9X![�ο��n̙媾����6\��	x��i���#���e�q���Q����ކ[�I-u>3VzFr+=�#��Le��ke� ���ŉ�p| Z)�T��{��  )k<���Hp#،_�%|��W��w�؝y��um�~���?���Q�~0��Ʀ_��[��Nw��縻��/���y1���k#پ�'T3�5�����r+�v���D�K�x�B���?Y�%ȣ@�u�JVl��w@�����`r4��TX�	6s�	-�8�:I�����{��	�x����
{������P�:U��l�T44�>�F�oq4#\��ߤW� ް��U�S@uX_"��sF���rG'��Ä�����\gbe9��>� �B�H��`���YE"[����`��Ry�=��٤��ó�K���~m�����T��3@E)�-/Ǜ��yC-��y��r��0�I�j,Ꞩ6V�g��Bgp3}z�'��\\\�g+X4l�	vN��_b�<�`(�~�kS���Q!�ڏ�3��x9Ua��q8f1C���o�)̪��-Ƅ��ݜw?��F})��&D�:��vi%�а;�G:�Ht�0�]�]��
�$;L[X�]p������@���&�OͼFg	P�������Zy��{|�I[�A�h��ơM��p��9���Y��(�z��L�� �F<�;���mr���t��sC�+X�w���޷�8Rz��r�����r�X��7�������A�\	)�8�ٚ�3�Dz݊" 	ty���Z9�rzX��^3).;>7��[_��A�u�V_���ҩ2	.X�F>q�xe߂���o젺Y��QAm'P�L=��%ENk���B ,f�iL�y��9\�?�?�F���7=z�����#o~�{��^hj� ��7�|��hI%��vz���7c4-��>���\�����'��c���s��V��wo2.���T�y�����#w~	<Y��S�o���^�P���D��� ~E&���hvu���\�:���C�L��읉Gi\vE5�u���M;�N5�y 
 ��@,@��9Q� �Nr�C���>[z�h.�-xBm���f|H�`�F�t���qD�>n��ӱ_��,�>ZAC��ӚVk�J�;iuW�<u����&1M=1���� ���ͤ'�xss3��dbxd��-L������];�9�b��r�$���otݏ#9����ˁ��G,5��ףo ��7	k?�x� :�����H�>Y>)���jkC���K!w��FC5ڴ�\&���I?��Zf N����_�x��C�� � �����I�ɳͯ�w4	��^�ت�x�7�*q����<Ef�<=s���vn���_�n^�z�)���<��c9��d�<�y9���TdCh�-)�-�F�<`	!p���Y�Q��$�:V�NR`l�l��ђ�EV���!�r��wD	T���)��0�P]�ޅ�~:t�B1Yi��$�Úr���g#.�un�ߗx\(�xq�Trd�����#���s����w�n"����(�L$*q�^=�z�E�ƕҪ)�#���-7�QL<�� e��X�]�19�NZF�NOñ����'y��d^�]$־$��V�]0NJR2x���=�BqE����ϟ?i1_�:��-��	{̈i�cw�)&�~�n�c.e����vk O�EO�5�X��!��xr�1��[v��i��t�T+��/��?il~W�3�}��t��u������9��o�����Tw���:v敭rվUNM���r���K�LR���{[��dT�ܚ�Y���E�G!��D��E�]��|��dm�ce��fp)QG���z~��g3큁?a�Y �XY�6�M�s���R��mm�YYYʯ�볈0M�7:��Du����
�ch11����'�CUT �X�&WĜ�K����߆�L��_#��-4:7��p�U$t���V/]�}C����m������׮�J>C:�N�6uM�O�|�hp�T���|��r�pS�9)Heq]�x]}�Z,�R���UZ�!Ӻ��e¡±�8a�p)�4��ϯ�~�wvv��T/�_g�J��f���<)((H�a���!��V\�|��ʏCMP�q"�M����h�H�%	�Xлo�ٯu[�6lJ��!~An�/��vC��x<�;�C�.�.�?ӊ4��jD��'L�<܂Eoy�6''m�ɱA�Q �lG��c�<��-�Tچ���L�)ljbTĮЂ�0�	�yx�d�b"Z'ަ3��ş��c��0�Xh��̠8�4nfk(I����p��ZXE���|�� e�Q%�F{�<%4@x����A_��}�u��\����_��J
�)�=��7�kF����h����9��w�S�=����]�(�z�Я�0����������5���DX�� IWWO<��� �6B�
����'���uu�^��Ո�r<���c��)�OD̪u~��F�vD���yq�F�}L(�(�/؜'o^;	�i����j�m5�����`K���M�=<��x���J�!���B4����R��g��V������+,cT���@w�Y6��c��!6ωʅC���b~?�45�'&x�P�KO�"Mæ�-x�XSY����ߩ1Z���LYC��(/N�*&�Zn�e�]�N?a��+�DN��.�o˅@l]��>�0-DGG?�]*�JDOL��7�h�%3�������!�4�F~���~kh���EH{�X�ܗK*�2����-��2�;��� �E;P�Լ��MNZl=����*#�Q�h���˶!����ф(���z�h�v��r� �������c�D~u��Ngo/�dL.�b�c�&�n}��r7髠����EZXR�H�}EN<=�+�L��-|\1�v���I�d�%�Q��n�r���??���W5.#Z/��*hr��=�>�޽�e%���~��n\��B2��cjj�!fHA�!�]:_���˼�r6&�ڢW�h�����g�m]���g�q�e��7�����|0�EE5-����g�*��r`��wڼ�*�,֬��%�����5L�{��%2�ٳ�W�v��.^dm�z�5]���$�Y�4�¶��,��lt5l5"�l�4%�q�����I�T��J�ǲuw�NS����te��B�⒭���7++&��ͺҞ+�J���}\�KX��<���«��B���w$?�rKD���(�t�|��#�i�]�Z���CE�8���%ܖ����X!����R5���quE�ћ��FNt�p���;/��K���9*�?X𕦆�t���4"z��$T1��������`�-FjjOd�cW�#旊�kX�2����v"N�ݵ6V�pw!ǫ���loo;��<B9{soɾA��%!����O�i19�y)�eV�#��PM�����읃��T���I!�B1��@M��g�ޅ{C�_烅�t���;��ˊ���k@)ҿ;S�X�8��X_�O�� ?~�p����ě���\Q� Pq� ��<X�XU��g��O�$���6��z/e��&蝭m�j�d�Д/�Y6��VA��� ��Ύ����~�A���f�'g����##���O�;x滀��4��\n]���T�C�f��uF��Ǭ�=;�o��$N*T�9����K{DXu'|��~�o�U��Z�t5:�Uuu?'p
S��Mx�S��ռ{&��ݻ|�-��gˏ/ �h �.,t��D�����W�?)����V��F�fd��N���m�E��]���A6P�3��{ �1���*_.������h�U#�P��b�F`ƁTE*�9��[6}L�V?��GC�Tמ����p
u���]����FJ��h�`տ�����V�?��x���ukb�f�{���{
~:r

�v��Q�H���-̰Wʟ���B�J����yRê�^�D#���M�3]�}�ڽ8ׅ�G�#��WO�i��'���(���S|�s��v[��}]��2rW����Х�_�s�O�<��i�% �&�����:�Ї9�c�̀xn��G�Š}�P��I�`Zx݃��;�Xww�cS�>�I�p)gz#$���P��l�X�rA�u8����E�������EL�V��.���toy>Y�!�/�d�M����Sx��	����`U4�J/ÚG�)��ԭ��i7�$MNN{��
d♳nxp�>%�2�(��>����WQmB�]~_:�*��-��6�
�N��st{��?�Y_ O
M�w�j]�g�)-�>*0��98�T�>� d�e�7�B Ȕ�+�88��F�*���с�=^|���W1��!\��7���,.u	ze7L�L� �J�C]\��q�X����i�ӌ��
�NN�m�{�҆ۯ���E�z��O��@Ą����9��Cy߂�@��c 4��w�'�mß�ȼ�c�u��eǫ9��g�3sy�Δ��اnH�H�",^�8���;P"�/(�I���+��S�o+b��и��<Y�U\��f�Th�Ȉ�Cp&V�HD�TD^a!���F���������0�#\B��N��EP�r%|-:�3�ϓ���I ΍�ϴw���픘��|WY׆�M�y�oP�6��[�8*�,g�EFr�@O��%�x ���r�,--�aH�o�)���:���H���\����U�FP+ ���6�c��� �N��؆�"�pq��o�C����-2B� �u�'�+�Kw���[.��H���+Z@;M�)-���ٰ����nS�dH῎�Y~Q)VS�����:�O�WH�|l�!-6�L�������|�sY�
z�Vxe�4�1k$�.;�"A�����Pn����~�^�J)�+�V^
a��aF� R��DEGlMe8	ļ���`e�4�w�N��c�6Y���Vm��it|R����کn�1;�� �6_o_�'�A�~cb;��+��y����#����t��-0��Ҁ�梬:���S��^?M��^��/~䥪jb�:8�'��`�0L�)>��y���:�>�g�qX�̔�ή^6��޺+�
]a�D2�+��}�-�tT^�$yzdf�@ŋ�<��H�z
��($�'K�w���7�w��.3� �E7�7{��fn��D5����"ab ����u(ryW��I狔�A
�8��8a�G�E��3G�p����w�% L�?F���G��0��Ȃ��uد�vq�p��X��1`��1��6�n�*���Pqs~d��2��>f����@#?|x��
Z88ڥL��(�E�s���m�%�x�j���Hgga��T�QRR�'����!Y���UP�T΍눨�4 -�TdCz�.)5ؗ���QGSB��L�-i��Ö^%,c_S!���-&3����q�lJr4?FNOO�I������!�F���&)~�����O�Q�e�-��(���7��ͼ腥� @�	r�yS����<�A��ϟ��P����^K�X�W�9+3!N��R�� )���S8�0�r°Z%��[E��c2(�ʪB��E=��n7����Y��J����sĲ��4�����*��â��)�п��
��(i���..f��l�"����Ͷ�� nplN��*����v�DX�0�󯣧L�$��ޝ�(����R�������d+�qܢ�h:��h�K��78(y��ԅPق*�kk'J�i�+�J�=޿���ZMg���@�*�ߙK&:���Pb���4�u�J�p
�*d >��?޽a`k,���9����0���Ha%--��s�B2���p�y����)s�ڍom�
T0�����B�_��ܷ?���K�}Rq"�6e�e��c�����q!�/R*U.x��3�.���G���ԓ�蒔�4�Dt����W��A�Ļ٭���و�XV�y��a��& Rn��M�FN>H?��W����9���X03��_^9QF z�S��k�Q���-ݡ �e>o�����~t�����iE"�+����3�"��ݡ&�>I�7����T�v��m.̀G#�wG��4�\HX����m��;s���7'������耵|.l���o��٪jh��߰�i�g�C+�}�e�C�M�~��3b�<G��آ����7���jT��Ը��_p�3`{!ɣ��K.��j�|#�0"���D�n{K'g2�·\�7�����!�\�_�P��n�	;2̵#�c;�إ#t��(�(��3��ӟ'n,����wޡ{ĹXbE��v&�|p�oƬ������0- �%�+Φ����|����^1�B�N����݌��މ�=g؞D6�>��� !ԭ�~.��J���j� ��D��Qe��H���u����,>Z�d�G�(�-M��;i��r�_o���T�˿���s;�=����&���UGP��65	2��,�wb }v%���G�p��:"x|0 ���VO:�;-fH.��F���eRA�@ ���s��\չ�1w*dӒ-	1q�o��Y�vD�Obe'p�O,�mT�=v;�l+-]��/��	�W�4
I�� �����j��إP(9�K;�e�$���w���G��RR�]�N��Xh�G\XYXj~�v�&�e���n�4�#�0b+�� �I�������V�wu�mǫ�H��P$)�35߼ɫ��v����Dμ�c�A���/�O�-�97��3|#�x��>h�=k��?9�~r���Sa�J�	�ODrΓ��&��>-Rc�O`f�!�u��eMz&[dQ��˃6Z�*�M�
��P=�(6���g:�����B.��d&��
�;��d0��~�)�w3�������q���7$�	��5�i�A��j{Q�W��S����8N�_�R�eO_�x�~GYo�y�j-JYV��pS0�~^�|-�����Л�
���JՂ#�m�0l��E�9w[V�Vk�O�I�$�[,Hԡ|X7��)z�P����}).fޠ@�:^�$2��a�cO���r~c�)G5�w�{)���B35]D�H��^9J� QKf�}�h��t���]����Z;g���������1"����O���fVV��5�2P�D樏����/�]��EX�s��4�N�����9 n.?���C�l1�> ?����S�Vpݑ��j�J��ULn���W:��p��W��[{<���F�cz�_}�O,�ހ�p�t;���dje�<�ު�5�����@��Ft�F���R�yY����g
l�TW�./jz��o.�`M������`�W)� tJ?3UT��		��Ox$⨨����ip4��>�Xhݗɜ��.�Hv��z�>�׋�%��יc�>"Ǯ��x�dԮo� ����������^~jɽ6�v��1O�r/������}<sͭ�������V��'��o�;�� ��)ߎd�{�V8�C-���s{�a[[S�#�̀��<�W)���b��?��|ٹ�8�ǻ���눎�D�D�,3�Sgy���	��uX��TA<�s��؏IX�ʳ����飼C��ỳ��lB���{w�����&����Z�4x4�oϽ� eo.����h}��3b4j**�m
e�w��f�_Ők"��Ë�j����	 E(�!���;;�6S,v��O���u�aa�rXGm�%�y�%q�W�9jܐ��z�G���#'�-~c7���RJ�H����BC�]Lu���{�^���/�P���zqp�pE�[[�Oɇ}D��(1��N�̱��D�H�7
��~��f6�#�@�W[Kx�p�5���tHQh��\U�H����cN�Aw��~-Ε'{�	�Q�ZZ�A,Ք2�{�`����swH	��@��������̔�V6E���Y�<M�����j]*���ū��U�g��g�7��w�Z��n�;@C�����4~�����R��S��2X齆@ �%�(T�����|��H]!�3Ծ���0M���>���&�b�ẗ��@���n�q�>�Bk@A�DJ�}r�~���ו5��U~;��C��L8���Jc^�;!>ʻW<�w��n�=JG(�7
6n��t�C��7��Ơ{n���G�N�o1ZW���3#�л9%g
�v�܌�c����A�n�]4$Y�0��}R?)4 �@��W���W���Q���ȲX 0X��f#V���@ {LM��ˈ���7������V��c�&S�k�o �hpN�Z��NS��Q��4�7�����g�>���2�`���k�B�hA;�
B�� NbMcnQ$�j`��b��3����	��������_���B3����-W��8?��ũ���:C�=���޺�&r�������������O������ZS���?4����C!�i�����p�ѹ���Z+�K�{WJ��C��̤��V#4�M�Ȏ�W��;�,����B~
�D�G��/hBյ�nn�FY�'JBU	���Ռ>���Ztj��I�:K��qT�{�q�ϻu	0c`�O��,�$͛����vy ���Ӕ4��e7H<������u�&/\I|/z@���P�I&��I���.W��H����X��;��cFfra���s�y�6�����#/J��.Rʒ!p(l�!H?��<޸�jE�
 ��V��5Ye5���!Q:���x�n/�E��L���)a�`՗\ب������A^OH۞$�9c��<p�Pѝ)���>
9��~a������m�\L���Z�u�P��I������'�R�8� �Ҵ0	� ��B:��$���2O�*\PP�pl�	�$Iҗ��8G�5�k��lM�t:��+�5�v�6��mќ`�B�6ʧ��F標oք����[�1�^��koś�[��vڢ�<yzu.�9�aL�_,��>��K�����p��U����Z?�^���y�$��~��~�L���H2��������C���� ���DH��e4X̎v���R{�����jڗ�%��M� Z��;���s��U�ײ�G��6��#?f��v�f���T�֔�=N��_�ˇ����m4���y=^9���� ^5��(����TU������B� .��q��m������e�'�;%��4�y��e�U*b�Xa���k��7���p|��ciԡ�0%�_x�:�=T�J���h�'hi����֭I|��H�E�
�^M��΍G��Ŷ׌�w|<��A��ۢ�j�%/{�w�Q�� �r�����Wv��-~��g��ǤTc�����z�e����j=������9�
�y/��|��o��i�ӑW�6�� �9p���t툙���=f*�I�闦j\�mϼ�S.д�ͮ�e{�P�}(�Ѷk��Kv��iB�l��AZ�U��AwTe�%���4�_`ʭ����U�<1���so��o���_�x�zq�@�l���$ZR�3�cBN$����&��]a3m���|d�t	?�@��J�WL��D2���js��m�^������94��ǔ1a>�z��Y��f�Ȼ~՛:X�㬹8�~Y�*�f£���S�P���$~Ţ�����Hg&�Ր���x#l��g6�����9չ����I��ʫn΀�s�����w��(����of&���X�O�j��-<��\D�� �'�F2�Ja�:�������+�)��]�5��L:�߹:��=�Z�Ug��G����i?�y�7!�IQ=n���h�dv���)�6��V�A��^	�l�E����.��G�8��1�k����I��|`oJ�8��`a�ȫ�D�Z ��u{:`�u�&��n��v��t��>���]!�0���I�E��`�N�:NfǨ� ����X��3��tt���PO
�EălD�_�c�z^e�`�;W�s��ω%W�*�g�-�o�OZq>Q���+~�WH�~���;�U�[�������g$�h�%�$��'M���U ��uD��ۧr.���r�̿9��&��L�Qݝ��	!.|�Ws��x��7]��wh>lS���� #�e QG�����4��D�9Hz���*x�M�E&��y�odL$s�'���]��|@�j�����v)���y�EVy����l�u�0�_��j���|=ɐ���L�{������`�Hr�`\(�ia;{�B:�*�0B%I�-�%����L'9Y�븟�y�Z�FA��,�C���)$E�$��z�w���2U���G\��4oS��CP�:ۯ�\���Iy�vv��h�!��Ъ�>?h�&�m���n΋��m��w���8r�t�B8���$s���=I�* ���x�Ch;vκ8���!�{*Ɖ�j<Sӗ�V9=�S�{�����{�Ö�Wq�F�_CA���^��(����
�:w�ᦴ���)I�5������j���ݻeM5�d��+�nX�}9^�Հ��^�N7!F�w�O%{�qn�s.��ISVӟC,�D��:�O��Y���Z�������H�k�z$�]	1k��ه��e٘q�gM�`圹x.����,�B̧��x)}�R��_&8,��Ŀ)sRwww�� ]5".�U�d`U�֖O�1�w�t�1��k ��9��D��ڣa�d-t�Y*^_����v�oiį����p��?��Y�^I�PiL���`2lЩ7#��/�V&��Z�cW,*����Լ�Ӯ�c7Q����'2G� �������5��@��vc��X+�F�[�"!JcN���Y�2�_g~�d�	����M��E������^t8�K��Q��_�3&�?����V�\�Щ���sW���^h=��6$��E%�|=K@��>���S$5�O��>�����v�-R�f�:��cy�>l�\�~g��^�#�څw�����Xe�K����M�i�q)'�6�;�>�3h�Jtc���w\,w�}g����]]�V�����'֬��̰~��;����Zv3��9ă�#2�[NE��c?���U� JjD���i�V�1���+a�)i��Ro�iZN�-����i>d��XY��qL��/��޺��38����jiC��iR��O�� JG��9�y��F���6�zwcm�׹j�~�~.��9���f�^�g�K�O��j%yj,��ᦻh���F�|o'�[�
_�{gw�l�xYj�d�7�g��n�F�n`��{�K�_��_�Q�	�2R�J.8u�T��mЏ�#��N=C�RjyV���$dⴝf�o�I+���%74����A�^6�v�������9�	�\kr^%����o��$A#'�2O�׫AE*9�4w���P����B2m���e��)n_��R���Ϳ��D$ҰD;�/K��Ũ0�������B�M�g�h�{�i��!��!e������'9�<8�4��h���;���O��m���J��L�;���A K��BC���͸��U���tt:�<�+r���#�\���A��k��#�袩����k(��Qu%�P���%{e_+��o�Iْ�Y��}��}/��%��}�E�3�}��c������w��s�q�y���s?����^-]���:~R��9��i�y?i�?=t^�\j�;ۯ�)ÿ~lL�ZT��iGcD�r{S�U��f�U�����3��o�G����� ]_�9 ����"PtwYK�އ���/X>���%b=2�}��r�g��ƛ�}�I�D���4�/��|�FX��N�)�x�m^�G�W�����}��z=��˟�C��_6��k���m�i�M�L��w�9��wHM����<Ece*9�o����� =t�],q��r��&��x��7��4	��$qAӾ������o� ���`���;��@�wr��?N�kv[e�d�[�#�]@����6���LK����JE�:[	%+�3y�EEEߘ��C�*����m�貍h
������/S<�5�i�({��N���E~��a�j&Y��T2fW-�����$�:=ܨާ�\{��
Y�����m��Lv4k ��[���#=]0T��s�'Q�
6���SnX���T��|Jl�iZߨ�Pd��dI(YQ{졣��@���^u�Ȩ��De7
0��~&��d�
�js�f3�)�p��&�N����E�S�2���JѤ���{gX!z�Q�m���lٹ�%>wc�MIwTSͶ�j�w]�i֨�(�A~�M��`
�ل0���7+�Z�KGw�^��=ê�C�g���zi�PPC2������	h���T�c�9�aQ��/��Lv��j�9�S�ܦ�f�L+g���k4!��l���~&K��esJ�S4���Չ���JS��E�J��`B~�Azzz�E7���f�X�w��P'�=���t�u� r���R��4m0+���p�?��-d��#��6�ǼQ��a}i,H��3#x4�t��hR�sY��6-U�t�j��ƙwENVT�/����܅���P�˲��;k'�����ҭ�3��N �(~Dx B/{��(W43�_%�׻+ h]M�߉DS9 ���|��ڱu]�,���߯�m��o5�'��0E���u���EeE<k��ZT��o0��L?�y�V�J�7�N]�^�E��	?��/]r��3)���0�彴�>�x|K�c{���d4^�\��ˣi���&XJlW*���q<�x��й0{vnDE��X��O�����;��,T�{��b��:�\����(Hc�չ�o�vG�t5��9�bB��2������/�v֤DM)M��8Ff:D[}���#�CQ��S�C����}�|[K���Y�v�d�g�l�ӵ[_�oQ+�"�_��|l�G&y�5&�ej�N�:G�^���w��^y�>�C3?.�(	6���Y��b��%���@�{gi���GHϴ C���[��I�3�l��җE'x���D�[�D����)�QFq|m���gSDRIAg�[DW�fI�8+Q2�3�D{�ͅ;nlӽ�NU�F%{���!��"�zEB;��߯5X,{�����ϐ^���'g����[��+o����1�&}v��Ԟy���у�6D�����n+� Js���(N�G��~��Ŷ�O]�K�q���6~~���l+�U����#�}�(s�1�J���V��a�҆�����"�V��g/�py�I[X\:���q��_]��[U�Z�R������b}�B�=�Xev׏ ���Y��p�#Uщ,(��ߖ�h�Q�Ff'	_K�uv ��ST�Sk.��'��59�d��d���~}� ��i�̀��e��kg#��r��F�9���g�}�|`�l���l+bzy
�+���mW	Q)NZx��D�D%��9D5ȼ=(�^�*�Qu����u�NVY����m:����so�����m���_.u	�>��ܝ�^�Ѳ��U���&�ON�RJ���L<̭W����\slX  ztں��(Ls`���є�R-1H�,K2��s��@���/(��0���fbm͑�k���sE5��/�֗�ntBZN�6���];&�jh��X����\�p�� F ����M4�$��{kIq�Dj�4=d4�|[2�&�|���M��û�_8��޷UJF܎�r���24��i+(^�e�,.�0���ٹ�p�� �σ���n0W'�BqE��9�OQ	%�����ͯ�-���B�[�#�ϗ�d�ѯ��0���]��Y�B�g>\o�|Vo;�壘�z�w�ϑ��.Ȓ`ae��q4<��7õ� ��f�I ��Ge%�=I��$���:}�����dv~�g�Q($����ol��7fƫҲ��l�$��]G���f���
�/���`��n���r�y�zdBP�)/v�͏��>xSl�y��
���rj;�@������S��<.{	���2����t]����ڕ��Q`��sAo�̀
rf�pZS�k`�g#��H�Ui{�!�XqE�m7����Γ�K	�� o5ޣ$�/���	�Ы7�6�f�8�mգ ��*ͲM?BL�K~����5��%޼�����MJңّǔW�s�l�أ>�T])�+����3��o���<|;�����i�߂v�dvi���z��~ׯ"�J�=�5U�P�XG'f:`��K�顛���U?�BÈ��ߔ����a!x�]� �M7�&�4w���S�>����
�xy����R�꽋w��3�z�2 �ƞ��og�SI���|O�A2x�D�ُ�=H����������������t**���Ҍ��K��ɣ$���	A�WR���y1�*Ɂ��L�+h��L<��A�G���Y�MD�}�k�&a�/��V�>��i�b9��i�r6��4�؈��ԥ��2���� ��:?A�K��g��'�{ �==X�qr�/���V��Bj�,Q�Ѷ�Wof�y@+���'?��A���`9����ǘh�^6H���·�|�������$$�E��iм���J�s�����+�ك4�tE�՟��^�(���ۆ�G�w��[���Axt��5�;mg���XO�Z�����Rs�6�F�����&�(�f�2�����>&�dg��l��6��o��o4���= �:-3sp�	�n���X{�uJ�Ol���^!�~��}pA�,䧙t�����H;��k��Դ M�R\�j�����i�=T���Zɕ�)��&SH�ݤ�>m�W��~F�Y�W�vik攕��=����D��?wqT?�@�I� ��ŁF��8����K�3%�r�]K�-���|lN��h
O�,��vd�x�
3���!����%}8a�#����3c��c�]��6�; ���Z�?~���Rv�S=�e6��>}�f:��}����24�/��AȢ������'�$9:�t���Dgm������@_�P٦O܊]t��Y�:�Е��~��Uҧ+䈿SiCT{&jѥ��\��(3��H���ʓ�BȞpPz-�A�ުY޼ݤ��n�qe�Ėm�~0�{��*���sl���hq��2/��c��9���a#��دE]����df6�+p?%�l(K�n��9ҞKLy�ɴ�R�׎I��əI��jy]u�,�py�(o,]�)2�l���:Qp��*I��5 |5q���6�]Ia��t��@���98l��o-���p�Ќ8T�_q�#�rS��Pb?���(�A���w12b�m�}���OX�QYI���M�$�_fg��^5�-�gI��z�ʾ�ԡ#�.�Wo�.q" T�����k^u�ZƄ �����C�B����2�[~�_t��A�q�g�	�3�"����~0�{]|ZWW��G�Hp��:���̟R�O:����P@�sgqOx��*�s^�
��ˋ3��s%��)���4'�mo�`�#5��?7�i�H,���䝥y����Vl�Wp��>�����c��b�w�R�a��yHIY+k`���r���g*������ ��i ����pE+��Z�)X;�zd(u:�d6A��ʌ�P#�<?�#��N���>�'5����fEp-#H�]�n��V�^��D0�v�6e��Sg�����ILǱ���1l���zKk1S�U�r��ɃJ�:���&�4O�Ϸ��ɐ8p�&S���::����޽cW���KV�q���x Sc��]^y��}Tzn�)���0��8�������9��l�0f.�US[�y�RKg�Ǔ���>�x�z֊�U�t8i+X��E&ji�3&����.��a�$̠(��X�eg{h�.����N|bǐ	v�)`,w�.��f�[�����hd��|�m�����<b�}��2}9A&{�V��HF��> ��`�7V�ז��*i��p���^lED�눝x�_S�'����(/6R�Z{���uG����嚞~~�'A6+kG��Z4x�[��Z�Y�C�I8�<),�� �@������o�����7��{>ߧR�c�,�]9xIɖ�)�`r?����Z:���re�m��BW�K63v�"��$��i�MD�
�ԿLr�nɯ��P����j=v���:��@$x��:�FS!c��j��#vt����e��*��!SX��*��UŊOܥ�?U.v�dz�'��z�d�E8.�ƅ�>�AH�ְ�G�w���-�h)�OJ�Q�E�>fӶ�������Z��j _"�]�Z�Fs�*w�����{=����-w�1�#�KHG]��ߣ4����v
�/H����
�"�UG=D�B��6�3�p��쐶*�;�!�y���$b]ֆ3��^�]2�:֔� �	E�F=2#��4{4y�aᶋ�r냮`p
��
&d��*C���a�����ٯ:��r�&92%9���	2���	����x����_�B��C^6����/��P������?���l�M8��dvgCX$�*�r^���,P��G=�1
�s�ˢ9���w.���(o�Z�HrF93�D58�����q9�˫�ݫ��*�_��������=xBzPg�t�9~.>��T�uʄQ��jn��5��&�њ��U���4P6Q_Y.�m���C���\�<[-j��^��*{�c��Θ�h#$�qK�sY��-?�<MZk1��Q���߼[�D/q�k��YӀC���\��$�"3�B��܍��+:�?�������0eJ��u�Vfo��T�)L*�]��M�5�sǐ����lvW��W����E�y�M"��榘��ͮIh|�	e8FD�����ueW��=����|��� w#��@�O����.��z~�����ҳ����mFG��E��Iq�n;��Y�~�o_��W\�X�O'.��b��E��8��=�G֑��n�2^nLX��5�<-U<��J��	��&��oeN�ݥ�9x��ܣTlb}{�1Rh��j����l���B75M���ވ��ӏ����Ӂ.��>��l�]<i�����9"��ͣi??��">���_�(����9����h����7�POE�;eڳ�����GG�@T�$|W`�~D�d�dA��6��=��)P�CF��;���>l��ˁ'���1O��HSn�yz�:��Xw��L3��W��5����T~��PmB��*L$���LĖ
��/� 7)�Z(�5��j0O0�i!�9d��5rK���*�|=��;�.Xn������U��6G��>�-�QlY�vg?_{�k zy@^���{�;P�s�m����ϓ�vd]����t�\[/Oǲ-`��u�,�	��~��k�1N�v}ann^Y\����sA4{�燐G�-"�hVz��k��5���_B�I˯2v�F���h���+y�epe�����z'�aJ�=֮�,@�r-���K�F/ V�B�����N��ofEe��x?>��n�^�x��	:}��﹘���(��[����W��:|oz���mh��V��Ǔ����� E:�����C@��1�3��?���[�
��
_���3�d�{�_��Ť|���8��aJ�92�Q�ʊ晃�A�F��%	��E��ϫm�^�6V��";�Ya��atl��v�*�{]����J�z������x�.�c�p��,����R�)�!���{��::ȵ���=����B=ͭo�%�<�S���� 7�M�8f[��A��N��ۯ� ��Yd$�{-�^��J��x���V�mJ�� u�7��L��TI�0l��s|��-|�g�y���Ư"L�j��P�E5����b��T��zTH5���\N�hR��Z��i���� u)��SkD��oFN��_i���*��i���G���	1��Mv��mBmd�<n2h��o�g:���$dG�2� �W?p�O�=��i7��/��+� �go�:�l����:f誌e/��`�6L�>G�qt��K��v����ϽI��r..tz,/�P���~�.E ��0��)���] 1~$�y�{g����hH�a.�ZC�D�T#	կ�TKQ�T��:f�o]�A�}0����!:��1��b`d��0�d��څ���0��z�W>K{d/�V'^Uo�@��-'��.m��W���a�3J���[.�h�$g�7�h#��.c}���M��)P'�$	��c��~��z�%Npg�-��Uv9�}�ـ�\<����Y�^�0ω��s��0�2���*�_�6�gJ����aH���q�C�G���.�E6;f���A�N�=�v9�%�sl�}~>�����D՜�����~�\LN�ǁ1�v\YP]�^`�C!��t~�>&sMq��׌c#{�^�[m���꧑:�;�
�,5��:���M3y1f�|g:�<�*5e���8g�9wH[S��#9�~�nG�Ѐ��RC�n<7_�w�����F���*�E�{���
�{a9���$&�^:��ظ�����9��H��z��>�Q[*ƙAr9g���o�ZDĸq�L�cT��n"c|0��װV��&.�~�u�A���1#���R/���L0_%�^P����dA`$�ݫ�� ېՏ��6��;d�sq~�~)I�R��6��F������f���ĮO����m�MZ#"� ר��%\wV�f�x����A�W���Ɍ��/e��-鹿�5�k�1J�o���C��G���o��a1x��^�o���J�$=_a�+,i�X�NGn��4L��{��&��DZ��Ҙ�0��/??���>�)��q~��/��k	5�!b&�d#�$_��C"â�w��v{�=�^�J'��{<�}nz��F'�Ι�m`�G&5� �=���+D�5��AM��R$)}��~���Ϣ�nx��J��ڟ��m#�	\Wy�pݱ�8`�@�����q ւ`''�{�o�Ä��Բe�}||��ȹ��j�\�/�����c�wT���3rbu$OɃ>���z�N岈�Xm��X�!�ov#�!�s��Zn�'��$)׉9s�'ջ)ՙ���^q��U�T�F����ˡ�$�]�5lT�8�����:_7��4�؞ �Z͊W3,�D�BȂ�ވ'v	�MM]<G��۝�6�X6A=ޕG�X��P�7̟�!x�wq����){F��il����������:���5���t�'���o���j�ކ�w-��-P	���ٟ��. �隘�(
��T���qT��?\���6��c�F-�t���>�c/II&*Gٺ�"wpP��m�k�USB���~�3΄�T�۠8a��!��2�_Gӛ�č��ݽ�
@��e�D"�m���q��}W|�ݎ�*���E����\q�PL�w���.qm,	�t��m�T�ۦG����w����s����	A�r�$�S�,��{j����2�c?ݫ<xl#��|���c-�L�^�{��.-M��e�Q���k�Io�s�������/.)-�(į����=xnꃷ7r� ����o�P������6��=4$����Ll}�9�U���%F�U�����Zֶy�1l����z�篛t�~:����)s�1-͢��8XTX�cBEEe�=���5x�~-F��T�h�ԡ����5
�m�g:ٜ��x�?�?3<Q������R�`V����s�w�R�� u�}�  I����|���ڤO�6���=o��\��P�P����8RCa���28��W ���)[��g�v�1;2R|f�h�ݓ�+#�]GT���\Nr�%.ڿ�OBʡ7���qIp2( �}���>��)'��sG�7�Y�ꖇ��g���~h)�~ŧ�	A`ߋ:�@n^����]��bMz���h�%6�b"�'xG���g��;KR��_��J��g��IW _d�n�z'������;�"� ��
���I�tA�|�ڶ1�e�/tF��Lg[T"J4F�4w��գ��`$���-��~�<��|P=)��yw�H�Hɢ��	K�y<�,K��y,fN��.��Yk�E Nm�,����>�����Ãa���r[�>?A��T��4�1c��	��z��~˞�ϵ1���챷9<�ߺ5���2w�e�^�ͬ�������o;�0;��n��\��
��S88+)I��'-���L�5�AKLL�iC"+�ȠcH����N��W�z�R�kT4˷���6��Es�V5jj�����_��W���4 �en����WZ��������{0-m���D�2g죕��h '��}�S��1�t$��?L�J�����h��"�/�f��XTg�»�������x ��t�ǝ�9^4k=*L��@�����ym�
<<��D��դ��/X���!��Igʩ�>�r~,}����]�-�Iܘ𵟹ߓ �롬z���U?B�5��oz@��G�*3��_?(I@��-�X���#9����īW+=Q2��zx���Z�~�q\Q'E8W�#+��R�N�6:|�~>բ�DT���Nd�u|l����@���3[��i6��Ͱ#�JD�)�|�Cro�� ������X�4Z�)��̼컓�Y�g�pq��I��K�㼆�HF~���N]髬`%���1q�)�8�-���r���Ztm����iq�9��w角��xx��)��&V�9�X��&Cj�����\���R4m�6�77<�h��78��dL)�Ĥj���`p��_�6v�~�âg�������_����.�fO����&�(�U���_af2�j��E�D�`9�ͫ��p*kM��G]��ks��E@�*/_?�5>�r�����u�\�����tzc�P#3�ccb��b�t�5`�9fnGI.�-����L��!���{�^8ފɟ�ty�����*MC�ex��
���a�6��?�:X�pۆ����U��?���T�s�~~�t�X����"
�Z޳?��T�`'x]	Q�㳳���.�_�?��IMֽ���hX23,Wg����a�<�=�����^7?��L��ݔ�1M�����GY}�~Ҷョ�.(	�eV dO�4?3'�c���嵴�HGx������vj�Ȳ�^�&�m���a?�V��ű��w[��}���� Ө��1������_�}w�J^��/�S���=���3�x�,Z������.���9i
��ΐp�m���KT��s��nH�ow�W�W��V�o.Ƙ�WR��I��0��P���k1����X��
�� _��i)������^���G �G%Jnw4yl��B8�BSM�<S]����1��/k8B��3�<8tO���^�l6�S��ړ�����X�3��B��L������_O�uԏĲ˄��k���k�EDEQ��(��\��`M�@�����=�CBW|د_��<�S�������������<6�_�x[0p�,�h�`����:e��������vs�꛰�_����Vʋ�#����kfܛ���\��;xv`����tjg~��d��������z��t�i��1:�2޲
���==��DAW7=(I��om���C��r��؞x��ś�����KY���gF�������Pd��+DV��*���S�j��Ym#�H�9�-}D�u��1uќ����D������U�[���%��A�I���<�y`�p�4c�!��$�V5A�>�췻�O�`���G7$i��.�MFٲ�0�L0�mwf�t1�+�g"6}��>���O�U$��$��ׁ��;�����KO~�����g϶�B�f)*���}�!�����x�M��&\�S�n\���zy_,w�I����,����M�g���W��Է��fe��ަ��v�����Ļ7����e?I]Bj��Fm}��Em=G��ؽ{w� b��a-q
�fdq1����ƋkzQ�sc��d���4L[��W��[Ee�������4�������Ֆ#�����x��n�-��	�^g1��A�P��c�+����G�_#�>�=�2��y���g���P������5�4�=��}�c�0��
(4��h�^��4�d�f2 Ҭa%˯��R/7MRI�{�z�Y��[�5�;�^++���y������ĳ��?7^�'�2��v�"�7�fpZ����!�����Ӥ�����c�8t;�<�{���B�;v��hpA�� ����U�,ޟ`C�`yg��J(#6�_��E��XQ�u%��]�zY����TV�z��W.�)+�K����+� ���p����&�`�k��/Qb�y��.d����R>~�V�jl������_&��Q���lL��Q�,��]o�Tf��O�����e�rn�l�Rb���Qm�� 1�(J@��%ҳ�ETBa#��ٖ����1�>�'de��o�����?K!���)p#�3��ݖ��;]�<n2��l�hB4���],��ڙD����N��.x)���� T�6�wA4IJ�?U�}�;����}�$�(��.�_ޏ�n�|���� �u�n^�+�w^x��������z]��;��\x!|�Q��Z�=c�J���+vnǴ��#�m/9y���A]�~�pr�,,ڔՏ�A�����B�ɠ	ߜ�ރ�^\;91�� �m�!�ZIm?O�t(Xu��b����l�ɟ
�<*���Aj���� 3��9�5�7^p���״up숥�ޮ̤nGk��ͬC�7��� 0��9��`��������B�B�-v[*���EB��<���GL�'�ٮ���h�%����C*��	:��#�;��ַ��L��欈'����6�J�]<�M�6-�立�>\�5~j{L�ymA���ٹ~��F�p��=��1r�"�v����P]�l�cb��ȁU.--e&�H_���(�M��� {����T��ඎIf�!p� H8��
������<z{���|%���n:7ɻ��^� �n0�XjT?�ba��m8uX��/l�aO&���$�H�i�9������_Y-Z�@Ѹ����:��+����*����)�W� ;�zh�/� �Y���%�´��Z��p�ɉ}�S���Nkd��2���)d/P���8���E��2�&����Ӊ���bX�v���qN{�$�I��l��K�ɿ���n+�$i���&�%�!����*��$:4��$�I�Qԩ'�50z�����Wa;�i���5�o�K՘ħ��̆�Ɩ՘��~1u:�X��N�4�H1�{���!�s]�Rݍ�Ħ������CE@���j�c�w�]��U�F�]��5mc20263���4WD���z���N�AD�'Ԟh�>x��Jj��o9e@��NP����\���譶<���nE�ިc\��"��F��������aYBk=͠H|%8�!n��_�<�Q��+~�L.��j�t�i��U��@R7,ǪP�[�;���K�P�U�������@xێ�̔:3��@ޛS��ٜ����^ĎF,���;.-cc_cݜ����88-<o�Vu���utP��Z��R�$���e�AoFmA�>�r"/?s���9����E�i����o�#/S��?���2�Q΀��U��ǻ0a�� �t���MNB�QG��"xnͰIې�{�K���4�FU�^48/r6(Ғ�H����3��S߲��� ��&7�cvn|���Ƀ�'`e�F!C,M��e>̤&F
Y˯�1y� �f?q>�f"�3����Υ�ݽ)1����-Y��ęq�|�L�|�y�vA���G�"�]���A41
�Nt�����Ck�k���sӨF�����/"��B){���MQ�O�y�֯����v�H!��Kq�c~�� ;��|/ |�X�&,?�$��U�x����֝ ��v�*n��4�Z�,i�G^8�,I�Ƃ��Y��)�Nf_�RD�j#�bRxC�6�ac��,I�;3X��{�3,��ṝ�Q8���s2�5ed�2�f
8c}8گk?��£R���h�K��-��=~�l���(R�G>�2��2���dGl��[� a�2 ���̫��f 3%]~+ÖQ})��𫜼�=74��o�ͭ��z�}j�ؿd�W���E���o@D�͗C6w�]���� �N<S=�n��h�[�-���%��,~D�i���U	]Q����l"r}@<�wCq�3�Q�6�`Fmg"�ɰ�g��_Z(}p��ew�o J������v0������zGf�W���cptiii�x21r 0��e�m9�ԒbC��p5��9���g��[�S�n�	1����}�/���౳�!�F�[t�FGG^������ħTK�8c�p�P�<2ٌ��f4��nu��i�#�=����f�,����F׵�fJ��6��cx�
^d�zy ��Wo�a�鹁�l�Kl֡��?h�S�M�����#'�~@UW����Ձ�R����{���6�d�5&��[i�O>h%BR�V�	xN��@�!4&/ϩ�M��xB����kB�����t��yZ�_6$t�MtJt�kNN�D%�e\GO��w�ɯ�q���k��S�#h���N�V�-�T���>q��d��!F&�K����|PQ�Ƒ�B�;��A���-A:RWp{��Ƅ��nG��޼"��q�9�ov0W��-��u�"G)ݱ�֦��Q�J����(�D��S��}��]�`�땴�P��3S�4�l�P��s���~O����L|���0�cnh�x�?�݋�uZ;}�+�|����Z
����E������(���[r�[��L�M[�q�{��l�6W���߃8��rJf��y%B�B�����R18t����@����=K�� ]W��p�ym#q�+��[/ �6��s��1_s]EG�a�#f�~�JR}�m/�i�~)[�q���"�>:l`>��o�W�]�`��4�V|X�vl�jl�#�X|��¦W1�i�VbL�N���O9Y����ȱ�B�/I���m�����q_�c(g:z��p���abDg����&��'��bS�{M�H?�E�l�tm�p����p��j�,"~��i�I6��D���fk^�4a�l��U3{4]��턭:�;ٓ�����S�MZ���$����ʶ������C�u�n3�����G-�lAhH
O�/��ו�.L�^ ����D�>�iC��x�� �.oZ	:Ș���+������ǅ�~(�ֲ����N�tP���.0�M�KE���gZ�P@;F�S��x�i?��.N�cĦmH8-5����{9����:��Պ��9h�����?O�M�uk��V9�����'����s\eL���@��ޱ��>����E+��lB����A�+���HW�?-pc�x�${~ �c-%��aU\��
?6��XM��C5g&´~|-�[D�
Z��z-d9g���xJ���iA�>D�dvπ�� O)猶@�%��~��U�iO���B�N��zU��Y���VN����>����������P7���q��Fח(�D��#�`�{sj�ߏ �<fj��&�*����MK%�H���N߻�~���JZ�B
��o�2���z:�{�L@��cr�D�g��	~P঑��f�k�RՎR6������dzA�~%�@��ޱ7�%F��Y_�����2W_2�Ѡ���Ѹ�
c�Q������О�2G����T��m�$�V�K�'bΫW��<�>�����utPQ�%��Vl\}r��q;2���AW�,:�A�"[���_����q}����=�WHJ�\�7E|?�Y��9cs��?5M�1
�q�@\`��s���{1�R��xʥ������!t�o�,&��2��䏜���:j��=��j�SE�	}6_�_�#sL�K�ۥeexl���f&�[�sN;_��M��5�'�DZvtt�Sǣ\��~�?��q;E����� �Xh�8&S���[��9J�9K�
��&�L�U��]m �8���}E��ؼ��6�"���\�5޲��kː�Ǿ��ߌ�=1w��s~]�G��lV�,m���8�<�J}#DJcBμY��uuХc����v�s?�qa���������4����g���o�I����A����[�d�)Y��*��⾬f&������1
jTݞQ���yׅA�Bk�'�<��g�v��r�{���/nJ�M[r��ta�="F�'��c8X�f�y7l��8�)U�P��Jm�
��L�\)��Q~��,~��y��^��e�ڿE�kP�9&X+����� �6�q/g2H,�V�i��\��)}�?$��yls6�sm�g[�o^
#V�W��j�lJ?�����������w)��1E���\o��[�?e/�����H�J$^x�Y�6φ&7=76.%�V�^l|�u���u�L���WR$=X���u�4�7��*�M~6���X��d��s9՜z�p5r 28��p,uvr7��	�t�%����x5bL�!�N��	!tM�~�_�-��/�j�.D���J�Өש���=��k��֜ت�Z���wű�Q
�M�Y���a��⛝J�F"�k�3��fA=yZvOc1�qa�A���Gl(�w�7e9s�ٍt��r���Xx�W�[f��k+z��L�i��?�.,�s��lM�g҂����"5�0���K�P��>=�l�����큽 �u�tP��d�w�c�wVT������k㼫x���B+D��E�g!���p�G����U�>0$y�>�F"sa����V�/,�K�k���ԣ3���k�EWq_�Gƥ��o~��?�p!��C�M>�͇بurtg��Hs�;)����kVƙ��s��u#���[ p,8��y���$�=/�!��l{כ6����C+��3�Ǽ4�?��S��[�����n!����[�pGQK��SH&(�I�D�
�%��=g�h#�:q3��Sr�+2լg�i���w�\���,q;6g�1J�*n3KEs�h���捬�*��1Q����~"��R�M#� �	��N����Fo�%2;�J��Z6R/����0���w�E��y�-����R���mI���a*Úȕ	CQ���Oz� �,
r������4�_K�]#� ����= ^�=EE��`�'NbK��E��̕�?���)d��/N��0�����G���U��-G�cm�.N�Q̽��ӈTh��MA) .���r:���HC7�fTf}�\�;%�R�����$�i� Ut�.�Uwi�Y)j�}��&�-�io��� 'a=�^����	f���/Mq�qhj�D:+���F k�����F�J�� Gv��.)�b��P[��*�bF�\4K�Ir�ۊ����Ty���@W$�<�z�w�@�r���(���l�w�JY:�ou�G~�4�n]�5"��e䣘vfmC3�{��� ���ҹi���B:6e� ��8*Z9�����n����Aۻ!W��`��c;;.`u��{�m,�����m+���1��(q5m��#]rJ�͛C#6�O���LObC&�����ĕ�x<��"�>�Q����/q�he-l�Ax
M����:�(YDn�/-�܌��7��F�պ�@t�n�׮�
|;��;�M�\�pZT�-�%�Y��h(KS��:� '^��.ϟ��8|*��8��c�� �1[¨��zL�t_X�� ���k��tMh��������\��v-[��U�RXB"�P}ɣ���Ә7��b����P%�*�4��K{ё0��u�py�f�A�c��C_��W:*�BB 7?�ي��
����Y��<��Kd��ed�q�aMye�&(��=������D�Û�$X����afxy�5��+h��JX�����5��������[��[Me^,�S��G۟� �-����g�]x��� 5�哛t�n�l�~8��>�ޖD�w $��^[�ls�_ C��@�kD.FF�2<H[��.$�'ꐁbZG�zsՊ��UE31g
�ӗH*��#o�D`=O"��-���m�y��6�u�@"əӵV�6$ ^�^y���\���ϩ�p��܎�um*�q��aW��ٯ��f/����ѹ�����y�Q"�-8o`��E5��ww6��W�{�������{&�m��7,I�{���%�?�B�X��#Ci�����2�]��!�G����Y�X�����/#��h8���?�h*ؐKCn=61���\.���@����"/�Bs�T��+�z���I�������t%7�fp����ku�^��>N���ƿ�_ɕQ�]\a�j�s`{�43�,���E�k�כ�Z{d�����|n���b|��蓥�d�R��oXkQ`d�3$���3J`�$��k��e����r���[Ʌ����[[[��u�	dE��>{��z[VV6�$����[���2 ��y���J�p�Z?������C斛�����8gh��Z���b]������	"Cވ�bhhx�_0b�Py����A�X!humە~�=����Q�Z�����ɦ���l>��^��������KL�^���K���L9�9�w�n���꺏����-}����ѯȢ�Wpq�hi?>]�t7V�bQ��442z���m��ڊ���P��"�XƮ�s�m�'ػ�ֱI�#�*��U'�: �Me����g�;��	yh�R̠���q�ʤ4yw��_e���:�����e�+�j�~�\��Ow�j�S��N���^:ck�3���~~~�k��Me]��O�?_QTT�TD�*�RS�Y� X�S��u�-*b+��u���3,+`%�W^_���sb��؉%J���#��t����o�}2��R���d=�%��H�9fM���D}w ����Re��2"d˵�̌Kdĵ�][�L"{�*��J.���u�l������������u���|>�9�u^��>Z��x��p�����b�q1���yٗd�q��`����tg�Yh�����SӮ�Om�ƳU����/���>"��|6�CI� l5�{�[��o�~a���%!W�:Ǐi7.��Ds���N4q�4���)�u�#<�������.�
P	R����2e��M�V���!�o�t�r60<�K�mc��<������"�0S��u�8��d���@�?��K��G?D�s	��g��&�Ӡn�_GME��l�1��Z����Pn���H���d5�)�a>Z�W�ezk��|�{��c�I/���
�-�C�7���B��k� 67\����A#�Ʒ ��ǭ�B�@���.��w�� ��aN1/�F�f|��y���v�.��]����u��3���V�՛��O�}�]��֦�lծ�lJ*�
��4* 08�^cN�R/���]>�yo���7�v��2=�M���o���C�\��=��,�{�	��wN�@CL�uDP����X�@��v�~-%�L3g�`�J�wo�}��r��ST[{�tC- ��W�Nl�sB��S�$�v�-���m[U���꾹����K���<�~�?����bߋ�G����Sa}= |��Jj��w�_]�{G(����	����- �fa1�ز��+8���T�w��oS�7*�L�c��=�k]Z�B�M���p�$Iڐ[�z�Mf�1�tt%�����'j�rΉI�r��o�S���3�ș�?3��rb�K�\\�~����P4)�[��� V�B����\���9#|yb��H��q��!��Cp�yS�!��N���Ԋ�=Z��&���ږ�}����-obB���	�`�g��p��ӧOW��.��gʭ�I)4J�n���h��Z���nD�*���a�2���Խ
$�(c� ����'~�i���8�2$��(Do���������Ǣ�{M�r�� t�����I"��,E�/�g'�_���>�{q���B�ʶ�,���"=�'�u�ݬ-H�֋*Cjb�L҈�c_ɡ�&,r��`M�"^��9�7����}R��K�r�;�$F�:�je�G��|8_i����am�
� M7�4������{�p;M��-����FK�#�m~h���l����ۻ"��o�{��<���Ш�n�q��������nJ�-G�]��$���ҡ0ᬷ��3jb�Yl1��NO��r#��.[�:����5?�U.�����\�b�W�/�?������e&����VQm�bZ��W��Lbg��&V-՛�/ �[{�>��=�H�j��4Ͻ[0�/���v�[��A�7���O��i��gF���}w���	
\��RY:�� &�jϴ��_�Ďu��Mc�G���M�^���{<�/�����F�P·�	�LK�P�������~�%��G�%��s���[�?~(�j�e�v��kZ���s���=�y���E��=_z1���봺f�	��|s�?�w��K��[qr�'��ZKi����
�X�7A+�(���e[1�R��'�W�����U�6(ն�g/��]$ҢU�L/��!��q<�7���}#R�s����7�O}!Nl/�\ha*��Щ�{���i��l/�/�.��y�`LFi�U�ݾ�Q�K�����Ĺ��T������he�7r�O�'|�UM���>J��o$�u%�E� ��%��rGe����آ�a5��:���-qWB�!ڟ��)���{E���R����s�#�����J�j����Z���Ø�Z&����2(RR҅݀����m�e��(),����d� �T�~�Ck��d�_���ߟK���~���b��E2��h@���;�ke�S�)����zG+�إ�ܼ��E�u�r��jd��:Y�@ڍ=�5��.��ԣkI3>rT�Q��b��u�o�%)��gM,Lo�Jɏ_��4�������S�?Vp��_�@��R���f�r ��o�'�B�O* p��qÎd��+S���ʻ����GI�y�����M�a��Q���^`~��Ȑ������?��Kxd��QZezz��y��P��U�Ѻ�+ؚ��~zM\�b��r���k	��{'=J���h=����9�n=����ˑ��4E���--W�������2>�N�K�t�9ʝ݁�/3i"��q�< ��7&�=)��k+?cX��| |�-N��М>ӷ�E��?�� ��lV�{�,��m�wѴ^�dt�}�M��'�bf�Na��,e���nQ%� K��\��i�8����@�]����Ё����@��zB���cQ7z<S9�����YT[�]JAR����]�/&�w(o��V�d8�|�J�K!B�	�~�D�L�T���j�jmjdW��`+*�X�Rdl�0׉>�pϊ�m:�2ǧ<�D�^�L�{/|�Vc'� ñt�8�09ڶ`(��PmK��naGk�ch�ѭ������J��ϫZ��Ն�]�wU`(���B�[xr]�/2����1\�zǸ��������������/��g�-�DD��r sTTT����ms��L,}�+n ��0��A	�+nz��Nhį��9ܛ��s�O]�^7�D/O�@\��7n�,?�
�I�9��i��ó�Q��]�TC3;�6��xL��P��W����?\d�h����K�5���S���{�p�%#C��) �����M�`���\;ui��(��Cb���ѳ6@ϳ��B�����ɟ�NTӈ��aE���Fz�@.d�NM�����M���6­"܉�4�*��t����T؅��V$%X���B��tt~��,�ciצu�:^%PJ�T�_<M���9����=��2��3r��BR{#L� � ��%Ӗn�a�Ǒ��f����?���G�C���$}h���j�U�� VO(U��� C�'eދ̥��-p�:�=3V�A⒝ݘ��}K�3���/��R�ݫt�哗,2m�i���N�#&����؃I�gD�WZC�=�s�+�%�c!��]K(����7Ef�}�����Ү����={'�e�����mf��
�EZ��0Vi�$i}9J�Q���u��F`�!�<��x���ə�<x��+�z|�fL�t���#.��r:�Ť�n\N_�RӦ�>c1�79�����޷�~^ ���Kn>�j���Go݈�#��5ߑ�'ofn(���+���܅Z%@W�k&0��Y��`��&2A�x.�j;e<)�XW���՝1�}�~�	�)��q��s��)f�.�u5��{�J��c�70��҈�3mk=y�s�hp ���G@��(��{{]p����vB#���$k�$�rM;���mbiQb�ʿ� �릆�OoXo�ִp�Y���\{s�k1� )-v�����������Tz��0��u���]D5@MI���$�Z_]M^�כv�I�4�V)� ��O��D?:��J5<�{��v�Lg�S��wf��T���/�+~-���B���M.�u�+K��$e�B�.�K��È}I�$E���c�h�n���s�}�m�7��1�-���Jw�Z�^gb���"%5z���^�:z�-���������/���H��;R�b~$qr�ml��\z�o��T�"�H]���e�����D��5b�K�`͹����˙�$a�|,���iOj,l<5&b���p�E2c�$%@ �� ��a_kI�5P�%'�}��h0�Y����]^+Ù3,�VF
�=]��j���{�S�t�/k>��A	����{��Ӑc:X!��ߺ;����J,��?=M�svr�˯s��rSC����@p9�GD'�u���蟼������c�2Ծ\>�\V6���ȣY�s���7����|N���3�릦��3z�>f�����~##��Y����8��H�a��8�y��"�GK��W�?�qm��9�M���Z�����l����>�~�,m��5xYy�40k7v�|�1���$?�ϟ?;��Ti5� ���ߟ���D���� ��x����WH# |�3P�h��74�L���O��+��w�2�m?���Z��(�Zļ�����X���1t����)\�5w�G�m�����)�3vsᦗ'?3��3����[���f��ֵ�P���;D��sD����=��L?�9�**Ĭ��9R7Q�곩3�������ڍ�R�!��ΘH@:����H�"+�e��܅�0�%R�F�����M�J
u��n')�=�~��D���kF���O��� X���A��F9�� R����<,��ג�_7����-���W�ϲ��.T�m�L
0u���|U���J�+s���8������̯�Y�)���L��6���|n�K��<q`J0�qm�`*?Mc-��А����,�]�5��#n:?�z�?d�a�ߣ'}�&�g?k{����x/�.:��[3�dK(rAݺ"�w��|!���s�����O��k�R��2 �Ս�$Ǹ�΅$�.�.y�I��_F����#�뒢���#�"44p!ǘ����-���M�� �wn ��C_-5���(����������:5;50!a��U췮A(�-7�L�
�_|����<��1�%�?�w��(9�"-z��j�%��4��J� k���o�J���bB�]1���rE�H�e��~0�q�[��?wuF�yn7.�g��p�0��9��s_���_-Z�k9e�9��>��|F���:��+�&�����`���Q=K�rYZv�����������Gf+>ʄE�.;�����a���3p��/�����;����
��A�G���� �T�)��&�
��Q� j�x)�+1R���trW��{�V��_kE�Ķ,�D���,-��*�������>��"RQ	�Θ��Ӗ�V�?3������._�<W-��)H��N���T~�+���Ke�x�L��,�gi�>�����5�}4���s4M��]��R��5ɐ���˵(����`�	�M���R��n�ġ�_=� �y#3��z���:�%tE-&R�R������KYw���w�
��|�8\t�8|j�T�Z��DD$�!?�Ϙ?7|���pčJ'�`%�5�G�W�uE�[H��&7%/�Ff(QM%�E�Ē�����ڮ55]X$�)o$�0"�0@'|��z��HQ�ScȪ>��LqeIh����/w��N%P�"7Ŵ#��}3�����)�un�WT {��]}��:>;/�p5lh�Z��o*ߩ ������˚��â�q)�Я��B}�6���DUW1Q��)x`uy���eU��S��vWN|)2������9�����N�e1�KӅ6������Q�ғk�i�7N��_@Y�H��1&>ʽ:���yp+�\Ӹ�嵕T�1��@�jQ8�����ʼkƬ�2�5]<`�?Z�&N�떼�`xI��NN�@�� ��I}ܴ��E�B��^eE|DD����%]��LKg���U����1n`�|�:��s���yc������`C��co{'ה�,ZYTC�Z"y�R�Ѩ(l��eqGp�c��B�k0Hr�����k��ǃ���=rbRG�v*P��VC�ٟf�'C���| �������t�ˮ���V	���K�O�O<\k&<���VT����;�vڡ�f��:�(��#�0:�I�{ y(��?���2��DvUd�ؕ�ǟ������+ۙ���v�*)F�Yj\��Q5!�A[����&��cPhOC��{w��5��yO����P���i�-���(qJaԹs�EW�u�p<��.du�t��.¯K��'U=��v�Y��r�{4�Rw/®K�����Q���}>�r��g�j�@i}�q������w���ӫ�Ƞ�K ƹ�]�==���_IK�;cO�sO_E�r��%��#_���,m�?��POM ���bޟUu��X#�DS�}C�H�h���u�6��?fD�,�i��*jzb�D�}߶jm||&�<�6���d�T���J�m�7硽�")Иx�U�
�-"�hr��~�!<�bb��8|[��
���/=�j�7��� �����&R:i�2��%���1d��k�G�z���!���m���:5�a9�bJZ���Ftv��,fEتB�N����f�{�W����/��9`ֿ���Qu�>�<lQџ)�ؐm���M(g:�G�$U�h[���gN.V�7� ���{{,�~� ���JoA�i}�$3�Ō߃�@zw�����g�i=׍��+E-NS��w6�wH`�{���ǻ�E�~��H�|@�l�CҦ���~��U8��-��M�@G?���;�JGN��)�T=�Q3�J�\��I��d�l��^�"����|bT5%>7FS�_t�=Mc\�����f���Z|��ASV�&7O]a��e��Y��Km�߼/]0a�G3!�W n����ܕ�-���������o̫�"B��|����Z�o9�>�Y��g��+�U��g��T��g��555�����Y��P�\?�c�cm��FV�c�Ӂ�Ӆ�o��c?j?��G���d��V�՜�(\Ma�`������rWT�8����lؑ��ԩDr�e�򸉶�I^.\�-95HvΞ�'飵���]9n�������@���q|�Fl�-[��F�ȼ:��������A��v�dO
ː$@�Wp���S��$���`a-��l�^���o���r�l"�/c����l\D��"���g�8���4M�����p�'���������Sӳ��^����ci����K��K���VgS�W	i#��4>��n�"����i���l�n~��-4W8Xu� 4!_%�9?3;����1V2f�ؽW��,���Oҙ�v9��(ڵa gr�)��:K��GR{�4��u��p)�z����-��/Dg�]��޽���E�5=zP�q�{�tjvv6��|�s���s����է�~���a&�����R��u����x����Za�I_���t�������%ǈ�:^y�o�mn�SK-�-�m9���(xtn�aĨ����l�N�޻ٌ�k��n(̪���
H���ΖC���z�x�?����*��N�X��A�cc鞡_��3��y)te^+�`X{=g0n�R���$�h��{�(�8��N/��o ^	5�&�[K�F�ݗL��N�e�����k!��5o��WV	�E_^�ŜNN��fLϺ=�������C�y=}���E~�$Լ�{�Cfj�;�.>
aO^��ȟݺ��z̰A�K����Үzn�@:�s�%�uc�a�\G�_"� �W?� �pm�`���hq^G�&:����+d���=?~m<��{)*-�8���#QQ��49W;���ʟ���������3}���Γ�ۘ;��&軃�$���
NvE����,�8!�@7�"��H�¬�ך�H�	=!U�������Y�))������j���Ŵ�Ba=��L�V�M�Q���*5Z���l>��Z�H<&Zn�����cƨ��t)K�_۬��O�Zba3����������vp���l"홞�4�x�g��d�����:���O⢚6�EO��a>$a�<���A���uU0�v�n.�G��FZ>�� �>�sh�w���>.��O���! �luS�>������Y�]��g٥;�u��!�7Yn��Hx��a�*�3w	������̸�^�@�GK�5Å�`3�tC6���=��s�ɽ,gFȏ�B���X�"��[�O�t����t{��Y$����t`�Ġ9Э��|��@f�7On�ή��`J��"#2��
��$Lj��y:��#���`�뤯�TC�86*զd^g�}TY�%�K�?(ɪr�]��)��TX^~?�PkYH����	�O�&}�x��$������u�,��~1�S��.�w���PW���LpWL�e��_z53:drů1ۻ��`85"lM�)x��f+���]��b|�Z|���� ��<�5����	�K�[4|_��z�D���V:Ֆn�ӟ�{���5Lт�5�:�N��葯��N��N	�:�<���#�'lz���<#��A���l|�"��k~�Ñ0���~�^���7k���Iq*�Z��͇�~��a�˶�@�Δ�_ i�7ɀ�Qۊö��&� ��!��)��������1�/��������%�w���&�hc�|����|�����HE��r?����펲ۜS��c���MY�^�;��1>u��-u\����&�U5������'>��c�F�ph��Y�Ȝ��VVσV�gRѿ��i��&G_/K9�*����5�'�@�r��p��нl��J�v:'bԞ!��G�����k��dm%
9d��I^��U��Ws�ߍ���/�5������a��#ZpՃ�RZ�j���N�G7%[���Kࡡ�5��z�tG�3��[fJ���y��'}C{C��LoC�1/}[���d\%%y�ؾ�RӁ֏��ʅ��Щ�cP=;�����7۷��4���n�քw���*Z��l��F_��<���}rs[�݂�y5`g�nH]c��(�!���dEv�i����O7vAϲL��[����55
Z�*N�	(:O�����lno��ոu����a(�.Bi+#I����ə�5wУ��K0Qf[�(!�R�o���=����2,�ך�P��qʦ��^s���ō�'y�Q���@fn�gy_��S�q	�YK��dp�H9')���P}@��z���4����ݱ2�=Y��j0�B�uU���6���(NNLdx��r@m �lW�X,{	�s�|��~4�;Y�HpA��/�@(?�1	]������Yю��9m�+�<�=�[@��Os�VW���{&�U�S����ħ���q��T�H��-՛x�����.�8fm��[�&����I^�diN'��nchTv�p�C�qJJ'h�;�+��b�4z&R�_9���X�Bɞ��8��2��(�៛����?
�c���Ľ��]���f�m�����z�/�1�`0�w+�����@��+dK5���T�*��7.B�<�=�98I����8Ҟ���
N�X37���D�$�H���_T#!�@њI��5�R�8Y�pv�1��m��Yd��d@��>�UbH�f���*��88��B~�ap��Γ�z���'h>)��[�$-����k�6؂o������P��GW�0"S�+�(�޿,S�*�5�kI&<�IƆ��i���yu�ڙgXɦ�c?�!��+_?��p�l��Ȅ��<�2�����:�z����.���:��$b]ᕚGq��J!#<O�'�[�*����m�}�fW�+���c�e����m��P"��&y��{Ph_�s��U��h��c9A�b�A,O�*
&2�eF�;Q��G�F�w����b��*#`&�Q���G+
4^{��g��e�x�oY9��;�
����!�{3�#r	RY��a�݀�Т�0dKzt#�C�˨]n�w��X����)�b���Я�eK~��"�r~�G���|�F�������|1���D�I��棈b)��l�����[�8o���J��l\�7
�(�$_'��r�����`����k���(�Ͷ������É��!�T��u���xk�6`]��Y3x���e=�Q`�� d������h�I�.'j�f�m�wS%w���\l5H6��A>�
.���,c���5�Tm�s�\k��|���<s�n�����݌�w2b�I �XhV7kk�1�+s�lb
��6!0<�����j��dW��z\�^��3��LIM��r �M���q�=^�7t�������<�#(���'�����tO�T�#d�~A�*w'Wgޣ�bO,������7�O$FR�'FM���7�����vٗtA����;�`c�����{��\���slM�x�HaU�J��H.	��صO�;�.u��TVŅ�<�7��_z7�����g%4C��R94�A��,��=||u����
�IM�}�8Z�!�S�7��N��Ǽ}�3���Z�驺"0k�<�:D���� u�:6i}�9�f1 �B��(T$/�9�J|��w�d�!q����/�^����|��j��.���싌�����61�)����k>���1�~g�qI�aY��j^k�kyX;��H������S�a��}�Z�S��yGI�$��	��Ə�*�W]�!��X�E�]��>�?Q�L��j����k'q�z�;���J(IMc��Jϖ������5��#Wn)�R<����.���[Y�`�k��9m�!O�M����������c�'S���FK�E��~:C���P5q����U-���@�JOG?<ņ���d6H������"_*9�B���֖�-��rjE5�,1�U�0���y�l��Ho��a�>4w����k+�_�����7�^�CM} -ֺq�o0桙c��س�.A�n� $�X�c�ȹ��ލ�"f�MQ��,���P��ߋ��!�Κ~^��B`��q�W�^E�+��N3qR7�u�sG�� �?r�h���!�ϟ(�X��<��w޸���1O��q�W�F��F���z�@��hu�Ϫ{0�N۹�����Ĕ0�Lv)uhǜ��t�����!�7�ШL���\�����AKQk�pp��*N�F(x�W�bg�P{�g!�A��6��O�`�д|�x��]�]I��2�2nkrt6�G�N��a����%ߝ�P��+��;�ƔG?4Uù�w��jj=_YE �j��Z�`�k4��#R���.c������)���(z����<�P�(4G�S@+?(����yˊg����9;#U��`����GD�� f����dNGӟ���r����8���=^��7������SXk
v@٨�����j�)@�f:�Ij�q�K�uN_LMBw
��p���0�������k�QXUEfڪ�)r" ���Ez����H�'�JR��Y�1�S���<��/�L���F���HU�{?$^�W)s�T��9��gCk�w[]���߭����y�.�=��I��w�W�.A���A�d�2�g�Kn�c����gvZ�q�㛗z����_k���_�"Ҡ�&�~+����B�=y�~��$�ntm��������]�k���.A�4�~��U
�C��e�Y�D��S�Lk�,�ԦZ��;bN^Rf뮩���e�a�T�Qov�U��N4�)1ޠ��H�ךgc�ڒ�1��Qn�$�zڒ��AO�>y��my���*��C�:�y4.@h��\�]gV�
��Z(:<�`�{f�14T\�0C �+�O���D��r S�����C=w+�VfH��N�Vӄ^
��f��M���vry^���vA?$g�� 6�Z�ľ�n�*��t�^��$eHJ��$���������/=]gL�v���g���Br�cD��p*@UW���O�p܉	� ʓ�������6�n��&B{U܋��/�![ҵ6'���>O|�t?��D^tH�A��ڝ���=�&��7��F�fg-���	Ո��N�G�컿GM6������f:f���&5���8M��.���|�F2t�{WR���څ Yhf1 �����-��8I�����l��X�ۘ���|�|GG�B4��x�����<yn26o�wO�y����i��y���=�
�μk0���~zk""I�W&w�x��.���Ծ%X�{\~����ì_�)���[�>ś���� li/����V���Q6�1X<�8R�1GX�N��F�9sGD�A����ɖ=9_՞��2R�����G��l+[�Kเ�x�#�Z�Ϳ���tt��ul�3��M� \��M+踧yc!�7�K��z��Gɼ����"��*y/�2`��S}�B)�k�-D��{HIK�T��pQ��H�J�L�Ç�Q��~3��ym�ll����r-����6�[S� ԩ}6����(��ǋ� X1P�L��;e���f���^�J�pE�mo3�3<}08/g q�a	�{F5LO}29�����P{+6�
�1������}��j�9"��!�-�[��% 3j���+|l�?�n:;B�<�3�zG�Շ�ښ��,���Q1`M H���\�9EN6�~�Da��i�>ab����5�����#�>���� ���r.>�@a�r&�I	mĹ!�i@A�O_�-g����J��0	�+��K���Yfa=\
�����͙��Z�a-\7���W���e�:����Ă��6U������Znz���ѻ�a�W��1��f�ޙ�>?��X���ٱ�<czi,��ˉlw��n�?�Hz����=j�k��-L	i���X;1u|-����%�o���F�3��$yGH��B�K���S�Vh"�l�qҷ�s���D ������}�bbb}u�4�9�0���F �r���R��Ȳ Y1���b����ȭ�V�����X�k�Gל��/��^$��/3(AX�pW]�v��yd%���C���T�LS(�#�(K�3v$t�*�i'��Z~x��X*h��oӺ�t����1v�B�ۓ�����_c[C�<}���dL���1Lq�B��t��`�}Ds6k�2�  r��-�t��D�S����yreJo""�NB��焊���:��&C���\�C����v	R��΃,uTO{�#�4h"���� �:���D!������i+�w~2�5\��\]��FEg%}�eɞ�V�lV���)���I�Ѥ�8o|���!�֨���ڿ��FD]�K����c8�l�5v�5Mz{��Z��B��t������O߇��m",R�]؁Q�Q�_^$r��g�Ѭ����
�oGl"����eN�N��ܷ�zo���"��ٟ��k#�=��LLLb濐�R���d2�o�(C�v
�S�
������[W�ƥѢ��%���PQ�4�g��<*:�0���M�{�'��|�5�H��w=a�Y+K�|��n y} �t�$G��q��+A�QA��ܯ�Z{M�9Xȕm�3�_
�uYm%�v�r�\1��6v�ޫ�̐z�6��5i��)���y��pt)����~6(]Sx廄Ѿ����4y�B���<|Ge��u���S��8\�֍���g}6�p+��s�^��I�lf �4�4|}���A�{��^�r!�\�9��`�?�=�Y�m�-�H���������0z_A�h;V�S�KDw_$HK���\�)��y�~�G��ߓū�q����
}tWE/��p�V7����D۱]F&wܧ�8?k�*���F���T���I`���)�"�47�-[?'�p\�!�[��T�Q+��-���x��#ɡ����_~y5��3�'3ɫ�l^GWִp�:1?�:X���:(ac]��k�qmgG�t�.Y��/�����&}C���,�S��=�^" ���?h��۽{��� �Į��lv�oAP�������M��8��������p�9Q�7������Wv�Sج��Ș
�����*���'.�&�gi�`5����5�U>�ʨ^b��6$Y����0t�f�6��.[P�c�<�c���6��.�����Q���0�yw[ﲼ ��r��%@�&����K���Sx�t �{ 6[��8\�C��>.��{����+��,�ħ5e�����8�����:�ǜu|�6h?��˧�z��u��J\0��Ƒ�.�[��zt�6F��W4U'x5omz�w����Y}Oye+�1��La�k����÷�V��3���>�F�1Ќe�������7�1��i}\�g��ǏC�o�q�EO��|�P[�j8'����B������Q�r].��9�r��0�op���'3ͮo���I��?�L&�	nI��}��ߺ�sd1w�70��r���K%c�������r��e-��,�ג\���9��e:؞����/�7�6k��k�Me��/��$�N\Fg��X}�cp���EB�o%FESx���a[%��:�`� ��-̪�3�{�2�y+�%x�NL�(���L�1@&o��Ҭ�=q!	���S��)�+����PLG�s�u�S��ON���؂*!�����U�/Zܺ��{b՛'et�9��_��YD�U2�Օ����k�����5�_߫*�2lm�������ͤp����}��	�m԰\�&Kc��,r̮�x��m�*iE�<���eÍ�/�#Z��@"� m��-���	ĩqY���Mo��J�h�c�{:�8�,�ܙ+P�� �bnחd_E���F�Gw]�m���LLkkk���'�/��|�N�]��T��/	۳*ΰ������� �mP��y��cz@: m�_��J볙 &�5e:}��pp��)��'�Mz3�L�LL�P�!)R��W��0s"u�󰀪f�xu0�l�Bsɱ�Q�yA$ߙ�UW�R^�3��ot�0���P��-OY��E��kC�z���|�Iz���*�%�5���k�ZW�� 
�Aj�GT�F^�����}�P�(hҗEZ� g�ؐg�����$�J�O�{����IDl4J�Z�t���(�����RM�=�3��O���Ѧ� 9ڙ�7��)D�{g#���5�B�� j`�p!��ZG�`Ӿ��8�k�n��k�H�~�DO}䂰|y��jkk���ޡBP�	6Ҏىz�*}Dh����ZYO�������ܽ��^�����ǳ�c����qD#w@w�NY{����D��Ё�?JZ�۰T`X*��a	]Oe�Xq  '����C�<�&���<�����d���U܊�M{������!��)�g����N��|��
<�\�u�����C�E<<��2%q�c�8��8��6 � g0�`��a�Vnȓ�j�GX0���)��N������{vY�8ΓE�B���Aq�A�IF=/��r'�-�%~��f�����9���W���L2j
�1D�7T�Z����'{�K���4��J^l|<?6�Zg�Q�3d�xJt9�agu|5"�o��(����K~_�d��f���ss�O�(2�'m�3c��!�������s�]��̷Gd⧰��n���m������3�xA��Hw|����L��y��[��T�d���UW���D¾�>����P�.ЯEݴ?�Eտ�3Hn`��-�[�f=_2����@H���i� ��(_(4�nЉӸf���?�6b�"��k%�?jc�r���� 0I�~ u7'CJ ���Ev̋K��l���#���ͼ��>Z_RSvNa���_���FT�W��<k8�
a��~���([���6��yp)��|
zf:����
d�Ϸ��U�Г����'Wt��Nkm��͋�F˰l�&��8OX����?ܳ�Su��A!�)��nz���b,6BJ���.J�셚� �2��ls���;>,J��B|��v���dG<B�^���?��L����T��O4*�l��d"�}�.���*��[�a�J�1ׇ�T�Y��(�]=��y�͒"�=���<M�Ħ�[��Mj����0U��Y֙���0M����d��o�*.rS.\�ص����f �e�D|�p*�g�s��fן.=��[�M�8�א�6��W��E��5Ç��Q�<*��U H	)n�E��J)ۥ� .ϖ3��RiD���\y�/��-��db�0zHE�����Iߋ����>y�͉xl۝G�C{g�.8���Gi/�kxo0Lq�e% �h�ol���ˀ��޴~��Ox���ϐ�p[��b̃qz��&4��3��gZu�X}�Q>����B,�7�Ra���ܲ���� ��}��C���n�x,)FMUD�qu��f��'W�ٿ՘T=����v��5ƞ�$�z�f�S���}p-�x�����C�֤̏0-��X~x�3,���n �4���n�_�NBF)�;@� ���oM0�b�B�)����P[�x�8"ӫ�g����6�A`D,|R$��.ٜF����s���JD|����o|�/I�O4�M��_tp��Z�߶�εA}�s���|�~�o��Ӂ�����Nݗ�Bnͦ��c�tɕ�5��������Ӯhe�5B�=٥i�2Mj��x:��	�HH�!L�K@�Vskf�9�8�I"I�x����Ĕ546NR�K$Y�MKTp�֒���ٹ9��8,���N�5�x�ģ����C�y�g.��9�	X��RG]d5>p8�=�7Cˬ6(G��Ա�՛ �yDYO�4�}}�qy��[���1e}�f|v��W�}�Z�滠���6$�W�Ip׬[6�X�.�|�͛�n��ʇn�"ay��0va�ވFE�-{���r��^.q-��$�m��''i���3lrɺ�� �W�����4�������>��ʊH��Aq��X�+L #df[
)�G�s�!�$�YD�.*�����j`�v2��uW08�c���N��)rЅ%�I�wqVe`��f|$ϴ ����DK(�v�i:�{C�Zז\>��C��ށ�UZs?�_��g�X���?�_�TA�bA�`�$CF�C��i�����k��pG��'̸��6��D�9��N��!��#��a�����r��|t]��/Ο#�5��-��l)�[`�H�5�ʼ���ڣ�㾘e�T2}\�ȴʖW�3*,y�u��9�&��n��9W�5����<U|��W��kM��!���>����C
�ɳG��(��D�0F��?WX����F:��|������9\y���߳ߛ{�/ًz�PS:P�d��;kwE�k�H��h�-�n��о�W�����Gb�
\D�\����ٞ]ʱ�yMF}��Y��t	2����z����{x 	i�AB�$d�N���$�nj(�A�aHi@bh�;����ֻ�,\˥̽�9g�����{Tu��Mˠ��6�=�[�Α��>{	���~
��~���M8��.�;��?�nZT��{�4��n��4ゑEA��iY�٬	li� �}�O�|���+;! �ѽ%ƱV��ݖ9Lrpi[y_L��;I�+E��dgc�s>:\�����0+ʮ�W-�����;2��p5���8�mݬWTh E���~�����k�\ |	@��+��I�Zn{a5?�4LĲQ&%ג����/�������w6K���N�Z_g�o9j���v�l撒Q�#��f�y��l���A�Xn����"7�	tӜ���U$}8V虥p��������,�������
��m���ˌ% ��q�)����-���}�v� ���Z�6v�Jc��) uЍOt�n��P�N��F��N��J$	����l�^H�!�<�.p���ˬ�o�O(6�ɥF��-����s����k傚\Їr
A����݈ܺ�!v�i4�o}�u5�+��ɔe\k���}��r��I9sc<R	R�a�M"�?P��uz罾��6��3*��\��g�����`����T[u=d�$�n򗽫骽%��O���U5?�L�O\y>����흝����+*R<z���tP�:i�JBǹ0h
4��)X!����GE�|\��ª�7���䤪�DR�a�����7�]��~��HSHų�N%����/���z�3N�&�����b��q�G3""G<Q�F�g۬���������D'E�qڻ�#����ӌ�3�@�m�*O���{�\M��r�,�+>B�T�B�Hn��7.�[�&ǜ�CO\�C�O�@IQn%�R
}H=,�@p}Ԙ�A��=�K����f�ţ�s?=0�H�)6D6���" �4�N@�1vs�z:���5f�Yܐ��V�Ep�6h>�
lWQ9ԟ�����4�EA#����F���	j��s��9��k��`T�0lɏI��R1��9��*���B�}]vIf��Ō�ۋ����CW���t2^��K�ʥ�5	��}4]��}gi��x=���V���j�fa�\�༢@��x乱�8z!�5J<�����5�q�^�s��U���@�d(cY+U?U�QO\<.9S00��1;=?��<����+��출�1�B%;��O����q�ƃ�`�uo������c_�⁂6E
�}�/�Fi`�x����K�~�4�l�_UK4O���];�z(�%e�G��$Tr"֛�Ӻ���l���6I�i�QRD)�E�THm�/�\�g�"�I�-�ve��?�zX�2�]U��?��l�2����=u!�NƋ���ӝ�4�P��s(�L��}}Fm ���b.A�tkHT �ea�9��mT�`ց�PO9�9�;�3�s�5����D�����<�=ow.���Ѩ[���#��>�׬�b0��
����ꁾ�ؠ_���)g�g5��U}Zsgb�+NI��/��4}�zg��NtW�#]��Mѷ'��:����{8�~��@B����г�ʴ�{	4�_�+�;��V�����%Pb���J���?�l��Gk���9��zĪ�&�;#��<���N�Q�P�ב7�M3����ƺ�yD롁1Vr��~�N�eNZ�?W�~�	��r��H�y�p2�#����4��w��X���ý���l��\O���=c��gj�=HX�}*l������:(g�<����j����^wsI����pffj�!�:��)�6iyJ����T���Ix�����Ԏ�-n�l۴�߱sj����OX���/�#�Lg�(M�PX�5*4p��.ژ�3�% t�9�����vF�8�(k�b����2�q���N�?�7TTP '�x��>4����
t�*��)�~���[�cd�iȎ.o�Q����ϛl�!��?sj�m���} 5>{�#�Dp��`�oʢ�ͭ{A��I�A)�A)+�٪���$�O�[˘G& �A��o	5��W9�u-����PӉ_䴈�A�W��;�JkS�"3�����{��,�����h��?,��j��n!Y�����>7L�	��l?an��_u7I�Z�:��A6��:�AL�ϻ�%�3"Z��J�G[j�b�|=r��b1d�Fd�#�k$봘j�T��$�`L��B^9��T�	��@��pп�B����2���-&�H�OZ
�uZ���伖����d����#�	0��ʪ�B@��b��>�,$�tp�lr^��,��4ir�I%�&ű�.�r���eY�ke�u��-u�l�S�Q<�DlJ�4Az� ����y�Ćɿ���4�u��ܹ�
�$�;�ǈ����L�:������[��x�����	���Q��;)�h! �H)�<G�����ج�)<��`.7�V�'�6C un]�0)LB��� �[�Ş
<S��pd�+L��7I��6�� ����I�,�����X�5��sw�V��Q�Z�9�e����B��[7�`𛶪�7�k�@���i�����{��xRm.H�Z*)8�~�����<`�u�4k�ݾj(+���W�kxTv�eE��R�$U�#Nbf�npϭ�z��˻F5��X	����b���Zo�~�!��B���_���;����^��$����(���
� �0��s�i����Wtq�k�w�6���u�����)~�6��R��pU���IHB6�dk�P�-�PB5J"


r���	 "/�Qz�=�&��{��Pc�m�'�c�A��^��uǓ�(l����M.p�l�ӳ3�����ٌg���zO��ƧE]Hk4�X� j*�R��f?T��Ё�=��[��ǿ
�L���ks����ؔ�B�.���o����U���ُu6��9�U�/'[s�</�!C�|���n�Jt���7/_�b������m�z�C+�]a �U�'�c�&���Ӈ6~����%U�H�����i3���Wb^cʟLv�~f�,�Sm���Т.ZV!��9���'C��V��@v-U������i_u�ڦ��w�̼�Q�*Ii�O� ��32�7��ϛ�H|3��9�E�j�aa*�$�k;�����\������ט]�� ~������RF	-Z�94o�kr��]ރ�,hmx@*l�mmmG�����ʮ��e@VлY.��*�	�['!s'�z�`A|wA��皔�������7�Ķ<�@��n#f`,��]ť��ٽ�j����%O�Ɛ`E�����:��8��|?S-}�<B���"'�="��;!�A7(�;:]ctttQ�X	��|�S|XXX�L����8񑶺u�{�c����Ùg��[y�����iz@^�I���6��U��"CI������T�|��NB�!/�����NH���{+�ݰ��|A�MMk߫z���D����p,� O]gBU{$��+Wr����)L�]�����<����2����SBd�#z^��[�
��j�/�=���K(��Q��/���돆��o]+BJ�����ܭ�|{@�Jg2�0	���i����m�á[�Qs��ɰ0=}ў�Ԏ�8|r~���	��˗��s�ǅ�o�M�zoQ]2��JA~�,�]V�%j�?g͋�i'XY����D#( 8 8�wr�� ����d��5oJ���<m�ʓ�kM��V_� ��i�M�)��y��k�2��e霾��gf�1O�|fo�E�x�o���'���Ҷ>�6@T�7: nhSc�fh���<Tu����4�]w	�ԫ�R>�]���Cz�� ��#�$�W�ˎ�mR����CD?�]�Ι�}������M�7���u����S����:�6��� 񨓑#n�Q�dh��yq�T�<�o�$� ���U����<|Y���A��8d/L"�m�=4��ʑ�)*@&����>a/���'���,>	�P�-�Tn�ET ����+�K�_��J�M���r�SQ�[l��n_t����s%$ɸ�cV_��Q�X
�l2��[X�G��[
�461�EǏ�X������WN(�ա؈r������ݷ�V��+u�Ʈn�UC��@�a7�]ݰޞ=�:�r� ������� 6��B��v9sDgY ��NQ�o��� �9���1O��t�0�B�Q�G~�����4������Z�4���LkׁҲ�?�������L��_nRmS�H޷��^[!��=4�O�\r�5�#|���dh��	�j�{�he�"��aQ��y�k��?�GMq�b|+[���yr�����S�7u���F"±pC�I&��ۄRu᫣��ܙ߯��{&tÖp�;0����s��o4��\]8ULL�\	�LBx����Ϟ�.�c�m�r���黖b��,E�`%���r�_ ?� ��j�q�~�!���O���p��tc�n"������7�-�G��u��8M�u�UhR)3WK��8��t2hl��X�2A�h�(ff`k\�r="��j�.��UI���|/�۫�⸃���Y������F��p��i�V=�-Mp�W�|m��*�p���i���&�� 5�eB1C�D�F/�T��WM�䊊P��8�i,����̃����T���/�:7̑��[�p/��=(t����G?�l#%��7&�9M���˃A2��dpe���yϿ�2`Y�Q�¸�|d���~k���B	��$# �41����{��B 
&tn�e~��}\���،kF)�k���GO�����U;��}��L28��wq�CmpV;���c�,��+w�B�h����9��B���Tz���l�����<I��H��� C�w��:WO'1�|�Q���$��wE��֍(�[d]�Ǩ^�۲S�{��%u������
��V!�R�{39e�Ї
��2�y������p��>�Yt,@�]���_^�
N���k��6^vi�AhMW���g���);/Ӵ�U�2�>{����Xމh1%�,���;�>f�}�6�����������^NN��W�v<����|�����h%2V81�,~�6Q�f���^	H�
��F�W�fّ��R.�L~���\	��Aa�2~H\�QP`� ���f�=���ǀ�E?I5v�q�� ���||`\c��t�({�G�r��;99�hR&�,�鎛��ǺP{"5�+�<�n��G���|��]�_-/Ϥ�;b��)޷�:�?G��1�c���A�*~�Do_�Ouh8��*��N����P#��k�w�I��>�IBV�Rq����~�,R8N �,�rq����\�����i/Î��"N�=��!�%����G����J����f�f� �.9�\]-����nNɭ��
��:_�o��o6�����uo�t˄�e��wų5@;��X����c0�;�Ć��ٿys�����E���^��t� ���a�Csa�I���yMr�4�5�g�ʃ��F���O�L>�E������TH��ǣ�����"���2'��m��1�}>�iL
���;��O�(;L�@�����Q~�L�Oof����8䟍?QW|	�WUh��Ӛv�T�^]��%�5V��x���G]6K�e���RQqn�yf�H�EJF+�����b7tCvV6���SZF��n�
�"�c�<��b�bJ������㲦�?�n�M
�[��m�P6O>!4�>4���O�����?씳5F�.)�%�ļ��1��q���)��sp�Ee_�.Q�B��=i����R���Г��F%��hv\r�$O���i�n9�_�!@#� ^� NNN��\��������PD[C�`![�m�ȗ)9���Xy�ܓr�k�ޝq���'&�ѻ�5�|԰/�;�R�Î�
��k~� ����hr��"�"~hW�PR����g���a|rhbPe/�Jp�ˠ3��i�q�p?�+k{���sT|��8��[��H�=k'Պ��/���1JZ��F����:��,x4�:%��P<�����z��~|�Qb}�1��i�(k�R���/�l$�K3!�ε���ל4j�(P����Z^5��|щV��6J���in%z���sj�ㄏ��^[L����UN����T�y���lU��f�V�j���η.u���}	�Ʒ���zog�d{ovw�nd�f�Ld��,�������l�I�v�߼y�ή�+���Vu��T+J���,8S�K��}I�O�߸����I[/���-A�Y2^����H�'S��i"I_N�{�k%�Ŧ�w�'5s\�&�U�w)Ȫ�bC^%��.���v���6�$![aZ�W�eӎ�(�P��s �wn/^�=9��`�t���
a�!�I��\#��4��Q���镶����m���[��������7ѹ���t�����/k��̭��ٳ�z3���!b���o]� ���:5��֋�p��A�v�C�}$K!M�%�u3/4�K>�+d
(I@�����VTXx2lU��z<��L�Fûn��k�����?�.������3�4�2|�z1����wQ�l��i�r��DE>jz�YvF�����j%��ҭ���7�HA�W"���逕�&�|_cu���gJǝ�M~y�.	h�ݨHb��!��s1���k�Y�	lT���X^N�O�-0�=�O�%�OU�2��CG?�rP��U��>���O��'�����։N����u��P�������-j�`DթLbT>@�����������c_/�Ȕ��{�ͺ4�\�����.�o}X\�0�j�����#�D��/Z�x�mb&4��qQP��|m,�K_e�cUAﮣ���\\�dj"��k�-%H�y�C��ی���sE��Qc `��b<pq��ɕ���h��������҇�%T�ղ��u��0Ic��n�[N���i�9?�\�D�jQ�c2�"QU�)%���@�~�=,����pwx|�{��ռ�5���P-��k5�'�ۻ���|&�M#KKz[����dc�ʏ�;�y'�y'�F���?%�x�\�
�_e�[�?i���>{k�$a�����L���D���!��?�d>ٱ���z=T�}�T���v���ʗ �TT��KXF��tC�E�1�q���_s��)�e~������ZcL
���bM]�48 ��Ƕ	E+�x xDT�v���� �����Dۺd�X�	��(�;��HMY��P���k�X-/�L����~��`�硔p0����ϥ��eM��hհ�Z����-��&G��.L�kS�y��o��ϟ?5�L��j�z�+�X��(�����q �5���r�M>ѫ�Q�4C��*U1���V��E���{mNd��`P�x��������c��*��AN�PE`	��OY=���`�����������>e�|5`�k�����+y��O�+�	���d%�:i)�R�Ir�|��:`��ΐ�^�M�Lr�E��2F����zZ����jh���=>� !V�:!��[l0�����ZD!�Xa,8��b��aD��qz��l�ֈJX��ɮިҴ��=���%�b�p����h¤�j���n��.����vF튱?Ȕ�^'''�&;�ͻ���I���ު�z�����vE�Vk9��mM]�s�!O�|�'�����l&N�ݦ9!���FN�I��m_�0U��O�ڗi�����)�7�s��X+�www����	�+�C�M.̺�3��sL��d7.�=�`|P^��k
���AO?FT�(�>��](�ߐ�~*h��BL=-Fm(.�~�~&!���˧(�g����I���靶�OOsx��c+������1�����[E8�声\J�ˆRG��bAx�2n?�f��9v��ڪ[~��j}d���W�]���Z�:�:����g�,��t�د��R�V��+�ޟ6䇦�5������>��v1�44@�^ɋ��ڐR��x�;�8_� 1��}#�|������C�`�UE�di4k>v�j�|�xN��5+
��9𭎑��.l6��`ܛ�G����<���&�	��;���-L�E����M�C�����=���?L��,,�M���mJoHcC��T0̸�P���;u�E�C~=�c-�i�	�I��'S�>z"x���U�˽�x��pIt^_�j`0�q�ɮ��T���W//��J����̃c�R�7���#�%D [Y�XF���� �?�CY�ǌZ^��tC�<K�I���D�yʍ\2�T�ra�z�V�Fҭ�b��a��f�@�D��@��+ᱷ�̳Z�o{�PR/�f�Un�I	��ꄎB~E�����l���N�,���u,�[��j_��ϒ81�nδ#�J*�G�=|�*@�I�D�8�w�^�}A�
����%tNld�L f	���sX��ƿo[bB=�{R«{�?�`3H3 �7�dBU��M�^���Sk�X��kx���J�D�ع���"����o�!��l���6dr�U���ѷ�3\��G��{g!=�M�R��ڪq�9�^NWKcďm�Q�<rR4Eƭ�,A��YHkx�㤚�W<wT������� �z����A�m�!{^�%�_�EU�.�p�Ly@����o�L�M��}���- ��<�OeuFIi�%���� gFDK��U{�E%�yZ5d���:��<X�**d�ͯ��nAa;�,U�~{xS-`�W_ى|�؝67�ߦ�Qf����M�M��QH�����A��6�.pҳ��:���#"��@�pR�t�|D&Y>k�a({�5����Q�����k�"j�ir���'M��_]���u[Û\�Q��B���DH��� ��<#?\�2����y%�[y
�=������]~��_���m9���s<����5�	�B7سc�<�:����DR����q�����1C�ãۿ�-�?W�Y�`�˃����5�݄���#¸Q�,N>�PI�	Iφx}���� e/4�n�.����N���
�G4��|BV�V��@jJ��ھn^��ԣ��4��;� !
�?�7��w�t(�}|)T���BCU ��J�a�l����ֽ�Ԉ�s5���r�=D=���{&��'��.;h�/�6�w�M�!�%Lʾ��'�(d���}̻��?X� ��U	]^����q��� �;�(wɃ�z��������?��H#**���� ��Yl��r*:��%P��޾�V?([po.�z�A3��ъ�#6�ǒu��%#�`��<�!�2g��{��&V�_�-{U���r( �ǔYH!��x᥎�1��XZ��/w�!�4����&�j�i��F�lAb����%E��<�dn�;o0�b�6ӛWS�Xe��`�<mN��0V�	G�E�K����t��n�~�wq��FD+��i���.G�����!���%��(N���o;��d�S�&�R{M쐣�'�Цkޱ�ѯ]jx�::��k���eH��<{�?_�����g�SrJ	�/���"��nx�ɕ2ɔ:Zb�	-�h�
 �XN�'�́�u|��(�k���@�~!�7��NH��E:�����T��+��C��Fj�cƍ�P�9�~ɔ=����S�^\%�3"H�������K����
���H� `�Dݰ�%/�Oh����Ĩ�#֏eIX�L���P���T"A�)ĸ��YV���=A��bj�O9���OU|����iU�����i�0�r�ߗҋ@K�G�a��R�OQ~?a��^��%/��t���a��_�~C��J�� �v�	V
�3ZB&��B�I���K��C%D�j1�]�����x|��:����j�� ��> ��S�{gUe��֟�z�	��K��/�C9��L�*	�(	�"['mG���8J��]�0�Zj�q������G��:.��ts~��v�92����ۦ>�``SKg��n1�z����e�����"���6���1[	���/��.y��aDV{v�۩F��a��8x��R���Hf
�"���=(H�c=
�ƀ�Jc�y�zZ�a����٧\!]��:���#����?
�e��NOMn#$k7U�;�8kj4�Z}l���l��7���X�����&3����"(y�O	�伷'^����	-�Y�Ɗ��z\��@�F��U�d`�1�eQ��|��������zR��l�1ee?����-bId�@�) [ ��з~��-�Kz��}Qz�C֕3%h2b�)�dBp����J@'�,1})�5���r�����^_�:��H�Y.!l����F-�RАk�hz���pk��e	E�r;W��U��ʡ|,�Q��q�������I�i|��}X��؀�������V-IR9995�ƕ�P:@��j>#�.ɕL�S$�-�/4�����ilF� Si{�����X
������Q	���|sg�#}��S�'��>^�'W��_1(A�ڠ8����%�`a���;��/8˩��	���(�Va�?!���Ѩq��:�1i�@�~fӶ�Ը�����"ݓ�W��,���Ӷy����>�GI͊>>	����K���b�0��0��h��Fg9�/Ң,�)щ�9�;j�B�P��%���M�Ac���ئ�+F�7�-��F��M�?�Tw1p��BH��0�oQ-��ϟ��Ȉ+��0,�X������'���Uڰ�6���	��4��m�LR�ʦ/�z8b�#�)�qa4%D��Tm{e�tz��RG ����{��m���>���WW>�-��k;!'����;���\�̑:6�����L��L��<��O���&��Vu�Z�ھ�C�i	�d��|���$]�KN1A' �9�O�v�<�)j2=�~���8Bn^0��O�4N��|�>��'��l�B�������v�9+��VS$���nLR���-���َ`�cu��&,���7��k�ovD@=gqMw�5MO/~�ͱ�e}���>e��q/��Ju�-����ܳRt,�p�ۦ0�Ј��I ����4���:/I��鋦6�3qmŮ��H	�����j�sF4�'y��F:X�"��~�r�A>�s�ӡ��_P0d�T��Rou͡H�a�F8��peL�`�A(�e�ϗ�	������}�(K�Q�<'�RM&����6ο�E�������&��&���x����<Q�[X�Gކo,;���L����:��`��1cj��ŀ2g'����	f�x��*�{1H���q�F�%�hEp�g�LR\��>K�/�߂\V8fDD���_-+�R��H��^�t�[�gJn�� \�'0���]�(b���l�a3��`�>���k'wĤ�����ʀ�Q���_���?���0%Ԣ��A�+��`�@����;��xׅ~Ff����x&ݞ��u8#^� ;���������Q����y��Ջ�u�Hv�@������P���y��(/]Qz��.�G^�a���b��Lm�?�*cm4wUt�)�SU'��R˕M5�9��`Z-�E�v6��J�J�F��RY�u�ٻK����T+�xm]p.uQ�����w�=�&�#rϟc��lZ*s��P�˚	�v ,�s�w��kyF�!������v-S�,�WdX�vF1�ï)�l��<d�Ê;�����^;ҡ����V����{u� ���?��זSUfC�bh�M���ON@�eڸ�a��vD�%%%-W��k�����~�o���8�eb�k��K��	�Mz�պ%�V��� �I$](*~�P=��� �}_@�0?׮��"�/{��R767s^�	j�c�̖]C]sVT\Q�7�)��kt�g���ԫ�{���8�Ԓ�z�w�N,/%�+��!�܆sL�Ѯ\�yPk1�P�qX3�  �T��I��6��������M)�3 K�0P���g�_8���Q���<����X0����׆��G�������:���G�Y>u�9{�T����$9<XLm�=��.#G7��3�s�]9����� *؛�J���¿R�7�9d��Ӵ�_�4�2��l:@`d��W#��	i9����q�>�姖;$a�to����暭��I�5������i��E�m�e�3��(0��d��쿘D�L�w�d ~C���`������N�6��z��]�"3+A�S��:I�����i�����C�����G!�)���i�Z6��tc��
v��7<�����&�(�#�e��˂�1��s�����oO���\d�aw��u-u#�!W;�?<���QP�nG�*�/�vς��ּ�XD�$�	�2����?=��*<y�B��q[�nQ��&��l�:��L�w���oU=��u�κ;��ɫ�ցM�Y�[�|��9ph�]��s��,���E�hvu�[>�H������ff���F�[�⡦<z���ݱut�Q�z���Ö�2
 ��[��l�$Q%������+���r"B�K����\�ά$o���U�!�t�I1�̰�zg��96^��x�(�r[�9��T@�+]}`C�����	�O}�K$U�-P:|&�1����*����G�O4M��w7�}����k�t���zN��4@\F|�x��ӡ8���F�7`�j��#��cVQ��3h��ٜ�ǲOФ�w�:'�qzO�X��Ԏ(��433����PX!)Ͼ1BO"�<k�~IF�7b�,Pᝋ��&�� o��0�-YIC�0m7;hƾڅk=������G�RB���'i�4���H���fq���[��ڍ��[�
�]��A�o�_��2k�KS�c��U��s���D{�@��y9D����p�� �[�լ���Dp�0�3g�~YF'^��Qh��?d����⬶laaN�1��+C>�߭����Z�v"�&�e�Gd�:�K�x��_;w��V)��q�q���_q����e��#P}�g��D��d>���eɗd d�d =��u�@���9��҅�̘��c-��
p����h����cZK�����!�D���^�������WD@�[@�!x�c(��|���q'���p�\��å����w@ج!�������C(���vr���d|p	
�2�0�.��n'!��0�
��=�-dk�{"P�}�Z����wV2�<�{o�6[}���A��Wܦ����u1�L� �D6+*�H�Hˠ��_Xs�\9�" ��?�#�]�l�p�����+౞�26�p����h�Ӌ `��&oH���)j���,�5�\��Co����Sk)�u��R�~p�3 mJ�������[N��!��b����1��^��a�L�.?heL����_����W�	7kԠ�X��'��3o�bMg6�8�6��ﮥ�m$��1EFX6y�U���{�I�><��~h��.<�OY-�j���k�h����?Pe־��k���m7δ�'M��e�R�M�׏%�]��1r�9Z�#rg2\@�_cGQiHQkz#�?��m~B�V;kX,b�R(c�6c
�(�5���U��E������6���7���ki D��՟��o���W1ʜcۏ��Bg�`�|�n�<sNn�P�wC3ghH�!��w�� ��ޝ����z�3���ŴL�z}c�pѥ'V�i�T��%��Ѐ�&=��?n���h}�x$��ʥ�]N�x�Sf1��b�=:��;� ~δWB��7H�C)&�ޚ�.��9���z���Va,�*�nV�!VoT�B��V`�k�A�.��p"��x�h�-i FYoy������0j�9��<p\[VqLC.7��GԄ+��5�W}�W݃��^U��ޞ���J����\n�r���\��I�R��+�k�q��\�6��_�å���w@�?$�0�-c$@$;��ks�vK���L��NGb#	�m�R�-� �;oe- ��k�s��4��4�@A8�Ҏ=|�_�:ܷ�
w	�ɦ����~ӑ�*���Sy�~���![Kv�u�iV�s��`m
��b �m0�SQ����r����$S��xrq4Y��@���zVV �R�d�^�;v�.���#��IJ~C�w8x�9�;��~��Z��\��`{�0h-4=kɑ;
Ԇ���P��b�#�*у�.>�����ĺ:᛭�;N��������,���hZڛ�4����a��X��F�\'��G#�j�G� �=���{�Ӟf���݁���*v5���uk_c��
���{ԖZ�t������H����vl\���3j3�GL����������ST�M��lEsO��+t��W�'ы��rF�	��p$� �����dL��+�F;����nx-Jw b��n;|Pf�:>��EA���U���$�����ˇ�0�I�@MW=0����j��8�]lR�h�- �������BEͥ��"ĝk�y�2f�0�#�a0	迨_�;X־:���f�5�t}��ѱ�tg:]�Z&_���k3}���@?�E^��^�j��C'7�����^�N��ҿ'�N9M�E�_%Ch��G���2!�"݊��i�30s��#���#�����-+�'��ڕ�PUd'Z��{�7��;��BN�La�w��M��;/\%<��A�������=�(��?rE������gJ�9�����a���KH�ʮ�}��"���RGLVvm�����+*�<L3�.���!\�Jjc���ic<kJSx%H�V�EC�sG�8椯��J~W9�_��-����̝a�kw��ҋ��d7�*�3��e  	v1c�0Z![���џ���m���j�[z������{9���um�=���p<V9��gטּ����0D�xr{μ�sCC��<}��Yu:�P�k,1�{��)��ِ�߭&!�o��)q�Y`L-P>��oB�U�`��(�wô�E+Hħ��Ƭq���z�ى��b���׉.�⁧o��|�I��D��IA�t)��x�37
�/�W��0��Y�_���� ���=Y����S������4O��l�IO����+�QS���� �4�l]&t���=Y�ɀK�-��ohl�H��\�t��,0?��މ"�Yg��Na�9�R�ow��yѓ ���n�.xbS��D�3I�D��\��rJ�q�f}�@|�6/�V7M���Sn�0�x]?$���n?}�_��7xyrl�/	y�R���!{l�A��o�C��$��mf{}5�x��J���mB���苨����HRL��ba��g����,��7!��̙_#�x���������SCW�9@�Vu��)�f�]�
>|S��(�-���YXZӤ�*����wO|1^�=(���~���!��kAm�Ϻ�5��x��sȅUa�����*�#(�lN�#��))�᪀�21�K;??�B���N�u�L��C^_���߹�L[����s���4�򨃇���!�'5s�}g��,ǲ��]Tw�.Y�$C���L�2\�N_�)�[��:��o��*=�[<�Ů.\����o�������q��o�2�|���4=]��C��3g6�H �P^3G���!BXv���/��>�jh@����fɬ �L���ݱ�)��)Uԡ�J�TO���v��a�K$�G�K��H�'�j�Z�Ydffܻ�͝gp�y[l�U���*���v�Q8����U�J��v ��%mL-^3\.��NX-��U4e��k�>�*�hBe~?橖a~3>tk�o:���k	O�Az�A[PK"�*�a�X�A.���k���������U��-(hYh��>D�=�W���A:��2K4�?������hk�C[��9�Ԉ[������]Ħx��Y��S��	x�2��x"�������>�@)�|���)�	���؞Y4�7�
���?�9m��X�,���-�E�<��[GC�~�k/�D ܙ�h5�����XJN&��3�I(�+aj�]� �����=��d��g��K��ߝ��)�P�?��};04>�{zZ�-%u!�'&��ݚ��z���ygY�B��
���˖j��nVIB%�k�ػ���/�H �����e�vvv���|������u8�Yo�sv����� �V/ Բ���LBM��d
��4��拙�h�z{��9��ڜ���\q�֤��['&�m�)򖽏4Q�i�4̩���HN�B���2Ȏ;��d�& �������#�H=�)���y��2�Ϡ����6u�ߌ�[�0�	H8��~�=7�)��
�[xYGAr&U=6�fB�	&a�v�[�dn ۟���'J��]Ņ/-#�ȭju�"�[��8�h���mo]nz�3;`ְ�����d�w#�׬����]m�`R�u�JCQ��j̪o��%�����~�1�I�� �,8�Q��`���뾻��K�@Z�4q�Yp(L���*p�� !l����`}�,���5��Dc/��Z@���R,G8~"W���87�V��θ������ �{m2��:���ﾡ���Mi3h7�]�e�n��gri)%_Ư48��v� ���r����&�Ю2���
LPCcP�� ��'x����Y��ZAt���c�����|�z�F�\9��cM��z�q���!�Hab`�o�3��p�
� �]G���W��G�E��U�}�ߟ�D2\	qj_bI���d<�K6�~���u��D�aJK|��(��Q}�h�Y�:F~��	�{hx�6on��O����)SL;��$���~S�RՎ�C-F��ɐ���m��|��S�M�T=��"zXd�H�˞��;��e�&X����q$7���N/-� 4.n���_�Or�D?5U�y�4''G7���]x�t�|x�
w�B�uͽɧk�lRn�յ�"i�{�W.4�x���0A9�P�WT�a�j�0� ����cꬣ���pOwII#��� HKJwJw*1HK7Hw�0")�5J!�u����]��_�>g?���y�6�e�h�7��W BM��Z��7�v!������V�3���7r�dC'����#�1�0@?��VBҡ���d�	�͕���������VVW�����P���ν�h�m�#�p�v�p�O��F�.��Ƹ��]�0�x1�L��{�)*����"���$(�LX�]���^��������O�Tx�I�2I�3"������2a�4[��ޓbR2�[��;I'?��p.m�F�z{�&��f�f/5�&�Ɖ ��9ū~g-6JgT���Z�]� 8��k�ߚHk/�!�*1L��`�J�n�~�F�c޾`� �m�Aᖡ�tHL{���b�I�]��CQ촻ι�3�ѱ��#f�I*P�d6�rb����$5oK	����V���5BBB�t�V�^R\\���Y�&���^I��G�����0%�z���.,@��$�S���A��F���i��b:���=G���|�:t�t�qް�Z���O+]T����BaʝXI�U=ݖ���V�.�j�e�2�z||<���J"s�n����Q��l��T�W�ZMW���8�S��J��MϏץU��A����$	�{��v�A?�}��<����0tٓ c>��ۓ�{�$��:֎���3N I�=��Ņ\��>�JC6��$J3�!�nq/�q>�Y��-�pst����l���@t!��<5��B%�g�l�wwwoo{|���n�.cu%C×����E@A޻�~�C��R�s�E�l�P�~5�dQs�w�`�C~��.��D���fq

@ךYv�v��e�g���H���H7!үS�k]l�41�^|Xw9����G�w�~J���z�tݟ�UR�����7�LL(Y���PO ���zh-�����0�Z��]�T�8a6h{6'~�y�J%��� y��g� ��������Ɛ[/��R�p�2�~FA��!6��ɩ���"���ӽ�n�m���I)V�UU��ܚ��TI4R���-�d®d����Ll��]���N.�p]hm�������I�w��z�|8��YY�@� x.�ñ����`�����c�:l�f������˗WN��d+�RdmPu��\!���D�	|E`-���{A�̉�<��a�e�@�B�WK��>�*��D?Zi��^�~@��Ɏ�AZ�Z?y��ۍ������Uw��O��;Z��:(��AG�����}v��Öě����ℱ���4)���/d�b�q6�- rG�4}Э������Z"��em3�%SNR��"�!�@u�t���z�G^(�����J���b�	.�%�'UL��^	���<¿���ȩ۪��^3��f�"<�#e�9,��rU�A���,��W�o�/����
�=���HB�i�]�p[�-��<UT�����<�Hy>.0�5���^�7'
V:��P�����.�|w�\ט1MӭȠ�UR�������o�N��U���/�\�ŏoF���gR�U�Oȳ����[���=z�p�|j7�������g��_����Q���L ���o �����l����pӰ����9���F�)�{�'�����'���6 �ܯn�txޮڈ�j^����"�y=V��<ipp�%��x�O����B{t��V�Դ�H@oV���]aV�2�)��2&($d�Pc(�9�ǫ��7�����R�Ws��4p-`�V�F�n�Tp9�|>"l�Y�e��%�Y,vd#F��^�"�z�"���ڏZ�:悆�_���m��h�E����4 �_m;�rE�@��A�6��X�����kiC���RÂ�W��"E]%6%Q*���+��v?�%8<E�jZq��]�9�����"�g
k����mo�~-/;��+f�X����.�(p��K��,)/G��/>�BE���_�s��4��������w��J'�)�YVS��]8�����JoL!�_��0���F�9=�%1��>� p"YOK^�V�[_���Ӳ�[8�5g'O=D��	�b�>/�`N�^-l͕��6�ɰ*Z�8�9�R�x8!x�%�!Zs�`puM��EY���=�){s��c��7qO�2]�H�e�T�(�8*�TՂ����|<�+	�L�98t��wvv�q��a�D�ʦ��D��O��/�ۦ�sw�Z����R�g����Q���H��<P?����KG�̓�����=� OVx�~�+u��;�͌[�L �(y�Gݸ�]�6�����¸^��M����cMk�!��H��T��DZ��S
��tqo�R���d��U*Q����<�#����@6Aj��hg�znn�r��rX��V������ôx�,�,�vPȞֶ�4�XYE"m�ս�H�t��Z薦+��M�P~�H�|����V%�������}����D�:kq�jl��f��S�Fx�t���.M���y�iA\&&�W�)��k���G�z�4a��p@�xw�\J�^������#�[u�n�+�x����z���F�֨n��W-��&@��)U�&=�S^� ��	ּ�Z�� ���m���L�&
��my̟��\gi4����M���U��J��pw.���N�[
�'��:|p|���P��7�/�7�d�]�2r����aZ�1�	|��:=�)���S*]� ���-;ꍭjWgd_M�X�8^5D�ʺAu�lN}���~���œ7���r]��}B��,;1�t(oK������h����~��%ϊn�k��L���]�X{�#y� l�:o"�*�pC4I�ʊn$�<���(��:��m�n#���Ŵ�Ɋ��\�&���|��'�Q/��7�1� t�f+����|��8� ㌃�g�s	2n>V9��~ס�L͖���_�$M5;�Z�����r�x}����)O�Y%����֨�W�/��͑�[��w���]z�HB���$��@��\p���ak<�M\s������z�S�g�
DZ��L�f����?>�[�7�R'�zo������O^�5Q��h"��*r�׻���p���<�4ٍ�CN'��*����Cg	+��8��ڔ��I\5�]`a�GhB܄��{�����4�&[̸������U�Ws����x�����Y�Ԗ��串Zdw�������^U����]���p1���'>�s���wk���K��<K����No��a�x)n�jIx �8Ց
ӫ��Э
F�-a�37s�IM��:��&� ��#��nx���S����qs?�Ϗ�~jv^��N�܆�;�ݴ*�5�1�ŀm�ukTڟ�C<cN�BW�:ڄS1[yOƠ�d����ʕ��Ծ3>����~T��K㒕������/�5>����E�C1��÷k2����"?�:F��ٹ~�"����e���_f�t�.�Fb̶GнY��������T4����iq�#�#�����'GflD�6 �p�Qﶇ�5n/ �ll|���]]�Ym>p��|�-���4F��b��ZT?$IL�[�5.k	V>���kz�sF8~\�������1h�O��g�� �{��eMdu�Z=uy��Z��biΥ�=���x�o]�aUm�;�r�q�Gp⍺��LF�к���J���燉����}�_E@�mA�XJ:[^�ԃW--����� ������t��:^a�!6�K�ȇ��.I���8lf�C�w���g���K����R��U��Aa� XokkLc�b1i _}��̋�р�_�t#������;݀�:���ʹ���:E�T(�x��=9�^������Z��O�ee�����?�NNN���KA�
N�UVa]4n�~F�r�W�Ǧ1�;z���Ӕ*�[n�jtQ5��t
5K_�q��u�����rV5��=����^�����٠�#�O*E��[�P `�����w��P���9�]�]4fe1~��۶�6�=����#w.�&����--GЇ=������<���.���,�l�+�1��B���<���E��N���΢2�D5x��j?��'4�v���b��=�������ޖM��o"5�G�f��E���
A~���1O1YM�Ep5�c���p)]��~e�m� X�S0^ɿ�ZWŞ�鰁B��!!��b�N'�B�v�,rY >�.�,#j�ȇ����0E$�JP�(��?^<։�9)[Z���Zt��|?�Cl���)��� O�����K֢��M��g�6ݹXݞK3�bZ���B�i���Qf�ݯ0�yYl�FL�u�{�Ϧ�I��h�����
�V��1�������]��:�@cD�7}�E�ET߻O���6.�l�0���P~4�}H���),�����U�͠o�'��5Ӿ�߫���!>�c���AS��T1�;��v�����aVO[��)���+]�Nɛ�
����R��?-�A>b�b�`��W�W$��xZ;L��s��Z��/���v���d���[������2G���j�(1�`ɵ-�M0�3�5Jn9y�[Բ}�.�Z9�$H:��0���j����ٞ�?���nL�n�-v9���yL���!���� G��lf���Œ�w�G:oߖ=�6��9�f�C�ۮ�1����~���^&�ҳn�~�=XoT��[YM��Wb%�1[w��y.ja�����"�A�D*	f�z.7�����F��J["Þ��ɩ��H�?T���?�wq�aF����l+����ٟ�f�pxqm%�}e��4�*�����j����xYL��ug��&�s^�_[����b��Ϫ��v�w9ҹ�ť�
�ޢT���JJ�XXXM~�~h>>>�zO�:y�~�^о#L����/�����k=�Z$�k��K�!�����m�^aXq�s���*�#��(�5���lD�W�je%�n�p��Y8N�}�/������� wz.�Uiߎ@��_/W�����P�ֿ3���?�0̜Zԡ�0$��z��~�ޢ���>��܎j̈́m�yi�6	o%������X���|Z/�nl���%h��¾Z���-<޿�'����?��f�)�|d�K��UX&-s�͖���]�D��ӿ~ʆ�k�j�b�W�9H��. ����c�}��s�����IF������7�*r��j9����>3��c�4)�n����Ϯ)d0Ke�#�*nnn�"'���9�I���=�먑���\WZT�9�Ux�>���Z"	":2�}@J?�<3#�|D�\�M���T{2-�lEv�����{��lq�{�Vv��@u�+V�DA�c�o�O�i8��߁��Ȣ<�
:�d��=�[|��`�-9pz1g�z���
�O]��]�fEU�	eP�lN+� ������Do�
O���}���� ���s�d+0�(����ڬ�,���Ou[��v�q��E)xam��Оg�^:��HH�0�x�b�CR�b�;;�ǧ�l�{c�>[���V,�"��kK�ļ�8�4�Y�%��ɐ���bn8&<��]ȥ2�-Br�刕��3�<ڗ�ه;��Q��5�"�a=nu���aE�/x��ⷽ+|\/�q*Y����d���4Qޢp�A6rr��G�_��`�������Eu�!G���+����/��qS$�{u�zS��8�׳�L�����Q��8X����0���Od��B;wՓJ�N~U�&p��{go��K�L������:��Q�比�6���,�##���h���i��F8
�%%�9�팕%i[���j�����6>]-� n�&����`�7����P go<�[��5���?�c��ÂYL��?�7�KHh`��(�98��]���|1@�8o?�����kH��aZ�R������B��b��ԩD�&)�g��ի�d�>�G�JË��rU�vs$K�Qd�M����f�vA���i�|>XD�B;���4S$����?��8V���`���(�մ�o����(=��B�6AA�/e���u�ߦ���`��~�T�zI�)\#B`��ը6�#S����g���%�;u����/��I�ڵ��6w��96�{�q�!J��|�¨��I�C�ʝ�f�a�ꇂX鰵燳O�ڶ����{�hab�[?u�'����'����|��$m�8V9W�=�[���L�?w��s��%>�莹ڪ��$�i�����.*�28���i|qk+���'�Ү�7L��::)�E���Fꋍ�8?�^�$�\�N8�l���	`�����
?Y�D�����F̤"LJ�
���f5n"����f��B3���x��Ŭ�z8�Y�Z�/=et�*G��z�#�2=����J�D�	��|�>	��a�NnI���Z״��YPqW�!����E�R�����n~�Q˳��Μ��&ƨ����K�I�wV t����.${�y�����:�T9�Щ�w,6k�VU�K籖}RF%&N��뭎� Rn��'����;/�J8\'{�H�1�5�륈i_($�b�"��G�H>Ċw�����M���IN9��4����.���m4�,�����q99����������_��h���ԇ?�p+����a�j�p�n��U�tj��Cu��.���W?�-Zd��v?��hE���B5��Fׁ��N�t?<tے1s��_!�}쯷pބF�˕5aj�	2� ����`|���GV�3� ���H��~%�Z�����\*vTd�^�k.����Z��ӓ�RL��SRPx�QK��c��i���1 S��_ֲ�v�ק����-�uN�uy�q��R�tt����4�,�)6��LފO� �Mn�k(hl
�\�{'��~����}H���V-:���ԺU��
0���|,��������� �/���NZ�o���^? ��[}=�׷h��J%��Aj���H�|��>�M�V?)�!QI�5�|W[�T��GF�U���g�s��FD�8�(>�'���{q�7����T����2'�
b�xwI&�e�f�>[�W�6���!3�=�
X;0b��>	�����lж�&�w�WH�
�$3Pi�3%M؏��(�@EBġ�^k�p� 7�F�h�����DL�5���.��{?F���!xc�����z�T��6��p��ʨ�1��yܤ��br,Y.q|�b8�1`�Q��'�KZ�UD�R�g�7ʙ/�Ӝ�3�4���Վ��4���y8�܏ ��8���%RO�[���Mʤ���4���@�e�'����<q%u�D��FF�W�f�~�&��EBT*ۃ�g�NS.?@f�s��p7S��";C�3'x��Pf���.��`J'��I���F"/�6��u�ʥ�^�� ��蔹?yq��L+E3ł��8@��
�/S�i��|KK���=�J��j�o���E31Z��%��_�Y&|������+�����N�]�C�|�J�jkk �b�N�|q���3@���}��1��_5��@O_�s6j�!��Q����@�o4fu���� F�����śs�_��l�)љ櫯��,�BYO���vD�Sf�	�XS]��lKf��}̺��lCin��U��6�v��@V⟢�Ĩ�C�/x6�*��K|�}W�9�O!Z�վ��C<ۗT�NO_�^�0�@��o�ux�L��N���6������fg^gE>��G_�J�n�z#�l��h����닉o`�O�T��me�?����yѴ�"��:
��qk��Yqّ�~4�Lo{� {`~�7;���7�˗+�H �>3�m���BI�&/�ɜB��5��i��ᖂ�gj�����O]����聒8=��􌌜.���������&#��-]w	vUӊ��"Hp��!j,V�.�nt�\?���34'0�&���� g�d��v}QBG%�!QjC%��%#a?w���S/�NV5E�l�(I�x�(!/�fD#79�����I��&Csm�i�#_�<��6m�7 l�����n�1�+RykX�J*#
�z-55�h�C�	ݷ�����/�C��\7qU�驰�l}��5+���-��>�|s��,v�"�Zqq�8�a�v<���9+�.���(Z�&w���t�%�ޗ��j^.��4���-�϶��H�"�#��Wbu�'�C^��F�_����4+���v��n�2���wd_�Cb`���=����ɏ�jH8l�O�O�[L5�R�����v}@����y3��;a������Y�ׯC����T�ɐY[�ٖ�g<������:���AF����^4U�+�2b��u����Lԓq�,���S��������f(��o�m�
����-�T��y�M���/�t`֦hd!���K�cj�iݡ���x���~�ʥ2ƯVlM�|Q�����s#������[���Vl�Z���iA\}��w�v�wT�GSM��u���	!�5��{���;����W}�0&V���\�c?�Iqoi�����g�D���f%�g�n
+�#�sl��Ďl���u
0E��ӯ0C�Ȍ�ǿ�[�̭�<�|A���oX �W��W��j4|s����,��Ԥ�:��ZU����!>{\���e�!ĳk��7!JX?m�r�`6� P�y�\U��
�qK/�O����c�N�[Z�y�B��aԕ�4�T���e�5��]�qw��-��{L/�W
�1K�,��=~-::>�#����-{,|j��~D?;)��?,�7{�����$.޴ʮ}:)+eA��Nih�Qw��Ev��-b�)����%���������a�^�_�ʙ���� �I��V���_��&k�oɖ��oEHx���f_#�*������9�}�o�m��e4&����hd��V;�M���uV68zt�`�΢���g���,)�8OW�Su� �˘���͚~�툌�yv?[_�F��gFLɩ���	�ȩ=��1%�,�$ӂ\�*)56*���D��ǫ���v�_��c�o�Z��H7`��7��c��!V�����	�RѠ`�� b�;�n(�-N��/��ݬ�	�j���&���F�,D.��e&֣@�"}�(㷪�;-��Gۑ�&�V�D-�1ʈ5�)����0?ETtz��&�9{�~�QU��,}���/o�	r�ߌbǴ��?a���Ҳ�&a)P�s�㪵_=#c�O���
��,H$�5 o�?��?�Tx����MMA�/'i�"�����^�#˘��������Q���*"�z)�\"�!�ܦ�W�֍�u~�����e����hZ(�]�V�y��%@mm�C�|@e*�,�z8%�5��cݍ��tz�O��9��CR��6�Q5�-:��Ž�F��㯕�����[Gh�H�k_��gY㐌3����Te�+�Ͻ�f���S�.��΅�1����P#�Hx�����m0c�%PI	,~ܐ�ul�<��{���� ��Nó�s})��������!bwU�>�����5������j;�e�$�l¯���Q{�YA����F���4l�.�#�3F����?��n�p?q����{�#��gA7������i����i� �;m+��q-�d���!8љDN@O)w��s
��{�m�?>+�`!l������ h���H0��#�)��%���ʨ��ٱ����A�^3�;%��&9�'-&�>��L��(r^a4,��������o^�l�|���غ�heO�yB>�x���VaV7����^�MX�U�R����y*��1ԓjq[�|�!cT]���mꅺ����I�tl�B)+{���QI���V����	�+��낔���N�~E���ٳ�����G�1�z��H��""�R|(�Suf7%}ҥ��)u�T>6y���P	*�%׶l�sQ��>�K�??3���ެ�
�����U
�hh�U^R2��d��S���\u�+E�}X��+|����t77mg([dY[�F<�z:j��\%�	ڧC�w0�M�^�"bӸ���q���+i|/�G������6b����#sRY���rz&���d���m��;^��L�Ƕ���A���Ze�Ъ��B�?É��積���M�˾*����O���,~��(�;\����̧�u��9�y�i<i�M!9=�����|d6=C�PԞHď�?,E!`�j�6��ջ�}�����/�:t����~���>����^r�1=���+�ؓC��OP�~1~fF�
�%��*����a/#�3X1�Ѷy9">��sό�0u�V �d�A����hZ@��u]�&�0|��þ�����Q��Ǣ�"�Kx��A�aq(������[�je��D�h���i�_��J-�?�H�4'�e>#�9M�<-�V���uvQi��I��q��f%�T)t�����w�r}
*g��o��O�;L��Ie;qU[|�w):�����-u6-fý;;H��eW���k�����;�ք��Rrν�F�o~2���P�	^-��?�&:dw����u��{T%&���뎘�^ѧ�Ū�îH?"�3��n�ث�?Z~�3ۆ�L	�h�D�[����(E��hOT�w
"�pR�j��B"�7�����[q>�����>[5%Q�1�lƞ���Á�|�w��p��q��n�(Q,���7�GY9��ɐ� I͌?n�ik�dlݡ�ĩ%M�k}�,�m�A	�~��fl��5�ıʛ@��5&��Ǳ�)<T�r'k*u�Ļ,�`ں2u|�{�Ę��siiӪ7�ER��#��U�b�vi�+'���~{�(�.�zp���H�����w�#˓�C��b�����W����J�߱i�0%<���o���z����|3��� �,�WO+���O�:�>bx(D4�ncܟO�G矫��_�z��,z�� �(e�=y7t�ƛ����F8F�6�?4��r�re+�2]U��¶U�i�V��E�Y��1r���qN����8������%�~��B�{�.W�7���dM�6+�N����]��::z%J�iZ��h��o���h�ۂ�BJ��ߥ��R��T�d�K�v���Im�LߪI�I��g{SV9W��ח�0�\rBQy�i�Qr�!C-g#K������>m��@���m�w>*���K���v �5���BU�p��/� '�&g�-�K�c����ҙ���Iv�v�t�V\���.Œ/��̘Fbb.���Dh��#�L�+�����H�7�+G�ǘ�\����|~����O���Ry�6y���`ee��~{���b��=���T����DBQT�]�Azָ��`�橲$��x�ܰ��gQ�U�,��/��3����)0B�(�h�ř��i����!(7�Ƀ
��	��4oߒ�(���)<�ׁ���|`��2Q2 @�����3B֐�

R7��YYy����Y��n8�#��O�ȍ5�Y1K�1Y8rƑ�x��Ա�B�S	t?8nW�?#ocn�W:։��X�d�y�m�s���a��#a,S����,�Έ�t��k)o]�u���7Y<�8"xS�X�>5�����(�FODѓw|\y�n�y�/$��;�l��������y��.��v�[���ǐ2j�g�j�I
�ƹ���ݢh�h*���d<\��T������Fz�{�QsҴ��T~8�$���뵨&ݮ�m�5�`RO��&�w��s��k������a�%�K�v�7�^�{2� �~J�zަ�]&���/Wm� �\�h��V�d6�oZ�~�
|zFn��p�;��d=�3�7�eߨ*��nM��,�}���'�P(�#�����⇭�w���[�(b}�_3���`J,hhh>�!�E��J�"ܢl��O�!��<��]�S%$�E�O�P��\�T����@% �f�꠾������5
�\�_D�ո�1�M��.�e�IM%T/�$OLLd��棊�*%%��7	��w�f�'�K����ߊ���q��m��X+�op$"s�B���S�<;gY��GX)�]y����q�{��A~���l��J#�j���̴���c�#��t]�������p)�S�=�<㇛��n'�!���#���dsg��cc�{ii�ӳnw���'��|�ܼ���߁��W���ʨ�j4�_�8����k_��\��h��_����9����N�ڱXX�+Q0F!��_;[��zy�󖪔��sZ'�<�rGc6`��J�&Yi�`�XeY����{��T̢n
������96�Ё��.+�WaJvlN#|Q*_I����1n#K��3m���+��o�9:���ǿP�0VgN}��R���`�_�z��F<�'w꽓��ףr#�/�]�8�.�Z����az6�.~ݡ��)܋-8h`��IK^���$��l{��k�$0r���:Fe�xr��<��n��!qO7,cZ��l����ŀ�]�7x[�^����-��fr�3T�!x�����\2���-_��X�u3��9�O
ۯ�3}�Ϫc��ϑD�+�O�K`�~9��{ ?�є ֈ���c�2�՘�-B���*<����Q0/�
R��27�ѿ��)1uQuJ�	��h��ng����z2b��S��[q���ɻ�N�-�F���oUO�]��<��\lJ'���oy\׽���SY#�Ǵ+��\�}$���<|ͽ�ݒ�'�M�0���Vb³�,B���˷sι`��m�ݝ��b�|�\��]89��7M�%�f��q���oZv(U�a��_omՙ\�<����OI����(���h��U�0����,���=`�Wf)`L7u;
�G�]Icw�HW�YzT�_\�#J��F�x���&�)		.&�6.X7�"�m7�S�e��ϤG;'P��6=P���.�.LcIRTKgV����&���@���x	v()�y���x'��&������茟�1rN�Q�e��v�\�Wk�&�K e8�ϧWɈy%��/���ph���u�Vru`��Pp������F��7���:�4�˜���|�x�3���f4갑
RI����h�L%��*�r>0I�`���P��~�w������i�_��I�<D4�i�K�GSI�8W*�������%��r_a`D˗ߘ$�2��R(I��f�\�D#�h1P�5�����M|`�t��$����5p��.-M�����8{��p)�=�\^ ��c2��%��u;�|�5��~]ը���{�w�u!U,�%@_\�R�'w�-S����It�sMM��HD� -�/�*B"��4��y˻�1�$	+?Ne�f�����}7d�v�F ov�oD�>tMJ���?�O�N�Gt�k�m�$��ߊ�>�A������Mϗ ��'�y ��gHSI�������
�3����{qxj蛔2=�=s�SE����5���Q�[�S�eXPjs2��S�g�2���(�^���_��x������q��Nk��dw58��v^�24�\��f�꿢\�-'#^>{���I%`���Bq�d��0�n�<Q�7�D�-�r#��(��"]��z7���㧴������+C2�����3��ǲd8#7��&�?a�b��)�@H��|4����CMA���}���̎���fx�ҕǴ����*��l��x�`l��2�Fw�݇���7{:��JF����ye��+��9>��ڀm���x-ɏD1xN���_�W�gM���Ć�S�ʜ���:�I�j���c N]|R.Euɕ�Xv��駊��f��h�I���ak��u���_��;��be�z��w��	博��؝��'�BZLQdΡ���C���^�~�f�����!wX�/��>&��%�uh�؋�\2�=���"�q`Bl��o�b�a�k�DM�?�@�C�������]����/&�*���[��9@JSP�n��.�6�h6@�����o�nr>l���H�^�;07(�s\�̻D�$�/>qI��4�������mw:Ƚ++����k��|��Q���;3Ǎ��R��B��j(��립�?���m��)d�8c�� �H���ՙ�_HZ7��P��99����G��an��!\_��={q�����(T��QdNc� +Ҭx��e�1��!7Q��<����)v�Mo��e���=�KEb�y\�7jj �6Vb�!��8������2ٯ�wK�=Y��[�y��I�4[E�L���C�;%A}�j�����o�!�j�齨�?�°@Ԧ����3�ckܳ,F'-���;qX�M_�U#��F>Zȩ��ࣰ�4�j�đ7��ï�׼���>W�����f��uխ�Ґې�E���IH�O(-�c<���UG�6oߎ��#���(�Xd�l�><qQ�m('	O�-��'F�CD�F}4��Mx�(�����3yE�:��vh�U:��B�C`�r���,�ZY��	��S>�ƽ��Ƞ��& �!�E�f��/�k>%�����<DC������_�/Btl7-x�5f�/fl�g��?��4���vV׺�	����4>�����{i ysYϠm�&����D8O�ҿi���E�S���9W�c^��~���4�������b?u��N�x}�.�)w^��z�Z�sIE~�4��M�n@�>� ;
J�P���a�g�n���zCǊ�1��6c�̝���8J�cz��^Ŏ�q�6vv�����c�R[3�T�O�=��D���k�?<*ν���"������/C������έ%_�*��z���������c �xQ�U���x�b��'У��>T�
o¼�1#ֿM��N�w
}�d�h��n��|	����s����l|�y�P*��|V�k��3����Ϻ���=�B��*�&G�d˟�܅c3*�e@����T|8*�7���.Jy�W_<7���DFE%�{!E�X�Ԥ;�����
�fW�r��=������|�,Z}��,��_zz���6�9+�Q���>�������Um�q&��><ZR�[��	�5�a����[7�^3�e����Xl�"u
e,[�eȫs�|��/�4yTU�q�OG�>LP��Z���Ʋ�WuV�:A~�	����G��C�5Y��,���WUW{���]�b��J&�Rƾf,���Oƥw1|�Au�i��*��W�ޏȰv�>�P�9�2i��|����]w}� �Q�Z�������t�pl�ӓ�O��+[l��7�ǘ9�9�@X�V�9�h�S�Xf!�	q�i���Y ��r��+y�DB�ICr%�^��b.����H���N�=�kJ!���p됤9�H��qǲ�O�a$�k����Pa�ƌ���D��������IP�o���fΞVʤ������J7Ӵwhb���,�`�?�-������2F=�-���n�u�	J� ���Z<W'[]����4 W�1��h~��/@��e6;Q��6 R0�%�ց�?����-K�K&�>��w�TW���^i!�9j��^��5�H�k��+�[.����|Ww�Ea!��9ʊ�	�c�,ē
I<`i��$���[���`�hc����l����cʅ��`�hބ<
��k����h��W)�_c��$S�*�5g�]-ZK6�Ly~��YwtR��^�.���`�{-��+\G�܃
��������W��8m��r+&�uhg�U���wY�j�������b�Hp.tV���$bނo�^ l�L-��s֘�-\+�r�SU�$����U{��<�᰿X���KѤ`=��~���2rڑ�(�(�<$A�N�g*��������Q�y�q���DCn2;��Ji���I���Q��KƓw�������ឤ-o�lI�u��E|*�3��~$���G����E=ۊ��o��P�h��j�5�J5��P���x��/Vw�r�"ӡ��h�~��Ɔ
�7�^��Kӆo!�����zZ�@�����
TtPFgl�L:7�� �R�J����(���ǎFL�(��
�<�P�=yq\J�B��t,@8F��q�X��y5�I�8t��+��f�0��>M)��[;%wV�+\�����/�w@����\^�?��d�GoC�cfc��J�XK�x�i|�]�6�_����r>By�9�(-�ɝG�%d��Y�L����u��ʁv��<F�㯍�1�vFN'����%S^�$hrG�ޭ��d��Y��d���z��:�L839�$
��m�v���3����\�ޟM�`�?՘.������:ލ%#K�^D����3�Myc��C�$2��cEs�(�w�uX0�ܔ�c\ߐ����y�o��8�ߛ6��M�0;�|�c���TYd��[K��]�CxL]�>]�XS��#-���Hy����V����͹���/�����FOr�ﮛD������-'q;kC$I�SҾ�V��C�F�cO�%Adddv�%b��FM�k���=�чr�f�E�������K.�ّ���RM��	|�crrR'�@��#sr U�a�>]9�������¯��b�|t����m�ޑET�j%��ȕ�V���UZ���S���2�Ũm� M�'B���d�[�]H����c?�M�6nw^$Q<׸57�����3@��nt�I�9$&���"��8O�`"c�7�D0Uؓ�����|�Ț'%�������ǫ �h�7W���&X[�3��R�y�@%��h�V�95U}���_�˘L�[IL�v�F�R�*O<\�4'1�_4U�7op"tqj'�q,�f��kFΖ�	����ͬ�6[�;Z3�l�3�]�Շ�C�[ U�}q�W�A�J��4����!)��HJ7(��J�%��tw�{����f�fd�{�^�{��Vp�+I��\X+���DS���j�\��f�w�ac"13�v�I� Q�ܣn�l񴴴ڴ_�4��\k��X�WPOC)1�J��/JLg�3K+XI]�SlJq�4�V�� ����͋���Ew�4�(w��݌��`@:1���pa�ˡ��Z�CE�^b��8�HެT��L��Θ{s�.M����L��?�zD�����^1Y�Tڤ��́����#��謌���Ȟ��:�FY7�7�~�:ƭ�/��?�����AH*ބCB)t �����f�T��%��i�zD��6'2�d9Z\��m���F��%E��U�M�dCR�6����n���V����"~�b�����g�KM�q��B.eءy����k���e<��'a	C]^b���j� [��wF��o��=��gBݷ���x���K}���c$\N������d����翫,����dCU��㰅�%�CE�������9C�7Wz�	��[��G��W��)E����Q��������E�N���\����~Uq����B4r\�ع�5���/;;A�~B�ĳ�u�"��<��	� v�a�9�x1�g|���s�������vxf���Ӵ��q}
$�ҏ��)7	�� dm��w!�l�@	��������Ä�^���p� �c̘�>�Ü6�/�m�X�k_���C�@�Vv�p�yoS�7�l?�[���ڠ˂.��d�I���I6��c��)<A���l��H�Z�.�����h�r��(�ߜ+.n����}�Ǳ��i��$�G�k�B�J)@ &�Y+�N��ߎx�ֿ��_ZiOXR��6�n��S�/I��LR�jg�hBcʚ�V�m�%f���{��ҭ'��~w��%6~�-���#���@��D� {���� F:��(�-q�M�OG���$~�����0���k-􇕏�B�����+���"�����#�����I����8ܞ�o=*�H�,�����O"��>�p��E�����ÿ�5�g�~�-�5a��ݝH�&r� ��-T������%��� i�	���� GG�2���$A�(A�_��S���)�N��?��MtΫ�x�Z��E�������ꅐ�l˛K���LL����`Ez\%Q`6��w477���5j�b���"D,�r��y�q���'\v{����<4Y�@Ṭ	�N���D�@CNp'&ڻ}�D�����O�Y���ߖk7��C@3h%�2�0��O79e�]���O �E�~�L1�AM��<.//�65i��������Nj���|a�n:�jh�h9��7�,�.^6f�e	+�ږ@��K���r�(�j�]�uu�o&V�]��7��KR�(B,�tK=_>�wk!G��iPz鹕��$�7���1�#���Z<u]������޷e��^�U>�j�	Y��BZ�˥��ku�j�9�����8]c ���領|���9=g�j�=����&�?.��(�E�<��*��;w�T�;���Z>�}C���q�]�zIX&Pf�p ���'> ^}�<xY��(Iҵ��dp���2�<� ���_v��s�ִr�@6�9���V����v,84��W�Vƚ.��NPf&@7&ܔ~��;i��T�������;�#��8b2��g��9�����PtX�᳗�[p�b��u����w��	�QZNV��1���f���7$< �T�zSTo�@�w����hV�+�Oͱ�s��uR-���2>�=Y��7��v��(�<�VG��FI�K~�%���^�SX<f-���Ţ
r���������@��jP7[��4�JYb��@�kռn������q��<�7.����s�ޕ6\�}������=���F��
�"�!<�\��+��P�v�˞��$�<r M��0{�֒�����x��I�H-�D��=���&wF׳_�r���8s���g�Z]��)R�쒬�38P2��2��6�O�Yj	
߹�n��W��,��֛��������gaQ+�!�Y>�8a��� .K_. �����A?ɍkn�¾P�|��(��G��#��e���o{=Q�˩v�`�\+�"p���H�"�����̾/[
���
qh���TP0�h>6�U����a�V3�/f��m�V07�1Ħ��3�E�.t|	�-LCv#@���涄�x���a�3*cl�}ID����mg"�br2$o�d>�K��~Ǽ[�K��{��Ff���~SZ�#N�袎QlxQ$*�=�l�YْkX�@ ؈j�������B�F''��:{	�{
���;�$��TxuGA��4�pbT����_� ������~Vu�6��Բ��&%�"��ξ���g����YD�HA �*���N����؀������.��J� <��GM<��J��`������bZ��xL�4>	��%��3�]�S��+�W�^h�ǔM�e��+V��T.oE�3�Yw�]s��p�e��
��o�ν����@�!-���1br�]�0exX�ŀX��~I�,.�q=C�Ŗ���b�:�VPR�~TU�8̠�Q�^��>1���J})�[�0v�R�oq}���H4v�p[]���pp/Y!���(��>kj�[�
�n���y$ъ��\`��Я�7�7��̿ZG?����U� �7:{F�V7~�ˢo9p���_ ����lS1B
�7��Dd1�%��f�P����7��e$j���nֈ�p��f Ε���sd�FN�����m+�k���X�@�k�3*��ա.x�Y�Ҽ��J�|���ծ����oqj�7�A��_�s7���UiW\{��c�O���%��
����V&?(�O���2k����{�
�w\k$�R��S�qվ���!K����C�i#I�Ĉkξ4ɐk���	)���x�QY��=_�4�
�Аk��g]5����`�G(ή�� �ks�\�7���m�s�K��s
(��x����F����b�����ϗ�����V�1�Z��K�\��а6_k�-hՎ���.��,����gl�a=	z���������%��k� �(�Y���ҜS�N0�9��ȊTqD~�|�|hxۖNq;��B�w�{��o2�{�iCN�+א?9則¦�����I�� zb�z睼AXW��v���/��$�'�ِ	��.�>�4f}6]B�˖��±6 ����TMU����`�pc3���i�Z�\�U�[������J++5�T'�g�N��Ã��{U�=5A��Uz��p��!�7��gP
Y=��N�M1�0m8��Gt'� 3.+MJ���"����i�� �AW��X� �s۝"�Ķ�b�,
�]"�2��;+w���E�黠A'QÛ�a�*A���C�f,��!����F�r�U�y��l�3���B7���ZZHKJ�L	���$�p��?+�ο�3e����~b90H�H
eE�]M΂a�ӊ��"$I򰝻|	�W������۾���/��m�w�O���Ĭ����g;���#�`���3��.d:��i���^�O�ߗx���gY���y����'�Y���<1JO�3���p��yhw���H���A��k�����AP�p��$� ��'i�tS_�K�b�]��i	%�r����zܫ��x�$��2b_��KCx}��1�.4��b�?��q�(�����������VR��8;��P��Ɵ���G���v�S:��M"��z��]Gfr��M�;{O�f�P����쒙�B��߿�랢V�^�P�P�/�y/|y�A�!�6�)��8������z�t�Ť��A�Ʈ�Ч��NT����ׅN9G�X�9��#	Ƃ�?���F�E�[/ј����<�fcd\|�g�j�o�[HK��;kU������z����`�oN���{��>9x
��afV7�M�1d�W��,!k�;��<w�;�QC�333.��k>]��&��2�V�3��,��4愄'���?�K�Ar���R�'��v�OD4y�z���)�bA���2[�����8Rw�{��m�̞�GAA������$���#GЌ&{��`��)l'�b���-���]S�tΈ���f�:���^F����j&4�7��?�o;W��ٟ�tr?���/��d��pd.Q���l��r��Ǝ��`.�B�^/�S�'Q�+<�f����w�|WiÄ�~VXu����.�W�r������k��ߛL�L��%�r��C�Z8����Wٴ�HX1S� wc;��'Z��pd�:�C/U4�%��L��Ȍ��V��=)�Dgp:�|��J���V��F�J�<4���Ŋ��-/�r71%�
�n��ʪR��KJJ*�8��]P�����0V__�o���R�h&į�&ze����&O�}uZf�^�퍉[Ա]�&������^�ժ����yڗ��'l��h墆��: ���@~�����V���Y�f!�n��7�i�bޙ�r�O�=�~��g�Bڬ�2V��:$�:,YMԻ7�~Të�f}�Z�7+텕\�]����^�����p����'�&��%~�2O��	�Az�J�9�*o�e����RoŴ+�啾'��Ξ�����湷��uv��W2.P.�1u����v	�f�˅��+8���;;Ђ	��?�;MU2 �ぉ����N&���M�����1��m�S�M��/�b�+��U��{Q�m۲x��q��Z�f�_S#칓��TO��+�E9~7�k�W�w���dH�l����@5�;�=-Ƈb������j�'Ain>��%#l��w���Nm�8�,��2OFff�
B
t���m�����Y��o��Q��7�L��I�f��L�f��\Ri����e���\�aF%/�1Dh�s:/t@g��,�t�h�^a�Ȩ��3<Æ_�0E�F�	~% �%hV�i6?%6ඞ��횗_c�v�\�����:�ki����5�l�Z ���E��yN"�~�(ͯs �.Tq���I��uE��C��z<�X䀺���Z�S������=���1v��Kqdo���u�. 著 �E�b�G �4	��qBg��qP��0���B�Ӛ�������:�nW���{�p�3o�v������%i��q��� ���kLt���g�)����rY��Z�%�|I�d
w��s�p*�˖q�Yq}�OX� /��0T&���=��_�F����?<�Z.�yd!x�d7+�[D����<�y�U@�K�{���1�"}�M�0���E�S�.Y�w8��r3�� Q��m%S��,T�f��ON.�L�K���a7�-�����C����Ye��U)|g�Ⱦ�1����n�J×W��ta�S���ɛ���`]Vò1'��6�z&&8��S�ȧ|QH͎��isգL*1�{D�j���y罤����a}�c��l7_=y�S����ש��[���"q��^n0�O�N�W�K��R.��Z�	��Cg�r1����������URR���$dbG��H�ʉ'�(3 ���+y���
6�W�U�i�<��A���g���U�s��G������[��*�j�r���{�&�6�9�g�.@rK�� ��5/Ɣ�o_�2�t��<u���P6����&���{���:�x75�g)M��`�*�W��b�ӆd�x$@2�mه��{�����X���s«ǧ�ڍ�X2梌�d����T���fq�qDT72�L?�p�D������/T��'���������1vc��s�/����!�-PL)�H��}߃p�c��,b��JB�H%?8/���U. ]���dƏ�R#�mJ|����{x(ňǥ	V��W`fv�ʊEn[{SHy%���ϩϵ7[m� �V� D��\���Z���3o�Q!CYyy�R~9K��{�X�\eX��i����>iv|��	�{�����5�˻�t����17ق��D��3�����h��x��\�{^�ʄ^�_ש�L��N��-�}�9�F����W�;�d��A9E�`��TZ��`G��wЃ���+��5�k��q�2�Ћ{�4�甲�����кZ��^b%��I���}?�d���l5TT�c�vgX��{L''�솏�jƺ�D;�I5-��S�F����^;u����w�f�.,����4h�����o,w�#�os#���}���ѫҾ}
�Q�������o{;�9����gt������3���G�\���.'����W�k�������L?8�7)��ĐM��̀�����|��bJG��A�)wP%��b�Eۇ�A�?ʒ��!�� q����fw�1	�U̠I�7N�+��6��9����DWW���u��Z_���n<��'9 ���|��*��3���۟ˀ��0#���ض;�Zp��T�����K�q[�xyq��'l��b�"��ؕ퐬i�o���)k�KQy�o�Ǵ���FRE����!ל�e��i�0�;k�B�D]X(S;M���-l8f	���(�bH_:i{�"����1O$���#BqL���Q}��\YŃ$ӳ��+3�J>x���C�fY��/����5fK�rw_�����g����Õ)��̮�v߾�o�=�6� ��N�ӻQ�E���lh�f�Ei��K2-�-Aپ�=Wꋦ?Xn6$b�	��L$D~,;��K��[4�Y�_�_���E@ U^�N�#��7���r�<�A#��ע��7��Xµ�F�\fB	���5'3\�IЖ ����&��	cK���
�J���c���8�Ƞ+}w4�q̵?��i�'�W�E���]΋<�T�fx�C�s���I���x��9���o7>�?Ϡ�F���\�͋quu\�����a8劂"����Qa��� H�����w�U��a'X��slnn�7�������$Ȅ��� @/�֑@�孖z���e/��M9�L.�+����髻�=��Yy�U��qQ���7*�x!C��@�JѼz���`4�g�c]�`�	��H��ج%Gۮ5����锌�X;��� �?+X�3 ��o��8�W�[��Hv�rao�A4'T�����/K.�N�J:���1R����<ׇB��-����Wv=3>��IfGąM�>y��2&�G��;!qt��<(}8����d?���O�l\����ͧ$����k��H�'C=�\R]��B �B q%y�.i����*ѱh4�q(���F+��6�Y�zڊ-o��_��ӏw��܇��>,K��H@��,/�b�/�B�N+W�V3\��>�}�z��m���~�>o�wp�e-��IMdܼ��Zw��پ�)+�Vw�ap[KKK3[N��ͺ���~�� ��|�2�~[r�����Q 0^�Fؼ�8a�-YS���L	�.Z�fb���ٯd��!c��Dا�^8��%���WEϐ�4�vއ}ɏ.�5�O����r��qa A�hq?KI����|�9R��"�{�~<<Kw9���JO�����P'O��Ҵ�Z��g.����#@���õ��N���ք��e�<��e�$LEn�B�Z����a��i��㩎�.�,%�H���m��F?�ᒝ�s��+����4K=�Nbo�`P��1kt���ܒ������浪�K}���0Tܳ�"���OI��Ն'	�Y�	R��� {/���8��p9n����H�2��IsVY�GG�{B_of�a�x���~���7��u��MB7�F�A#������+S~g�π�S �(dݹ�m~-����98JX[��rz�^:+�����9��R�E��M��S�,8k�XTh���}čf�A���L�_,
�	�sO/���z��;\6����Q�ө��x�WLх�,A��3�-�z=��Ⱦw���N˂�̎s���m��6��b�'=�d��ϪuSr�[Y���1�P�!a�}8nW����Ǝ�����C� Fl��

j�ꅭ�E�|��)[�����1�S�&���pZ�;&b��w
jڍ��a��|h
��pg�M�A=.fr��DA8��y~e��~�;Ta�o�7�@;3����F�g�=�'.:A�{g�]k; �������Ԏ�Ito��qv��v�MI�Z]ٗ3�~Z�(u��E���C�x'X��9�փ����ؿn�
59U�]5�{���� �����0s�uY���|A@�-_�w�M�$J�9�!Oz֦ 6jo�.�7�^��7�z" 3��$�O��p�'���<�g�Y�sW�bH���;��f�Ɓ�y�.��۟?�F�q HS$��������r�p��H�ο@���������m<K-�K,Bµ<c�&�4Ƥ;dO� V+J�ց��ms���~-,�$YdB }fE.i�;�����8�(�P���O@U��R�B=9'��q榝nV}�rS��a�Ya�����t3�e�PW2��E�/ "B�# �q?Ly˙�b��0��sym6�H�_3 �J�y���/(��!4�~u^��*�uTj��t�oZ9��y,C[�J�"��H�<�n���ݔ�Xd�"���jW��fLêb!{RVVt�ʹ�YY$�L<�+��pU7�'����Ԗ�;!�y>�P0���aHhJ����r���}�����\�Vn0�����y�$�ZXߓrp�P1#(��@��M�!C�;��|B�&�f>w��G�����8�=�]���#�	�s���I����������AKݷ�; %�o�ҏ��Ȇ��ր�-gU�x��e�lo���_�ek
1rk�f���66J��� V�5�u�	���G|��q��3�jF1��`�_!U��_�1��}�5��4\�QO+��	`�FZ	n`��
���^q�?�=��?��,ָ�!�OD]���6&cUf�óZ˗]��Ţ#F���c�����B\�S5�[
֦���m���gb�5:�������d�sؓ�3���	�aLM-�Bsw\/o�
����>u"�7�3 �(���HP}ڼ��C��U@���J�df'�?�9=^��ot�;�c�3���W��`������A��l$j���0�C=���@da�|��y��b���d=�e��%8��j{��-���ܩgGP]V���`�2iIz��I�E^(H)I�����>��ܬ�<�ʔ���1#�9|�ڋ�����|M�H�\��x���UiL���*ع^�c֒T8�vvv�-�8H�`��7&�Rƣ
e[66hŗ=��9����z�Ym��7'���e��>�3���X��@9XBL��Z��_���!�"��b�%�R�1��75� ���[�����޳!S�lKX
c�[�����~L\=G�c�6�˟�=�=-f�5��81���p����x�I�ƚW|{����h�@����>��������F�xh)�A̖9_�q�2�SG-!�����o��$�Sm��:�z���n�#P��K�����V��<B����-� ��_p�$+���s�%*O&$%�b`a��k�|WWta�M�M��M��l���f�[�d�l�k5m('�z��5�u��i��N��)�����3��m�+�e"����}��Q�w�˴AE�+�lγZ.�Y���n;�.Ǐ_�v�"�7��_��_-@!�32�M�X9�Xi_q�Νs��q���k����
�pIG��&��Kz�k��_�D&W��(L���^%��ZY5/*�b��Z�q��sx��i�ȼF8{~к]e�*�WH�0te��v�l&]�ɖL���Dl�&᠅���P���P@�uÓ=����J�Ⱦ��RF}�[,�d>X��ri�,�퟈
�u��Q�5��E��ȳ�*�����u}��M�J]�y����Ȫu�f�r<4b���;��"#jr-Smb
�Jr�NЏ
mqL�x�*��!D [�x*Gb�KHN ��]_Qo�x*~P���p6��=+YR�.�����}��g�SZD�h�ʎm��J����C��u�k������o�)N�RX'��s��U��� E�T���g<\2�2.�HS1	CE��^���j����q��Me�w)��1�6٘�G����`�z�6�E���טc�$_�偀:."��@x��祎��l��sJ�z��y���H����1�hF1��*�i,�iÆ��%<�{�\P��Kd/�sÌVj�����IŇ�g@���c]v�8�g����sq*Sݽ ��B�e[����<����4�[�a�=)k�x���m����$�	�*Yv�
���&��Ʒ3�S�����U��W�
fa
5�.A9��Jo��k�%�tF���.�!��[���#
�n6*��ݦ\�r����%�]�3�2��9�7��8�ܭne�Š��l�RN����wƬ��Z"1��~�8���u�1;W�bO�!`&���H N3ZF@�W�Vi����/;N~����u{tw��8�V6`k6�1f]t~^���h�t;�yc�խ��F�w��S#��b���!�)
�G���x�qI���qNj����Ќ�����ɰ�����x̔$�=B��籉신C/Y�$�ms@zZ�GX����#����j3�@6b�үsE)�H��Sܗ�7�HQ�@���tacxr���bb4�_�ighV�{�h��̜���|�l�;lT2���߇��)3���t��;��v�<1&[�/���o��/Ss��!��7T5�'CD���� ��)��_v�%��p�F����A�_����
` au�'��+�eR�Z��	����+�̂~�f
c�|��Bz
6N�tz*¾tb.g!�A�`�����v��t��|��P�l@Py�}�؍�1��A�*]� 4m���m�Rg0Q*�bU��+�Y�)��>�H/ɛ�D򮀨n1�<�U�*u����a��B�/�$yN�`��_��<�kv����W7"���ty6\�!���)g��*��i��	C�3���c4��	w�Ӭ�u Hd�#CFBR51�fc�����k�5fK�xh]W�0��2m�.����s2_�t��!��T&X�W����|��Vv��yH4�$Ձ��0���Y}vk4rl����kpzr�Kj(���R��
�䪊	,]� m(!��R�?�"x2SiQC�Tm��D�:���f�8��U,�G�Y�Z��Hk7S%c
Hv��~T|���a�\�;�y���`�����X)����P���7b6���Ƣ���RjR���)"i�\7�p�㌤]����\]^~-+��Y��׷�^\Ye'8�h���?TO� �,Z�{����B&tCI�G�)�������0�~~Uo�g���$��� ����7�vР�Nw�r(�a���/�M�3�udQ� �gt�nd�A�<���BJnM.`U�aN��\�B9)�VCMsq����	Q� c@�:�Ş�X�D��R�L��or�愭���G5Ú|�����`2��zm�xB>����,^eJ�l�D3u���_�Xw!
�ǫ�o�A���ػ��3�'g=;��� ��Q4��x����'d��{5������5�P�@�4'�M����?M���&"�a_�QBN;�o�D�/gؓ�_�Nn��F�O^U�Q�^fM��&5�,n�p����^�0���2f]&q�o^[�����6# �>���sHA���u�Y���Y�Ȗ�Q��N�c�����|�Wk��я��l���y���i2յZ�'!����UE�L�ɤY����!n��.3v�Z	�n$��ޟ-\3�$--�@�j��ZH�V��)k`�|�7��;7��Z��̩��~pT�������%v�|��'�����}��3o�OZ E��������qT�׾6h�Cc5s
G>�[�F��j�*��Q�~�p
ظy(��-KC������[x��]E��ʇx�km
�{�H�n��L�_�4_6����$M5�P?ꖠlF���캬�}�+EB�}{Ǝ8w�������g)�$�w8��sk��A+���3�M�ح	�.V�,��@��_�2w l���e���<���ޘ����w�E�Xya,	z��dCF8ac� A����$�p��ۙ��\�[8Tr����%l�x@@炙�Y�"`��(җF�W��t=�QŘ�ոS����-~���;�a
Q�����Ud�>M���l!����Q����X}c��4в��业NP@�7Kn�i�5m	��e�G^v`2�u>�s�/�$�����/ll4�>{zr�=��������7b���@䞞ʿ�Ǧ-ѓczF�vJ��V���6��� �O����63V�m��d��]��"��#L1!zy��g)��b�(!�<���cx���z�9���K~�vry��s�ʑ�3�ר��h$�B��tڌ�R=Z�h�7\��\�����L9ߤ�87%2�Kܸ��w���J��HS��?��9�V��)W�t����(�����?���V��M��L����$�+Ap���@�2�_	��� ΄�	��d����`2�$J��Ќ�~�����V�-�Ɛ2����Sk~N��Z���| ���zѭ˙�h�!��-����~%�$���3{����	Bco�����jr?ݵ�nI�T���o[{{���ZJr"<������K��XB��#?���g��Bf��@[j)��^�{��N�I�v�@K�T���|� Ə�,�s�%�Z�/PS���`E^���V^^^G�fo=	{�m1����83�O�����N��f��ֱP���r	���B��-�����[5��ʻ^���$�c� �jDt����܅��r{�1���_ϭãJ{{{�!7�6a����Xd�ge-�^�O���¼�^��l�d*�^��.;y��^��ڮ�Z�cX���I�Q"��2(����V���*~��Ay4��c���M�R|���������4t�߁H�������Gמ)�i�t�!C������U�E2E�Ƀ��(7����w�f���jER�Q���� �u�V݄ћ��^Ry���f��6���$��]5s�@L3��Kl�\� """�{p0�;%���� �j��u�����&C����#"������N�c� �RMM�ͧG��T�;���N8�d�7LL���RV�xt�KDEɴ��(FE)/'�Uʦ�}�1�T\��u����E�=�k��*�~�,*)������t��*���b�HH�gd_����^���綶�����.��u���#���-��#��u�6w;�����Cj-��?��1�Q)?�t�~#�FT�ZL|�� �u��(4�H<�W�o
$�U9 ���x(,��g"A.�s�sp�߆eT��m�X�u�m��
�8�_�E�<8`�)?��9z���a��2�o�6Y%�67�׸e�M��"c��se�0�L���m���khh�����&'M��I���������ٽw�w�(���emZ�.�厲��y�ä�7)�#�697gs�%�$99���_�]NP ��2�v�9#�����Wۣv�^���w��w�D_�Po�s`�5(���O����)(A�����fp^O��y���5�g4笁�%�v���x8�F%[��5B���ӝ!{�����	R>q�5]�$[��`���'
5�
%��ř'��&�f(��Xb��OV���rn�.�e��r�@d����\�7�n����W�\��b�����am9�q�r����E]Sn?.���̬�z�<^s��3��O�ȶ��v%��ϳ��\JZ3'p��q�^���p�&;J�(h�#��S�� �S�6����t���DL�FR�~��AMK+�*��߳p�Lמ� ��`����{*����Y���
�9��߼�I�Y�4j>�X^_��ۗSڪ���ޙ����a��æ��w�6#>>*B�]#��h��>�ɇLŘ|	�bB��uy���b�5C�]��jM�9%�R�0I�S]	Y��녑I� DӦD�2���F�݂H�>L���E�֝�z�n��(p�3�|��ʚ::�,A�@y�y�A7-FD'�_�`Q������Uή�X8��⢭��u����~�G�5�Q���P��*1��K�]i�?
u���HW�!Ǖ{�X�-r	�z��g/ںQ�%P"�|NXt��l�~[֭���S��f���s�O������w�K�I�֡�&hDi2i����@���`��E I}X0��lbʶ�o�<*��c�s��{��8����ܭ3�D��������9�_rx�k��Q������ ������󴀗$�~���;�&���X��X���2JJJ��*�����=:F`�ˍm�h@��ͅ�BW؈��/�G�L\�{��� vn���IG���9��_�-�662q$�7�@��l
wL+�{��d �f�f.B�'�����v:c����5�1�i�D��-c���߉��㹫m|q)�V3bRO�1��mj՚��q����|�t��`,qiU���[��+JF��ڙ����-z����eq*����'�b�N7�[��?�1��IT�X�sm&D���	�4���o, [c\��#vc1Gý�D��4�TB���9����X ��ڜ]d���7�?{�j��7WW�L*��WA^2��#7���Å��NL�@Y�{2nh�(p��4�f����Xv���/��.M��(lʹ��	���ZZZJ4?�7�5�t`�47i��ivs�0��ahu������bu�j5���
w�y;V��?$��~,iR���%�G�����W���C���(`2,�ClwZ�`���(��5� ~���۹��XN�r<�|��s�jO�%�w��:jR]��d��㐔�K)d�9h{F͊�|�bd��尔0�j��ߝW��*�mFdkk��79������H[Y���[�^�%'������H�tO������AbYYY�� �*�
����}�}o�p}����v����9<�Ӂ�}�`��ǟd7f=Rշ���|w�-/|��ok��s7 �(��IK�sq*U[;	����h֘
 �v����Vـ��l?�� �!�H�=����q���>"�k�u!�f�:Z�!��G�t}�ߍ���Ņz����CN�8�X��) ���F�LEk�n�f�wjx����!��'La�x9r:����tЋ���u��gԫFK�u��gVi�Z��1䖸Q�ɼ���4VI�M{}�h�]�w��C>��j���ٞ�p�Fi���x�Pf� p?�l�@��U$��&(�␆#�|�))F,%:&T������@�5�0�f}�ɳ~����\QWW��}���#s��}���Iv�p{ឤ�*Ů��_%J�ϟ�I�^5��;R]�Y���*C�cI���^M���=M6��`�)�w���,Ğ�Nm{�!	��� �cY���wu����MOO�]���L..�if�TG���TF��?��R�y�l���f�[�zF+�S',�K�_��3�<�'��ɜ��x�0tz�}������HI&���x"�^�X�۰^���-�`�r�ۏa������l���dXȽfnb�o�C ��ˣ ��;���o�2J�!�\��8]�#O�ܐ�-��qUn�d��\�c�m܆�(��I^�2|�{�(@����Qƞ]���������끍�e-$$!�.�\{7O����0P��҈�,G$�ScWWW@����v�w��W�hz�5��A�zY%�l }��ր�#h��&�w��M�fkmhTT�P��T�8�SE�!�����dd�lR;��!'��[�3�[�d�zܞ;	�f����{{���_����������x��$�@��}d,�F��R!�c8uơ�:-4��0��@���<�s9H|*�r=1Bk	�%��4 g��k�F���qe����_X��/���l��ǲ�gd&)���Rk�4��� �(Ķj|���0^��L $��i��!�^�'�[G�o)���m�4��}y~�N��K��_�Xȕ@&y0���T�f�?Q�`EZ�"���Ew��\�>�m�P�q0[H�]�>!gDej=�n��hє�8?�d�~��3�����#���Wرu������x����N%�\//~XG����;���8��U{�R%� J�;�b�̐l�6T!�CF3��?�G`gl�ʇg� [5�r��h�U|4�������\U5���u;�9��s>���hhr?Y�,���*��v�&���	E������6M�' �a3��#��$Z^x������؉�$k���fg����\�-�5���;��vp�(r\��ǈW�^���dFL�W�I3�bv
 � ��h��!)��G���wJ��|�b�S	���h�y�PC%�3�''�wRR���>��44vY�X���ΨG�rl<�Z���;7!|�9޼�����TɆ)�c�<-�	�D�.�-�:M�2�u��If���
jx`�����/w>�+�a�> ���VM�=v�4V/�ն�E	���R��|O(@�fh���]	Ywٜ6�3Ȝ��(���N��Ao�|��8���65��� ����Rǈ������t�y8j꽕�sz��|�g��ʤ>܍F�,�5sSY%	�T���}&�1���`;@�uX� *���
멽h[�<I�sˊ���-	��)��~�$Y�[��S�%!*bqR4j��g[|�4��:,�sg ֺ�]��t�3�t���xx
v	`�B��tt�+Xܔ��i�'�^��!��č.�@8(9�D��1Z��	??!
����33z�S�a8��}�]�zF�_����~�*�H�*��l�HS���57�-������j�H�5@YT������{먨�/|x 	%	I锐nABRi�[�aPZ:)	A�����������{����53K�b�=w�}��<��{����F*�!=V�P��k ��H�xN���d����^�I0^M��Q�?��vp��I�h�=���S�,��Cz ��V����5?����4���&P���H���Dް7_� Sg��IԻZ���{d��%[O�w���� �~\};h�����oI��:�|�R�߯�!��p̸��Y��M]��jx˭�"��.��;¬ϹY�ԟ�+�s����=^��"^�lHx6�֟���������a�*�I����h��lCI	���!�V�����;��_�/�	AE'�{Thb/�A�۷�{:3�������je#��aZ?�pA�z��װ�v��х���P�N�R�!X0v�ρ���/F ��� ���O��n�3�]�at��sy�u�b���{݋�=��p+#�ՠ��~њ.HP�\@-T�k��Q���tvl��nn6Wc׫h�-�K�|a��y������Տ��\�B��G:e�.�Ϯ�4p'�\.�Q;Kf|�Vν�o�zG?�;42r���b=�c�-����;!�b5�І���rbb"�4�O�@�����k ��r�`��N.e=Ű�!��.�h�4�MƑ�
�{���
�F:��ེ�I�R��ȗE+���M}�C��C�@=�leY������}��_��� �`���u~��0�wL�"�8X!�P@������Ww�QQQ����/�BՊ~��s=���$�P�.A5<,@��oB�]Wdg���^�6������pdGiZm휒���*�w�P���k��i�g��&������$��y�:��͡}D1}�ܭp43S�홝�|����)�3��_5ӆ�L �3�1 � �`x����i�`n@[nS6�ғ�fx��x�o) �
��S �*�n���{TQ�����#+Z��C�U �+Q����XGGG~	�۹�wy��z� ������"&ȧ��Hl�q᪝gEW:��HՊ���o����cKK�����7�D1w[�W--kՇh��mN0K��4Dg����^FM��t^a!���ݸ<���1U�l��E��{!�B@. 96�)��ykH�)��!�5k�;E������ZYKKF���tw�M�TnY���Zo����t�@���|$*��������H�Ɨsg/��>�:���*�"C}V"�����O�MB�ޮ�JWR���'WĲN�y�S�x��c�F��ڔ/(D�ּ�q���}����{h����Y�����x�{��CB'�d&��q��(������14 qF�~2����e��.�}z�u�;=g�12�ǜ�]����8�X�p�`ߌP�� �% �TY t���؟Q<Y���ap�
t��U ��π�G��ض����v��m[�zc�������'�����G����s���`=j�ҽ7A�J�����aN51vQ�Ȇ�e��R������y��`���r���̈́́��.��F������i-GA��A/���S}Y3��r��W9� }�ҥ��'m=q������@w��MC[#���L����|5t��i\���SH�#H$bb�߱	x�w���X?3vC�*����ՠ����y�Ųz�N299���2��(�M,o6��g�[�ia ����%8ZEg:3[@������߷G��nB��XF��Y�H����p�=�ޕ#��"���M@PM��� ak ��7��Y�[�͟Nz�ϑ��C��M��ڕ�K&5��0�Ĉp��\���'�����_!\�{�{�w��P����A�н���psԦ�)ʀR5 ��FO�c#ܩԛo Z��orF��Bk��n>�k�q&�=�W�<�S���%b�u"xcۼ_'I���.x7b����h+?,zLĶE*����h� �5��{ۛ�ב��Z]�鯚!Q�#oEO҆���k���ܞ*8h�5"�90q�P
g5�q�K&����u�8�%%f�%��6�P��1�4��Z��i�WrEɡ���������,o\-��\c�d^��ਯ4`����^�Og�Y�8w�r˲n,`L��l������ʋL���A�%��2���Q�,˅�$�����뭧�zJW|�Q���
*4t?�}nl�)�B�cQHZx�F��vp\����n�J��b���j����u��qT��6� �iA&��Ոۧ�5��X��"��|�z�b�]�����g}�X������Y����>� �vp���A���P"��z�����{m$���O������^�t�����$�n�����/`zY��`��Q��H:}��:?1?c)+/@$O1/���&� �;{,��N �.��%v��t�����ȐʛΑ�nLy�m�&�,����T�;�>}_I{������5�ݰ9t�;���0Zw��������0ou�O��{o��`Ā��P�Ǥ�^7� Λ���-~����=��S���[����T�z�+p!t�tn>�hM^��nF�yK��j/��
P		��Pc��������.q�y��!?�I-Oz�V�5YGFCy��r�ϑ�ė�x'�C��P`q�>�[���N5��y��D����֯�dw� lOcS���R 8uQ�����Xf�5*�	�(�y�<A�v܉}ʏez��������@7U^�;��<9��O�}�W_�?켍-���_q>������iH�CO�Y�iS�c����q;V/�d�G�޼��Cx�q��+Y�/x���9^6�;(��#,lx���^D��� �vC>�
�,~�2�3�B͔�@��|5f}��ig��q u�����H�Y�eu99M��wjj��>�{������}1�k0ȭ`Eۡ2�r�&��=��M�lQM
Θ,ʱ9fݫ������;0ȇ��+�K�R�vI�lhM��Dw�h�z�9E�z��"�$3�1�Ⱥ�g��x82$J�˯�C�ñz�o{�VhL�N9����+�s<�������N�N'_�w~�_b��:4��4���f
��i��W���v�rnV=߂��e�B����\j��1��W����4�A��a����J���6�g�WZ��?&�az5s~ޘSb?[Η�����5����P�w��,�m ����2Yp���S�%�}	Q����g�Q9555�u�]�w���*���qp�oE���|���6[b���g��j(]���� �^e��v��y���E���`���+F��!�%R��	�b��h]� A�d�R��:��x�V��D�ڎʸz�r���5X���Cgl�T>���e��HSq�3�ϑ�8�i�o�"������ۿW*����� }\=��3d?���ʺ{9�v�"V��Q� ���ͼY.O[�"���oBN5-�~���èzxn.��郜���hz��hR�jLT�>�}p�^U��m�+�Z-w��c��s�n�,�� (�8�G� ��g�W�Oϧ
��Q������a!?^T������d�{4F�����$E?j.�@/��"z`��v���&���?a[�]9@2�z��*''�����s�^hW�~s��K����g���@@�5s��N�Xy|��ĩ�����#K�b��W�w����q�ʬ�񳈝�9C*�t7z׿�y�%.�$�~����^�s��(P�i�p�w�p�g`�/f��q	��G�����[\^G���n@B|G_R�5�:�������ʍ.��%�!��g����[�����!
*{�/r��>�q?���|�h�Џn�����e��������!�P9�V �G���R;�T6a��ۍ* �|�\vv��W�u�b}3�:C<�ִr�nY=y��[\�}ˎK`�ׯd�Ã0g������ȟ�����Bt�i�%�Q���c	,�A�{�7.��{jZՕ
�vLI!g�_�:o�n_��$���#�4 ��;�}�M7ċ�kQ�&k��|���F&i+�0�]�(d�?lldu���T��_[�k{l+����{t���F�խD$Z/l�o��\�s�b�, �i-��qA@H�b0�Y��}��T|��$m=޻����H�x ��8
���;�E��xେ�_���#���;c�9J�ǥ�4ڱ-�=��O���V�E����8�0v�@��-ln.<K r���S��r_��}���p�:n|�+��ϟ��ڼaPhHc��Y�|X���if�7ca��	�MZ�&m�љ�դ���5���xK�L�n�֎���,p!���R��%k����$5��U���D�I5{l�VTd��P% �^��Z��kn�%��D��> `+��=fK �::�E]�Q��r���m�s0����N~����ƪ,Y����a%v�B��\�u�gAf��<���(k�PL�J��Ih��Nd��}��<�ez$bu�hh��T�Ɏb�kn��M�S�̴ɱ��p���#�m��&=9B ���R,!�L��:�i��/��5��=az��]����W��O7�:u����,���2E�k��Dy����ՠܿ��E�V.�((��pȱY�::Ə��!Kw��3P����<y��[=� ���nϥIJU4���b������k�۳GY.�_�NXC����xn�r�Y���}�$�����)����t�{HO�I@��Y�[!X`�����y���m٥�խ7�n��34���QP5nwe�3�]����j<l��w�B"&v�6.�_���ld�*�[W_o>Wc�s8�:9�n�VyAr}KEe=j�=���������v'�-@29��J������'iལ���8L�\F�މ�Kȕ�p>xBj6Ό��,_e����1(�H|�*>�?W$��u������C��RAWߔ��\Q�K+y�Ԩ�D�!�2ҋƹ�QK�t�s^�~�+� �xn4��XR�Y�#J>W�V�mG�����:�c/��Ud,H5�8ۨM>�I3$��5GF�t<@�����2�ˉV�4��@��(�s`1�)J�K�-��ի���@(�$E�~:��IT̠�>=�ګ���E�Ac������aG�9E�BޫE���Ӷq�Dj��&z�Y&�Aq.�	��y��v`C����|~��Ğux��w�
/��}�zf�m ���2V~�X�ZS�Cx������4(�|��A�,U®0"z�5�ZAxW!�e��Y��߯���?�W��.�.HG��=�����Y�5E|�����ӷvj�q���ƳV��5���MʀU�y�������a��F�ț�̻��1zP0۶��L�ZF�:B�ŵyBf��� g�զ2gx�q��t�ԋ��#S�Y��
(��A�n\)��hˏ�71��1� ��E�.�j}G �p�t��V�|��>�9--{���W�+�Z�B�`����X~2F���>�lqjeQ(����椈+Fp��i���� 9��4��-�M�B�Y����l������d����Hʛ�b�eCj�M�+c��ʺ� �7hX=���Z���ǋ�DUf@��R�+׻O�TB��qO��� /-AC�A���^�9'EF���f�*��'TWS���k�,���״���[��6���;񡮧���Qm���I:+��i�Z�zA��L���x�,}x�����G�:Y��z���^pO��ӯ�`���L!���z������O�U�+�+D����1,U�PE��殰� /���x����d
P�f�oC�i�W��0������f���[T�/�؄8�'��OL�0��+T0�0|k�Ӿ�	}��Nof�UO�Ǐ�	��o�}?x���CCL�<��})��:~e�f�q��~z��\�U����� ߙ�j� t�@<8�R�v�a-<ؼ�]�������}��4�e>�|��l#�A�4aZ���2�𜭖89�]�9J{�@���S�a^�T��z�n��vl� FO���o����vE�������u�}	ьH�
'l�����(���H���;^�o�e~��g����/)���O��� J��1�oFa;���3�s=��F�5(�9w)��uJJJ^�U���Ѧ���4����6�R�F҇+o����Oٕ�����\h>	�g��MR�/&Q�\H�B��0s,D������||���e����'�2�r@��� %%��Dr�x�x�=����}4�/EG.�ع��*�TJB�r�������V�s_��'?��oL$h#�����PQQ��-eF��M҂�o��;u���s¦g�PS��O[�	c�H������;<��z��B�����a1�-����� .��N���,�����Z�/QY��m��3��J(*7�w�\���9|�!]�?;%��_y�h�aω�@���ֻ̀wQ��4'��"z4\gQ[.��6����t�'�����_�f~<|�o��jW_��j�TŎ/�3���DGOӽ&�q�٦?b`��\H\C�t\�N�i���ǿ�e�"8'�fè��V���O�t�؃
��]rٖ4�lu+�����H�ib^ǳ�Qw�a���}f��C��K�M�r��E"j��3��U��AO�����8h��2	K]����&~B&v���͵�v�#˸�+���L3�J��N�~���]��K��ɧ\�	�����uYyyy�ָ0"L:F�ۗ�c闛2��b��isq�o,\a{Kңk�3���sr�7d���if���Y@d�{��� >_���-#�������Z��5:��HgZ�>{��ؚ@�fKe�}��G!t�ڗ}=�0��~.�:�ށ}<�����y��3������L9���V �W<?��nXt�m� ����B�m�fM�͋}�� ��h�^8��[_�ư���9l����b�d�Ӵ��<$%{��Ē)��L�YK�d c�:��8�����c3b���&�.-�����������E���\82�M��B��ѕA�j�{\�u��'h���|�|��m>�)��?N@��0s���������T��ٱ�}�yA����`%�~��@��<�[DFFݿ���U_�r��bŕ�����r���a�U��y����b��'O��������G[{:{yC������!����ª�]���+������Պl�Rj��^�Y  W�7�ö{f�F9�@�'�"��lM�W7�"� c�aqRB����\giq�6��E� �X�k�/�v73y���ߒ��N�|$*��߂�A�bc&;6�� ���n�K��-��C� E5�G 1,Tt�E���%�8����Lu�&ΏR�Yy-4�5�5�2�B���PpN���%V�󰿈�����RK�1ok�L���%��ܕ�0Rz��x�{����ɻ��1��O9fܩ���%/M}����pؗ���݂ksD�§�ĥ˩T!�"���dq�l��jq>Sg� T�+L��ʯ#фT��Y���3�v<�ҳ���;��$h@[��ڋ��� TMrr96��K��w�'��D�H�zUK�&j7�B��� 
�i��n���.m �Iu�.�j�mR�q�3�l���u`T��/��4�l"Fܥ��]����L��AZ��!�bƮ�i#Doՠ��"�T��%�������Ŝ<�aH���fMRi���|�A̶7be���Ը���+8���wg�J�?[D�_��Z� �����IՄ�8�*z�U����K���e#�e#�&���Oq��ƾ�8F�xa�&�N��=1�^a4#��;������.�Q�5=�̷�ٷ�g�{"g�oMUEǀ��N:��}�z�PH�¶֯��2>���W˴�� ����N� =��Ϊ�SߗcP�C�Z:����1�ᮊ S=ul�C���Il�%�w�x��8k\i8t����ԙ2Dƽ/G�,��=�6�/�?�:̡3" MM�H1�	o�A'GG9cc���i��t";P 澊��`x��}�"�=�9�����QV�r�.���K�Fa�/���p��/�Z��ɳ����Z���6���[�2��nǾ���V˾��lw�*�����&��oF�/#�K�(}.��j	ZB	��N糄�$�d�� � �������w\
�%U-�h�Ek��"��Ex.��YA���T�E�t< �wi"�vz#�w�˯Z�c��'̼Dm�x
�-�T��'����s��e|�D<W��l�(�L.�گ�L�44�B-l�,x��A��!9?7�6/����d���N^�L:4��Bu�3ŷ�/�4�.g��m����Ϻ�x7%%��;�d�'\%��o���g˙�\P}��y�($e;��`r��&%��
�kh ���Íx5��g.hӀ�iyCŔ� ���Ǥ,�%[�j�B�&�NK�v�G�Fv ��ߑ�z�I�/�p7O0u?�?\�󣒳���[��e�쭆���CE�yKe5�J*�7t~�L��<d�^��@��^��L���D�; na&�@�R~"�u�O�eۿ��YQ!���pTKU!�(+��i�_/��5պ���s����'vN���v�.XaE�5�{?%�1��H"̼�����'-�n��Фy`��!T�3C�-�5*��q&���XuK�&��qw�����g���C�{?�څ�����{S $8wč�?�m�yvH�.��Dk�N4m�M:N�pK���+�����^��,�VD��v�v&⇀v���( u|#d|����c3~�V�~��� ��e��#��=ĤQT�h�n�9�L�����E-����ܡ�>fA"�fN�_�e|��4}B���޲ l֠��1�n������TM���Rm��H�-.�P���r\h�۳4je�:` X�z%��g�u���ȡ
��nn�����1��%���Om�$$=8x���H5==�&�*6�1�ˆ� �gqq�Ҟ���?>�4�xS��F݄h����5)־c@�/�=L�W�����~��(�)�[CCq����H�G�%%b�����UY��?�A�?�H���{�8{\N��T���@\,����v������~�z������5]
��8�V�(a�K�7d#*���#%T��=&P�[����Yn�x��4����C>gGA?)aϛs�o	��'���gx�ζ�*-������Z�A�l�J8h�Ø�0��h�/ARٕ��bY
�������s_|u�'�]9@���ƈǱ%�;�E��e�y8��!�#M?n2�Ę
�w�s��6򉗺dr��ڪ~�ڏNv/RiȎEdd�2�ְ�v��J�cGjo��۰�˂Hʹ˞t���xw�����*Vڻ�ۤ�k�`V�:_,U���u���Z�	���w���T����J�x�z�o�Ռp��ѡ�& /���Y	Z�C=)�!�-��+�<A��^�a斓&>F��<��Q�zQ�AY���Jj9:8R�ʇfg^&l����k;io~��qWrK9�5�o�����������ዋSg<�Fe#�o(���X)i�QP ��ݹ_�JQ#za���u�������F��kV(6�H���:��]W������5�@x$L�����ug�%i���l�[J3$����k�K�i���`��1��s�~�x�������
]�	�)�u�7{�.��i1��[ިN!�ȅ�N�w�{Vb�ڌX&�+69z<S����_�ь��9r�\d#�?/j�v:�_c�`MN1�5�'����!z�i��j�~ /�A����o����wx�E9���t�r�q�S쾳���3[M�hqR�4�a�29cEr�uF��B��JG[[�m<#�g2I3�ڥ�bA�k���-�^�v��OM��&|/8�C�+a1f��S6kU�1��em��z��:*����w��,w)��S�mn�n~k���� Tt���h�M��:1?��w��� Ze����0[L�2�L�b�J�^�y�.h $A���Z�Ĕ����ù� ����XC��_^@)��%ϖ��Ի��%,��B^�w��^L���K wM&�y,K�p%�Ë���AFt�K4y��Gx="�*�ٙ��ퟅVy� %�j7s��H~3K t�3�@_��_x�j��{����M���Do�Ʈī/�Gm%�s�?P��6�ŕB�*\���/��/;��혪)eI�OR����'�����n+Ђ��
 8�4�.0���>��Ѩ���θ��q��,� �}�S�pd}.,5(����d�e�P�{����
��'A�
����Ѡ�ݷ�￤�uuH!w7{�f]�d t��oC.F]���m�$��$M��y��閻�_�U��>� �А�[V�a)��ʕ���qݼxï�*�
6x�dq��������4�iS�R#	�@Fڝ�8mgs��ה����j�c$o$��έ;U���۳��.�7�7j��dQh ]1*A^*�����
� ���&����*.���Qǹ����1rڈ͟����OQ�0��2|�y�������e*Q�I��:@������<X�)��%��q��p*��o�F���`"�:eC��]F���Y�����1,�~q%���� �+fp%̷�g�<Ü��&,��E��7�l���B$F��[5��0Ԡ9ȏ�mHd;�:����r3{�;+�}��2v�����鑷�D72B,& �`�-)i�`�ab���}�(������8蚋��{�~=�,���|��߼״j�k���3�_������"yI��/Ӛ�q��p���̊@]z�/�7��&��^�\=8W���r-Q�]@U.oR$�v��8��4Es���*o�;ECE����͂�q �~�nc�)��!������#Hp��}xpH��/�1IMK2Zm��'A\�署��;4���j��=�N�y;�.)	Ѓ�=U��J`i	�10WmU���B��B}$���wء�DY��Ϯ�൸��=��Ü�7�C�F,��/q��j�����D݇��r�@�Ռ��U�A�D8FX���0PluC����8��_�Lo�̀XI�Y�#k
���˵Wx=Z��ʊ�k���� &h���Ɍy%:w*�I%�s#|��=�e6`{���I+�P�ϩ�],H��7٩��t�T�z�7v��8���W�\80&��*���Ғ�G���G6���G: V#ù�Up�~Ȟ��A�/P���w/ By �	n�����C(�}7��3��)�?��d�������1�]7�M�0�nu���d���X��jlo�̏�O��료e#/C�(A���� �Z܇Ƌ/cS|3��=����zCSCM5�{��@m�zz8F�|�80C�O�!M�}�9��TοU�:	�jj$�s��~�S�y䇈H���W���ev &A�+j�@���{���xM�H+|Q'��|U��t��S�w�&�qo.��Q��=@��ɐ��z�(ӧ(�01��v��v��wmzv���h��,\�n���4���Q�H^�ϛ|��T8�Cy!� u�����}��� C�t���~&bv���5B�����>+���֪������~Q.��j�����O���7��a�~���*�u+|$H�V%ii�R��I��`��SO�O	������z���b��=`��z͡q���f>�~ڽq�-|w��?�	��$�b���]�t��m"5�����V�V���]5D�L����K7��ԙ�$�A0P۳?���p���{X�-L}W���˒�j��l@�K�64̒�^@�eKKTd�cz�dc��S��47f�f��M��K�xdS�X�_��c!C�*���g]X/p�2������Ft�����ޭO�Q��w�̰�g�8͵;���A�B�(;=Ubj�%zc*;b �����{su;TʋR���n�ƌu������^�~gGwQFz��$󽺨\aĎ]�9ߢ����Y�o����K'��=�AA-�@|��g~��|^э<�^�64���
�-⋵�H]YyK��t����Y����]ě���В>��X�Qle�:��E����Oq�Δ��J�����Y;Qr%�>�n��JV}�1|d�u�1HT�3�E����d1;�g�*�!�$���̶�vҍ*�s���U3�V��뫂U:#p�m�}�K�S=P�"9���{``�`с�}<��n�h��q�z�z�6e����U4U��߮r�<T�j*s1l�d�B}�(?;W� ��2��ak�{���7P ��n>�5{��z�X}��`��Mef	���^W�Wu���T�M��߉EY ���W� 2j�7|Dr���x�^�$��/�驰Wb�ur�ӖÃK�Fw�D�7���՟%;4�vd#���'��!?�Lc���&��\sݏۗh wׯ�φ�d#*������O����;���QЊ3��#�R*��K�@e�{�����(l�X�Ic �	���!����D�f~�|H�)�����h̡�C�i^D��?K��%���  оz��7@Mx��_u�ޙ�8���ج�����/�⭹87^���xˀ���'�R�������z�[��Q!ې#�:�+�D��#�|B�V�y�1��.�Ex����35�}G1�%� e���{�H���A�}�.��=��	�cĲ#X�A�C����nNẩ2B>�SJ�2O<8�=���U>v�
�!{��څ��C\i@� �/�Ĳe>.��˺c0��p��kT�H���X�����r�x���U�R�!����-9���=��M`C�e��I�+�u�.�<`E�>k�-/^�����;8�/�{E�y)$�Ei:�C�����rU�D���5`�?�g�aB���ZU'��;�	DN�)Fh�����4�6St>ԅ�b�Bk�M�k�A�ʭ���庸�M�O����A_ӄ�]�BȔU���¯,��FW?�LR�}tQU���!�ZF�%���BzG%&[�FXc�%��e�%�G����C�Y���L�Cc���b�M~_�M���~"�R�EI@���h�nyr���������B���D��]̸ɩd�1G~ ɳ���@&$a���M;
P�8�I��+Q%�)�a.o2���5V����
������+6$8mS{����;:�K�)q�t^qM��M���Wj��'*�A�o�0@���I[�Ҵ�l�x&������?�������a1�t`�����:�(���lCȬ�=8	j�Ol���:�k;�σ�2
����v.�F����\����1B�1wi�|4�6SR�X��N$�رsv5��P�޽y\�4z1R�L����X�k�kB�@������dFm��m.�b7=2��6U��;x������c�\ŚM��������9`�cl�*�tK�ǎ���l���`�<F[^:arJ�Ӎu���:S/ׅo�|L��Z��eg�R��ښ �T�
=8c~�R���U�M�ήtq���+}�(���ה�4D�O���2��3�����|]�O\L}24�����K�5��"�0�����'�x8����i��h��"��}k]�=[���ߚ����gSRI��!�ҥ�TC~���x���4�7����ɣL�X>c+��O_��i�_��4���I��Tiយ�I{��򛿖�4韤�F�౓҇t�H����Xf(���6��h[J����1�R�o�gw;�!&M:�����v@ן�I����]��{+��y��%�J`dI~����u�H'p)�������7����c
�J�x��	|SX�����ȯ�p��Ϭ䥄����4�>��P�{�akw|�K����߭];z�3���Rm�X>c##ճ�3B�L�YD��t+S:m?��e+`P�[�����|Q�$(��o�~F$�@�.�s[���]4O!�t�o���<e�//[�[��S_�֮l�^���� �a={�1׉�W���VV$��`��m�v�����Ņg@�T���?^�[o ��'*�Ҩ�*ɫ�UȚ}� PK   �X�X(rҪ15  ,5  /   images/48f3676a-8ce7-4f44-9cda-e384043a380e.png,5�ʉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  4�IDATx��]xTU�~��ɤ��BZ��CSA��RԵ��Vt������Z��6�HH�5Ԑ^HH�e&��ޓ���_Wq-�K��9�����9�;z�����lll.���rt����MMM������7��F9l-�7�a��F�)��t���Y--�g�O��)r����zݷ.VWW��v�����x�����&�9[^���/����{{{���\����`�?<��3�����555r�������}��#i�+���9	�G���ن��o������ a������k���;����[[�囚akk���u�3��q�{�OZF~�^�D����F#�|�^{m�낱�z`kcS���{��ƙ͍�J����d;;�u����c�ڽ����,�\��r�"�j6�cD��s��9r$�$mEFf�p�W��@��ƭG1{���?`�|Nb��ւ�%0����I���V�)S&���=��v)�vx�?~�"�!2����.����C0t������&%%����~�`0�c���r��&)�쟠�L��N��
�%��@9�-�^$����W_}5f̘�#F���)'v��g�DVv!n�e�j���7ET�	�-MB�VTVV@�[���燪�����􂳳��&�e�znO8��!�^�w�?ӹ�U]q�O�/ 
��:������Ouk֬���;H��Y����B92yӔ>2�喘��E�b�p�_EƑ����1q�DL�<]�v���7�$�<0�3���V��9e5�0���Ïנ����ҵ��Z�f%���_!�Q ��\��6cG�QTT6����A�A�Sgr��}3��$�mV��֭z����7n�ҥK�><O�?G��H��%����\���\��8!�ty8�A�a���=z4���A���N�(ޏp���5`��,����'�BPWkB�����S��:4�z���a���k��R�4�sr�J���v6�8
о4c��\̾�^��Z�<�C&����x�߿�|���͛�s0Kl�+r�/�Qc��?50?) �I77'��T
A����<d0��U8ѵO�>���A����*+))���hw�?_#݌�0��vv��9K��A��Ѹ�iصs#�}	4H��JMEҶmu�$T�Cy�z���H9_���p_l$��ԂkF�W��v��YUU��A��ENN�ܓ'���1l�0dff���v߽{���,3���y{�����WR�S���k[Q^^M0zEE/��)�oiY5Μ�Ŕ�Fb����P�������('�V89�1&�&L����?��Ct�-�B��y�񏩾��Oc}LA��,���	$�AIN�ɾ�������t���C����p��P����*�CYY�<K� d����0L�!�OC]CStLt𪌬�ōf��F�}	A�)A�р�WQbp����ǌ�C�]:�έ�3�j롩.N�J��
�����1��O=��[�w�V���㯿;����
���ZF��.�5ZoQ]E��p��(��b�Z`j6	�N�����ZJ:x�fQ-�E�UVT�@B�"#���
_�7O�[�bu��bתPSg]��ؙxrֺ͇���6�%��՚?��5BDwy�w��['�x�!,�wuyE������<�lܸ���?�#'��}||�͗������@����)m�m��B^�Q|�<��ux�i��%VqMM5���󲅋��-����O�]�`��n��'v"%���*�1{� 2IC�8{�6~�9FN��N~��J�Kl/�m^�(�
�e���5붋Ե�g\�KDG�e�Af6�:~�������ˏ�?�ѥ��&�w��t��HCz���q]�9WP: %5�fg�I�;�!�O��IT��7����q�)��MuV[q[��{�ꍗ^z���ö�����g���9TK&�	��
uo�<0(�^X�vzu�ǟ����B$�D����]�>
_?�	��D-R�Qe=r���$���р��6aܨ>8������r���6�� �M�������5�C��u���g��e�tw�у[���O<��Ț�����45��\�y�\�R���r�A��<j:��)jǈB��Е��No_e/|�;�w�h��s
F��t�GvR��^Պ�4ʆ��P��u��K�i��� �����Q|�H&��cL,���8�P� �`�
�$&��&�;u��^����ލ�_&�wv����0t�(������v�ԩPa�I����䆗	�yF�Lu:۶o����a��q�ꪫĵ͗��������;A���N�D���%�j��puk#4���R�/���l���vb���J:4��>��>' ��Ο/T���1x�1�C 	b�t:�Mհi�Dl����w�֭�������=0~t_�I�ǀ>0m����m��i��U����M�{�<[�
���Ftt�~ٲe���UDesv�P&�O6�С*$ ���O��v��oDii�" ���Hh//Į]��d�H �O9]X�22Μ9�*\�!��Ж�`\�h�-f~���!�v�Dj��	�/(r��s0+0J$��E�e�4#�>���(ooo,�t��L�b�n�P�~u fStF?�G��i��#�!o�����e�<o����b�A0$�E�����\�0�hH`Jƻ＃{�I�w��`�~�/�Ay[�T��l����ˇ;x�\���|�E�K~zJ�����6>c� �C��s�Αrt���nP^����gk������)��#i��@��ɛo-��t��і���>mڴ�W��J�F������ڃQZZ"��\�����J��K;v,.\(6�>�8�{�\t�0ss��̪_�����a֮]����#r��̾��TW�Y���.��� [��H�l!�j�N/D�-ߔ_|q��2t�P̜9���AuU�sQ,1���N�$�`|���&�o�ռ�<��Q;k�D	(k�Џ�k��&(i�G?v�5�7�B�p��#""���=��;ʹF�V��������8 ����>�����˕�m���9@p	���9��5��ۆ"��ϥTi�y�I�������D�'�^�z��z��:���GR�q��ho��ӯ�`�L��s:I,S v��b�m�K���8Q��%(�N�4� �7���UG��	�E�}>��c�x;�T�W7�#22T�E�;Q,* <B�Y-�d�>۩+*�Kq6�_X�n?V�?��L\�m�@ωI��.����}�\#�8 �r����˽L?y���y챎T�$�^������G��~$��v�h����},��$�S������BûH��kU%���pU�^xA�AcLB��Ers��/��{D4Ι[�s.����INBt�p�ꚼ�T
Ր#G$�/�Z�Z�%�˝���מO�J��#���̳FF��D��V�#ߓ�u�z�D3�;�����"��Ԩ&m(i�d�R:/w������Ԯ�]�wI@�Co/W�/,g��ɞ.F��U�JCF.��,++SI���G�Ѿ
�i0��K�HHH�����t;^.�g�[b��=:��ylOɱJ�����ڹ���?f��U�����f�Vi��e����PQW�z�TG���>^�����~9����B0��{w��{eU-*����f���K�\ ��w@���6�p�S�#Z�-ʖ�/�[n�Y+u�HǢ��լ����{� 2??��\�;���������̪,���6�����^�w7�.5ե8~x��^f����5|W��@���KJ.
��1�!,���Y7:�Ѳ�ע�8~�,��x�ͅj��V<�qS���P�ffd�K���H�M���)�A�:⾏��s5޿�����/�,���<��qQ��ݕ�-*,B�9ava
U=Kzi�$`߮/p���g!8�Eŕ��gЦ/����7��6��B������)5ŴUՑ����m�ݪ�@rS����i�q��1FAA�!�w���<��%��jL��}%���h�<�%���</�1���JuSr����U�E�Ɓ����P_����i���l��n�^��ߥ�:8:���p�b��<\pR���S�ѽ[>_�`a��[���Dx*���m&���ۧ��G �D��C�����(��1")k%^�d��?%��!���G͙s�rxt:��jjP]S/��y�N yQ�Z�0w�Ť��X� ��Y������c�3E5""���F���IE������O�������	�������kCk�@�-�LP6̘1Åꋆ�*��������I�7�`�k���K���Kg#�u
��S9�E�͖�>��i�.*!ƀ���C%2�<q�x�X��k:���?َ���͇��r�.*HCڙ}����͠������v�$
(3D}��g���bt_.�U^�!!����&��r�pø~�1c\\}���}x�)�\��i/% ������c�����Ϻ�r��D"^ǁCg���Vun�p�V�i���;*o���`3�Ok�Z�Ay���v;��^8�K��u��-U^�oJ�n�#FM����=��l�JNN��2�h������Ə�@qg��n���[��U��Se8&ޱC 
��DO��Ɋ]�K������7�kCk�@yM�N���f=��_���"v�(D��!q_�����2眹{x*;��J����4i��	z_����|��<aڴi���6��={�D�~�pN"ԍ_�GL�'�r���u�w(� �#�G����vn�\a��rD���a��^b��_`G��:wS�T������J6��oF
SO�}��
��tuu��!C���txee�� \]ݔG��b�q�����+ĝ+G���;N&�����Z��<e'*����9׫g��4l��qZ��T�����H�L��:&@!!!���kl�-���y+�eʥ��̔Á���M������d�"��h0��rV�U�[Ww_�;���@i�ɡ��7���k��[��@�����"���m��Όٹi��ac�9N�����J�?D�,A���*�n/ L�������U����#�`#n\u�n�9���# �F;��t
���"�X��\�M�X�u�K����Nu=c0&�]���T�=~Ϝ]fz:V.^�q��=D�;9:(骮�'�ꥼҙ�A��U�[��	 1Z�J���PR���&��+�"�PR׌T�,k���.�!ִ�4ڏ�o�w�r��_W��U�V�Ptc�+*&3��GDv�(���Z#23s�|�����X��C�r5���>�H�C��,�W�y3L�Y���n�^�.��-lՅ��o7H?	�w���I�[ʜ�˗��v�mjDѠ7@�CT�h:y �2[�7�&���v�ƍ��̀�����*b�$D{��	\�W�N��$Z��#G��z�uC���C;�;ث\�޽{9Aa�u����
�"��G�N�z��38'���Gj���`��k��F����@��؂���
��� ����8;��ж0����J͈�CTl,���PXT�������I����l3�O�.:�]�t��3Z��BPu�nx{+��r����UM��ֹs'2t�z9�^"�yO;��ƈa�%��Q�Z�	4��� �(9�^3��9������l�jVRrZ����F�={���jj��Ď@������@mu1�*
�i�
A�[�9�����ԗĤ�X�����c��<�w��7�f�Sv��8�$//�^<�5��T�/�b�
<���qi+�t�|}QiX�|vlߌ��18y:��e��4��Z	��lr��t��XAa^_�
�N(-���e���MS�L�M7�(:/X�MI���~��R����"m�HE�ʕ+]�m1�f�"q����j��	N�HM�T�t8Vb'a��S9����	]DP�g�I�� VYUmBډ'pD�zѹd<��pv�B®=ʠ�9[~O�ե����mr$++;�����	נ���>~_}�	A�>1��h�\���w´�#/�i]��+m�F�}���b���%���J:7�����z�A��ʵ;PVV�:�x�N�鵵�I��־%�����yس^2�9[ t�Cp�7n 8������;f˙vv�@��b?:744b����Q~���J5kB3H�̙ّp�&TT�Ү0Er�wpE]}��Ӵƚ��I��E���\Aj����|���/�ѫQWo�{��0�Rp��0��Q��N��W�(��NG�=|�Z���KEZ8�����S�{mVj����:���!0�C1uZ�y�����Pú�1��
/��g�'��Ћ���c����7�[��_=SM���YpU�����=c�y�X���+`\��Qȕ��Ǝ����⯾�2�$��BT���.��{�T��E�����?`�F��G�rYS�1[eԵ��
��g�Å�U��+�b�Vh����~����S��*��x�W+�qwNNo��썤})X�jUS'\�����+���h�l�9]5Nsa���T�9\imB�������TZ�
�*/��Fb��m7�����|(!J�QMrq��ey}}���f�T'R���l}QU�A�h+�^��df����ڌ�(-���=<<������1�lh�Cq�6��p�́��1Tu�t�t��R)΢�jp�]�Uk/Ȱdtgl\�)Ǐc���
���MoiD�
�tvvE\�A�l�	C��\��l��6X[4#�q�}��Ȥ�43��̀r�l�f�X��RM�nS,��^o���=�H��.Et׮5������&w]im����GQ����NM�2��0l�h1{��u>��X@T��4�����C����PKk�hi���ml~�b��z�bV{�=A)(,@�s������m��n�FQa!���ʆX$�L@8���3��";��'��<���YF���U: W�7�A���e0"�>:����l� �U��htQ�����-�ٹ����ƛ'�Jjf�BYIkr�_�.҄6>�k±%j �
��*drOOeе���	M�|�Lf�"۪�1P��څb8���Ղ���bS��H� �B-�U�L&oK��^���֖at��H//HLL����W������+�
T-���ޡ
Q����"�VT{h�T�J퀶�HujMb#���Csu�ʀ�Z�^�%� H˕������p�2؟���2<���/����)��H?���9��H����p����o,f���}��O�?LG��r���r�C15>��:����\��M����_Se�͍M)\�9���jB��w�/�s�̽��B��z�a����J�<Ԥa�0�p��ͦZ�9*v����@k�$jS+��?�����N-��ZQ�O>���'`�� �o4�N���C�n��+*k��3.⏧�潱#�b�;�Is��I�w��IW�g�8l�|��X�,�s%����^�6�M� �%?_�2u�h�b$$%��(Vޔj���>e�K��\��RS+�`��GLT`P^Ai*�f�p�ZMM-�����q�y��1�H>��z$#DTW_䂄脨�	΂�^���Aj5��˯/U�������jBZ��e$����w7��Ć�K�,�����ЦQ������`ΈwrrV#��ĦN�J@F��-7��jcgQ=�{����G(��;������O`7p6
�(P��=]Q^�f��m��z{{F�7l9�=�D���M��w݁��rt����1�;���lx��m�]����^rC�~�"ÿ�6NԸ��oV�]-Ţ�w�}7fϞ�Ĥ$�_��z!==�7�AVN1U�Z���k+-A���13o}^�a$�UUU*�Nb3R��URT�|j��b����{o� ����hޕ0��H�dN��3��:E��m5$��1|8Ǝ���5U�(���x_������[N6����"��uJ2�����V��R���+��	˖-�$�=+�+�Rb�3C��'��@^vv��2�'�AhD<�A��p�4���	Őa����'���UY)KggE�۴i�U��ֱcG%&G�(�ʀm�؜�X8x;���O�0.��ׯ_����'K����hY���ϡ��m%Sr0���dgὗ^�бc1H�ђ�wT�6l����^�@ ��֋�]Ś�O<�Z���_��"�yC�oA��H�1U�Uj�/S\�cǎ�D�>�NORb{Q'�P4��/D��kui���G����TkFZ-R�ߦ���v|����WbO}���9s�D���� iG7O�V�c����G�D����wg�GEť��N�>>�蘆+ ��v\
��TKs
�
�e�FGs ���E�0rYY��Y(��DN	@��zm>73��gϞ�m�6E�A�Bd���7����|m�Q��kΟ?�	�)��v�}�.#�Υ�\ȩ�	��	G��,qHL�pw	�qBh�Q�V�����/I���7B�br� �l�q�w�D���s{L��c�r�&�H.\�0J��#�S�&~ˠXI����f��)~���:8��������	���B�afBBBU	ڴ�4�0�2�ۯ��R��lRRR�ɓ'ѥK��ʘ*nQS;	XJ��L����D���UuN�Z%��o��SUs�9��E�E�ՠ%@m6 ���U�B��`���C����E3�Q%8���e�T�|�qMM�<�|�嗕G�J+�O/���/�A~:8m�i��D[[[�z�n�\p�p��&%tU����x�mv������%�g��0꺱��D�	������W�����R�7��o$�j6	:g�ڵj�����vS]]��?����T���ꤒfԉ�wBq�I�����|��~���(V`PL>�ꤓ����I��"��[�|�3�y���b���B����8&B����0}����}���XMΔ-��˛�:�ӧMFs�	�6-�c��WW�iG�jllU�X�&Ĝ{�B��~X��<���d�����.wk7�`��i�����Ǡ�4o�����U9Vj��x�b	�?�ߞ�#n��a����:�J��-..U��%An������������g���6hς\C������TUh�w�	�p|�~5}�駟~[��m���Ү��s�L��r@�?�d�5�_�Th�W�GKJJU`�u�va�:xz��U�PTT�Cl�Z�(�7�7 �wdI�����5�5��L:�U>���K��5"��{���i�RSϪ���MT���ЫI~�������\��qv�ZAig�0�$��E�͌��_\�b�QB��^շgY��pL�aP�Ѩ�޽�p��C)ܜ���i���wV��ᶺ�Wĥ�ѿOL̐�]�75-��!:���Q���m_�.�Q�Qrm;���������(�n�<��Z��%���E67#/�"g2%U���[�FV�yf�U�oz�3��i�ק�Į�B���9'&���QUmbE�]�J3}KeYْ���yb�VK�����`ɻ;���",�z;W�i1 j���U��*,/���AM�&(�<���f��(ڵ~����xN��)��!�fj��^%��I��+����Q	Zmml��#8ġ��ӗ�ͦ'X���{U%�n��Į9x4}q���C�x�֛�'�����܊�N�j�ڌIJJ�PZZ�<�<�r�s���ᡇ����Z%7��4��(-�$�Q��mc�&���D�:��ѧX��9=N�����SO=w�TW�����:'G��S)yU_'���)����ߨB��WK�( ��8����Ƈ�}�/z0���^zC��E�3YFѭ��BI�I�1((^�@�;wa��Ŧ�>��s���B[@U���P��"*��ћ�l�5W�:����"�'�Zx��-�@���yAaAV~����[u�ɭ��~����b���=�z�KJ��eߥ�V���Ά���
��oP�ZW���!(�Nppv���'�'�LT���#�h��;�6���V���x�Yr���O��ڵ�[�r ���0�3ΠkK5E����M�rИ߄�0D���<��J��5�������PS���:���ʫ�Q�wm��b|����x]}������jfM���6<�5U8��z��:��޽��Y�涭��F�;�ŅK皣��M��lڪ=�Z�� �&s����ֈ�:�:��jkc<|<]�:n���S���������Y:\D�	����oh4��[%^�^��ӆX� �����K�|2���	o���
�+@\\�*%+�5\}5��� 	��Qnn�(/+BF�~�L�-�˰1%�v9&
���n~[�P؞X?58� ��i&
��"1�*K�8#K\�Pń�!�!���2���	F�?�@�O�0_�:�ta���G�!��ov}�����@�l�r'�R�Ÿ��r�}����7�xc�e�����ؤ
e����	�1z�M�w�G.�ܵk��bk��5�e�"洖����hK(�j%�F�sؕ#}\���:�-�<e
L��*7�t#�QS�3f�kKo�i���p��)E׮��Neŗ/_�{ｗ���\�_?�t��L�=NP�-]��3?{U\<�7o���
�`U�[n����l��3���q�M7ހk�Ά�Qc�\��<�}W�^�HVV�����+���gD��%�[����y��0��}�����O��qp��L�3k�D!sSL�0���C��tm9i��p{?�.����fU9���[,������ �q��8y�E@���P�;�MP��رd̚5S�=_$�]mu���`��N$�R0���0⁩�e���F	6G:th�رj��#��4.��:���ľԋ���6�4����.��������Aۨ]�J���F����Er��jC�W^yEuL�V�Κ�TS�+0����*�����(ܧo���J@��@i��l���w_������O�(|�j7N��Qj�*��Z�����(��.�.�@̐2�,��lڴ)���<�2ˏhg
���3����l�+��,�3(.�k�V7��'ٿ6;��E�m�9{��4�)�ܞ)_}���ׯ��3���f�QPMi`���O0�:�Z����v�p������e˖ql@���ngN��U�� �C&'s�	G���-�F���m�Tk�*�bb�K1���T#���|�fΜ�v������.�~�[�rl����^[�����yStU]],����m�豘��+�4HOOG�Z�ߢ6()8���Y��R�i�i3��|}}o��/��C���g;P��aF
�|*2���}�Q^Z�Mێ*B|��v��_�۫�E6�{-�V+j�M�O7O�%
�.$u4u�A��a�UxgQ	F�~V�=�i+�����jſ�|k�o����n& T�g��s��1|��~�Fwq�Yg�*m��Q* <w.A����ѭ"���'��_�x��F^AX��6�@�],qxY i��D�1F�Ɩ-��l�6�r�mIWo8�W�^�^��	�riqil���si����E�>}��Q�.�3p�p��=w�>q=z�Z!Ty쇇Zz��|A��tm����Y8|䈚e~��5�e�wp���g��ܚ�E����Dx=�,�;vD��K�F�gS&6;٠��;�+|**I��dnl4������L~�͉ۃ"J~�ƣMM�/u���vDwѳ��g��0i� ̜u+��#�P�&$;�;.�ضf�6mRST#E�5�4q���yD��su6���G"4��A�F��6&c�t(�[�('WQ��pI g��s��j=>ϣޚUs�Q�
��0�0��Q�9���S�ƍ[@C�����~#�\��w��֙}�kM6�����������۩/���h
�*�MH:�=*2 ����������`��IдJq1�[���ٱ]DU�FF"<*J��6�D�����\Y��ŗ���^��DP�0��꜊ C��C��mND��@�~�����Q��Hr+	.	�,tN|���u�A�Z	������`�6����a�6o��!47�b��}ޞ.;^�n����c�+j���'�N�5=~l�Q�X߄����@����˾�����Ce�5:W#*���r�>(��������X%��N�f�� :���:y.9���衑��L�H���X�شq���u�����eX���A�E9�K!�N��Y��PJ��Q[g@i1��DO�^Bǂ����F��$gp��.�v�Y�ų�B|�+�~l�рhM�����y�E�_:8ؽ(Fu�϶ ��pp�UJۦ���Y�f�
)<�NgK�.S������r���p��[���Y	.�jFO��*�i������ ?w��܎�cHJ�-��p˪X�f�*ƈ�q�W�gf�R�����]YE��ƴ��n�i��jV���?U�� a�����zf6�2=!\>���C��;6�o߾**�R���PEm���[�J8v8QT��Z��o�]g�悇�ؠ�c������v�X�H���m[ML0��'�[�%Ǝ��՛��A]���f�H���PN�.,,��aW9i�8~N0.G�'DkֶE��^�8e��������v���ٜ�Gj����7�o$6l4��kX�uuqPHBk�%�k|�a�z����k�Z���l��/�Դ�\Q1>����;X�Ϡ��r]�>�(${��Ѧ����F�w�v9�o. l�m�pw�<�kB(�1%77���^z��{ｧ��q#1��3�O"q�QB��c�+/�͘��EDhmb�U9)���kX2�m��Ι*ns6N��AH�7�u��HM�B}m|���gΜQ�9ז�;9���ؤ�-�8����l�h�"5�����r��x53�x�ٸqc ����%��lGJj���ӆ�Av�ƭ�Q$�96]�1��T�*꨸B J�Re��B¢!c����㕝z��ϱv�n�	�0���v�l߾]�B��g�c���͓k���]v@�v`h���|�!��ĉ듓���,�Mn�(�ރg�I<��{]�*�Q�SZ��xhe	��`,"�*���K���z�nnN�c��Y���u��,�N��/�a��}�\�gDk�j�/���r!�j�����A^w�/�\I�w?��U����x}�
��Ӆ����5B�~��Zl�ڽ�h44�����ʪ��ʪڣv�9� ���4�X�O��=�7����h$��nf ��aU�^�{���`kgg�'��5���bt���@9X��e��k�Ag��{��p�HM���'Og涶&��x�j�0���_���Н4zl���    IEND�B`�PK   ���XdOv� +  �+  /   images/4b55d61a-3afb-42cc-8f41-c8483e8c29c3.pngE�TSM�)RC(���T�W�JT�4�*A@@��� "�M��t$�@�
�*��4#�zO>�o���bN�̜��������T���LEE64�u���
|�>��s����} �eʗ����&�T��-���ky������9u���n�pWs���`>����c^��~���N���4�7+z�+�}aO�����;�x���z�ˁِܕc˚w��w��-�`z�"�_[r\�����w_sɱ_����%�����I^���3|�����]/b�ݐ�		��t�!YO�~�1@��_Ǌ̢�_hDV���F"l��/�~,�kҙ&ڴ��݀�6Ғ?`�r+�.xc��=�3�Ma~#!����$��L;�AF.D���ڙo�j ��b�RN\lv��w�����Lq{7���P"w5�|~7\�VŇ�F H��d�T'�T�;����K��)��s��������
�H[�o��>���&��#�{���_6�oo�:$�N���ۜ������I�%{~�v�[�S����m\s0��V�̡~�N�S�tR�A��e��U��k�>�}��x���g�^m=͉����1�3V��k�iur���ޙ�T��b|u��ւ<Č��~]n��@KH�R"���a��.J�iy�-γ��i͢s���C��I9���l�	t�i�Wo~� �D�ڻ��ZI�����7���\{H�|�>2��k�s/�����긫�ݤu#ǧ�AV����2���%�)�.�������@�����k>5;�ׂ�����_�O�܉�*{�?!J��l���J�L0�I-ի���t�6wv=)/�w���p��':��p���?�7|Ω��}�m���ZT��\�΂߹�3���-��b�;�.7aғ��{9�V����+j��ř�ou��b࠮��O��{Y���õZL���ن���2�BJ�>�kλ�+7N�-}�z u'ǷnC��ʞ8���T�bFGv�� �8a��������u]���/���l�`2��'p��S�����n��:���=(�"����W�S���w8 +�o��Fn��� �u7/Y{�_7��+���c��⧟��T0��XyG��\����;�t����YZ���v���`kz��}o�s0H,�p��5G7T��Ͼ�H,5�����t����U����X���ʪ+:�M��]U�7��-�wP,[�F�빈�x�1�\��6Um�jy�""/�+��aI�^'���-k������0H�x�G�
]	L�%�1��	ܽ(��ʥ����w�#�����U�+�L�����$�X��6�_��>ޙ�%ְtS;崱R�_H���X2Y��8v��ڊ��'/7�er����f�S�<#N4�RV�h19CO��z��������"������l�.*�3��ޕC�K�;D�O�����/p%���U�ۡL<�23B��S<�SS�R����.�Rfw3G�F��@,hhѐ��m������O���U�3�CW�>a9����/�0��οW����I�����ͦ$��Z2B�UZ�;���7F&4���pz?�KbP�ʿ�K��F��،���1)5Lhp�Q�HRONW�{��o^<)���=_�l�#/z��%����$U���.��肿�Y)_����wz�+̂Waoc�C���a�
�IvEl�R?���:_���؟r���p�,�3���!V�:��1')�|�	E�Fu}�D�{�VC�6�z�Q�:c<�w;����۸S�q��,]�C�3��o����'��$UC�
X��E��G���:u�B�ҩ[�w�^��t嫬o�o�F
�01��lqwl ULCA��\F�m\��8?*�Ze�A�@^Ӷ�����aR&��NF�x���1EW�@��w��Z}��^�e����#(��%3CT�-Ń��}[l����%A0(���fY9���gIǃ��u�,�q�5�n&9���/I,���U�g�!�k��-C5H����Jm�/�ùHN%��p���*}[l��"+TBƟ��q��e�ƹJ~�g@-�5�G�9ꪳ�K�R�sl|�xD���~������@�ݯ�DL��"��oԳ�7m36�5V:��xǍ�Z�����Y��ӯ5��;r�:��퀃*�_�xx`Ϲ(� k��P��ڝ`��2��?�n~Ƒ,�!����0��/cFh���LȖ�o����e���t>� �~S�ɜ�����%q�XY�F%���OT��A����!����8���N�'�Lpvܜ���:K�Q���Sx�B��������FG���$���cRf���/��$�A����Vs/:�d�,_/�o{� S� �N��=ek�އ���DtĂK혃O%�ǬwƬ�f͗m���M?amO '�Ck�f>�d���Dú�&�iQ��qc�xg���ā��d���6Zl�v
	�	�+�m�l�3���-�v�v�^���ؾ	w2B��QB�2�qlK^n7%	��������D�l�䵫����X�~��S��S�Nw����r�8�"w��1��T�1��Zx�O�r�>�s��mA�B,kBX��4���:�WlW�f�o�^�X��@#$�p+�Kd�}�w;j��fS5��Rv��0K�Xo�fHУ�5�MQ�	���m�7�����2(x@�š�ǒ��RHC"m���d�'q�ʌarbp���5�T8=r\q��eEv�ݝ��'y�ۍoT
�:T� ��E�:�W	�����W�W��(�a!��K t�B�o�n�U�ĠˋO�.Ju:��$#vמu� ���t�>F``J����'�?��7Q\ՒNv.�:�|~��Z_�gyKd~���ow�,�ঔ�����^,�˅�6�&�x���1�˹j��6���ANjE�N#�%��[ƾ!s��B7>*鷖6h#���4z�k�h������16m}L#��;d�{��1U����ml\�/�i����@�8;�'��¾>��� �{^��@TZx�8q�slŻ��b�Aj�a���jdI���Ķ6��}��Nmu"�@/�#k2(!��"�	�
;�\�^<#��Eq���{Ģ=6�j)G�W?V�g<Lq[G2�X�9g�N̽x'�^:"׋�� d;z���HJ��Q�Ә������l�zPgF����[�b���T��׈�b��\+?s;(��W���7-���\����^�ğp�e��"=^�5um��q���ʠX烅�6=+=rf�li��G�oL�z:GF�#V5QH*�N�V��5��fR^��&��ٸ.YIa��kY�;56j��.^kr?��(�����u�ë���v}�0�M�j�:Ei��B�n6�~��� ��"+#e���8$п��j8����NFܞ菪^�O
(�����Ĝ��m%w	Ck�?N�gE���ڍ�W�$#�t뫖B�n,)2��H ��84�m�ݓ�>�g�p��\�A:Fʤ ́+��������6d�*��٥+�B�I�/�0��1�c����I��c�z��p�M&��
n[��?=��S�x�c��5Y��#�6�<������:�J<����g��
t�4?��
�ڭ�d����ћ6�˯;����~��
�26����2]z P���W�Z�N�z;�7�Ԕ6�]?�nW��������2����n-��m Ɯjk=P�k���?.���gf���<�KC�>C̏WA$��^"= ���X���r<�0�L�L�)>�x�)��ϔ�F�ˋ��=�W("�R���N�%wy�D�Qϓަ������1p�c�/�u*-�a�KK ���a��U��@t�.����D��Iw���E(e�1<SQ�q��|Q��{�b��S���z�� kV�>7M%L�Ypv�E�Kh��41�)�]���"�K�sاrQ��ܘ
}Y!���\Wq*�o"�u�t�d Y�{gE��Fz�F�������@�J.����mx@���J�h��X:-�4o�i&T�c��U���e�?�謫���� �n��E�*/���d#���X�uV���<��'#��H��ӛ��B$I5C�v��n��i`l����ҧK�-�Z��K�a�ts�K窋���4�
�C��p@�e��c����v��Ut��ge)Z�*�Yn~�OG��&�]�>6�d���v �m�"+h�R��>�1=�[�=ʾc>����?V��T�u��vp�qxoDl�Avr�5�hU�խK�5q�V\�M�-��9��tWu�@�=!D��\M���照��'l�J��J�;�d=X����5���+'Zy��XN+(>d	��}Ivѽ��]�ϟV˺�쿺n]��&���`A"UL g�>m	�?��O�?-�XU�/� ����!z�	=���ܫC��3�.��hׇ����{�rM�?�^J^��bb�a��H,"&�V:�,���,@�JVx�m:�H�59�6/�2N���W
?ʹ�]|��TISː�9�1^�w��ր�}=�{��e �~�����	!��n��)�V�����[�F�FϜ��K!��}�_:�5A+�>��As,¤���#Hc�f6y�����~�����l>��=�L
	_�*���_�3N��f����(� �ߢ���ń�ctY^)ôiI�H�L����s2j27s!�����f��!<�M�MkJt1<ū��4�l$�X�=����ۓk��Ͻ+�<��%���[+���e�T����k�&ȰG�g����^�̉�MC`��p'�g��n�M���N(e_WSГx���D��v{K�a1�F ����Z���[��%��^��?^
���Rj|?�|8�-8gC�������Ձ9� �0)nv���Q�� ��s������g(C�~�*�2ʽxq�n�֭Z@��(�W��U�Yx�2p��,hߧZ}B=D1.^\�w��]��mT���k6��qQ��X,�.��pYvF��,K�p�(�Q��ǠЬ�}S�����қt|���-�b�d���-�L��u���yB���ܨ�^ Z"W,��j{�3Ѥ�	�:�!��euk�^�VHnהB-2()󄸙��ڎ�f#�rW�"+2��G��4�K����$8)� ���K8z�k�J1U��>(/��5AOt��~���f��5s�o �\K�ʇ�ޫU,S�:I��v3|pjQR��m��ɔW9n��oK3��w�A��`I7b%H���"E��lwp�%�Yժ�Έ��_��B����Mu�E�5?����N�y�+^��"��P���*���]C �I��sw�N�S�M�Q�FPn���s�k	��j$��ٙa6T�r�G��/�emc����wO�h�5���oR�x��`���X�T5��D����qP��\��N��l@g��h��Zl[�y�+ r�`{��0�`��r��[�C�2E��<$vn	C���*���Q0uV���CF S���{��k{!V��l��5�=I����#����s:D6C�
b�s�߸�	So�%x==�����J�"�J1,��8�\T�g��i��V*�+ =���',y�Uat�e>�o�2���!�:\%m�݀D��k�EI��I�lSZjm�����O�~Z|dk\���J�	����|��� } }�.ӭ�}� ���@�`��	�F����$�W}�񞽕�(0����ai���޸S�{�i��82��{��}�����5�I�?������b��q��+�k�w���5r���eW�>tB��f�s�O�N���B!�I7 �L�D:4J7�x�oo�6l� ?�&�T�?�BЃU�N����tPK5w��Y7M�{%T�-G����� �7��N�T<�`H(ĮG��Hz�8z]$���K���pZ����w3W�c#���t(������П�-5���<������'����Św
���ְ���k��;�{8`�ЩIVn�6K���a��D������2j���.�4�'`. =2t��xK�D����J�^�>���/�E����~�9�W���@�5�FN��X�C�\&Z��{�cPb�P��������:���D,uQd����}���LT������qZ�m��K�O�L��\�7���h�N���%����J�!:�!���v{�h���$�(��hf�%}�,)2�����3�LКs>��s�a�e��+�)M���ҭh*zf[?��ؕ ���9�~�%�=k��%u�Y�r���Q�9�?���Ej$�i�a�+�Ȗ�����٣����qǍ�H��$+�q������Il����^���yVޟ�5*�X�DE�ֻ��3��M�.HV:v���Z.�� ���Lpc���A!藥W�C6�̟,i���te���p��a��`�Ö�њ�'���jW��#����oG�7��� \���Z&�63*�f������:XΔ���Ԩ#��i�md�Mo�O���	�U]\��$������� �ñ�S������ޑ1�F��C wS�&Vg�͘��m�z"zN,z�_"=���֯},��W�dK>M�le�S��8q�8������h�L��!���8C�vʽnJj7SM��4��;;��h��uP2V	ϊ�<��oq�c_>3Ur�}����� �&�=��O����z_�QJ��i�of�]���C�y�hicqf�-�5���</>�b*c��fߝ𩅛�hh��'Ȃ������j�}��!���Ea��\݄V����ɨ����ء�L[7D]������l�O���`AaR����=�{�wv~h��etٺ�;.Z���-�B�����X�O��9��$�9�����f���N5�*y����i-����Ԉ�VI��r�\����R��$��.�X���!W�K~�n�}L�Qo� ����7����Q�ORĹ���I'�=&�� q�L�����jA�����Y������5z#�fE3�g�2}��"tV�O�@�対�:��r��c�fT^{A�x��-CU=��� N_�{��e�p�����An�W�5�z:���x�����I@���U�E2,0(;m��呇�NL�x����A�&��eB#�PZ�\]���d�aPaI�m·�;(��ˎg[n.�9b	X@?㬰NMMU�S�&Ϸ~�Y� ��9k�7��{9��U�/>���/��5�//*}�-����������fIR���U��o)ٻ�KO�zy�N�"��SV3�B6�n5N�� �LFAJ"j{�_j�Ko��k6ϱE�k�U�x�Lm:<��r1R���[����,#^��z"
�OR}�]�x8c�� hI��'�S���$���#�(I�XXȗ]��\��*<@��o�����z�x�ތ�s,��gI$�6�id����x���OFh|�#�Pq:��N���☃a)�΅�[���{.q�y���1���^Gs��}(�J�-����a��Aq;Q��ȡm
:X�W$ ��V$����qQ�l��V��L�=zW��nSl����E�}�@��?c�ae=0|pV<°�ԫ��R5�\�k�ct�nO��-k~S��i�p�n��==,;�ҧw����
�w�mc��N��T/�tTj�������)ͿjIG�;�X:"�3�����r���� �4��r8���'��4����ue�i���<_��O��7W�����RX_�ȃ�v�X%O6F4��QƘ��lt��戹C)��0�G��ណ�j���P��m���!�u� �Ê�#[��L��t��X�ivY�B �6SÙ^��[l��D-����'���{�1EOK��,���Ԣ�s^���\�@�U�[r*lcF��/Oz�} �p�Ux�գԣ9��A�aA�4_��fQ�f!����������}ֿ��@Km�Z_��`3�����z�����^	�e��LG񾶽l������,P�̱�-��/�~bM	�̑���
���A	[z�9� )j�nW�aaڂh���)�9��]q�Dz`��:APwqB�R������bJ�����ƣG�F�Nk7}]e�#}[�_4����o cۿ��F����0��KA%�ZK~N�� @�Fw�Y�������'B�P,?�8�.�-B�\.Ր!#s
�t��I�r=�Ƞ����E])Y<� h#�=�h�-�_���I2�_��`�ɸ�aH(1"���2�� ������E�,�/��[��m��ֺ��zZB N�D��/�{[u��w�n���ii�2�M	wƇ�)U���`Ezq���������Q�,)�����J��ޚ|BHLX����`�c��m�˭u��f�lM|�RX�%�-��%�qW�cn�0�f�M�Y�X��r���>��~�+�`���۷n��#[��mf<�D����h�8�����b���X˫lS����ۛZ�R�{�����I����_J^�݂x���褔����'{�4��.	��κ=�*�輄����յ��LCE�JM��V��E�O����nޯ��۬���w��l��G/th
�C��Lx�Ȧ���B.���+f��o��:�f�(����P�>�1<�:5�`Sc��\Ot�ACR�%�O��CI�A���t��C���U�Y!T�<���(��:�Ǿ;���f0u��#��5���+��O�;k�g��@W��B��m��4�|�3B��y	�b�|��"JK4��:�R,�E��6��hD�8���1�(ג�v�C�ݹ�D��Up:����(VVW��gĴy3����п�y�U�����+������w��3���ZB���{b�kn݇�m-�;��2}#ܪ��r�-�R�/�(cH7e�Fw~XmD�=�ӷ��b�~��6��^g�o�c���LݣG�)h1�O�4�����p}���Z>5It���{U�(<�N�j㛩7x����_dia�쎯1�[�q�υ�յ�D�O���B�l݀)Z�*׆=��ӗo6��zyW�̓�nXX������4'o^?8�r�Nұ��'s�n����	�L�j#\�r��Z'Jӌi�"Ǘ�E��|�0�N�&Q�=k��[��;j���-�:¤@������Qǣ�͠a��H��l��%;/�-��T��wl|Y��������5b���=(��8A��"G���~	3�K����C��1��:���s_g�U�lj��0��5`�������V6��O_#)����A��`���밗c����W��i�H��$�s�!�W�qEגX�jt���)�/
5�<�T�w	��i���U*�0�CUu8v$2�a��M�Γ�<�@O�=�������s�����}�?wc%/��]q����ӻic��Y,�5;{K���b��?a������lN"ܧ���t�
��G��ңQ��S�V3I7ǈ� _�w
�thp<�H��}�vB3��<+�|7��2C�6V�b+��y��ڇvF4�����K`si'�V:g.NQ��~g�~"���]�p�)�$ٖ�u7��S�����u<��q'��z�k��T�ut����Z��?�jۚ���)$��{F >-\=̏R�8W���G���7y+9J4���� XX�m��;S��;��G"�TTbT�w�F���q�+3��7Xxv�+���`�i15>��YE��f/=��o�{��������ū�V�G1o$�I*=��MG���#�+� ۖV�1 ��@�2Q� j �������]W�CL�����B<�v��cd�Y��	����C�C�v������}Xn���o�������^<���z"� ����.�2��BGޖ�  ��nC/�h��Pd�ܕ����Sbe����(�_��R�M<�R����m�'ϋkY;�!���aLF��C�\W�]Ϧ����]�r*�D�X�R�?b��6Ë��w���D��rp�X��?|�қE0ll���;F��g�r��"XD?3�4�>b��f�.(]�3�|Ej��jj������X�i���S��)R�SFX\��'��k����9t�T�ב/����5��l����n*���E��a]y�u��na9Y�rs%vx^\�L�W�}�����_f(��3U[�.I�y����z��bԉ`����[8ʅǲ�'�2�n��2M�����]����T��������7����9�6r�ߕ"��.}���Cѩ��6ۘf������d���b���S$���]n�"�;ݶ�����}s���9��F����[��~K?�/9�O�MnX}.�PF���7��YH1 EP�%�D�V��eـ��~��sV�7�S]�'<��%��ڸ��Pv|�~y0�ʳ��<���'9b"����Q���������h�l�g���̤�K^\9��?�J���k�~W�G�T�!���A�$�
ˢ�T/��#w��J���.���c6��>��N�&��\�<n8kВ�D���|�ASR��Cw��6U>~76쾶�`oF�F��+3�in���7�n#
γ�2�����6<���7m5����5D������H����T���E�`�ࢳ}�秲"��3�U���EN��춃Kg�/�2"ѕ�78K ���m{�wc+���6�:]u�����2J>:]��Bj��֛7����+B+_�Di���<B�A��:���s�	��Ti���o-�1|dl���4�����s�j(Gջ���]L���Iv�]#���)ZS3�A���:).���
�F�h��̈�-�뉐��\�f�v�8T�Xc,�gp�IaU�]����=��v=�I�B��VaWTj}�����魚�O�PK   �X�Xh`Pҷ!  �!  /   images/4b60cb4e-ac73-4aba-afdc-1cf5937e57a1.png�!MމPNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  !?IDATx��}	��u�WK���hF�h4Z@�b��-˖B�b�����!���'�|b�CVs�3�q�#�lr�y/��`�1D�%����/�e$�F��=�VU�������Qk�A�{��U�]]]}����:.�<��c���7��;�a,�4�֭å��>M����O�Υ��KHQ�O���3)2�d��<���*g��{��y�>��2� 1-�C,χI�!z�����P	"�?RTbA��C��Œ��_�I��T�j<��0z�J�W72� ��O�Ua=QQ4?,����,�2>m!6��+����I�Z�U�����˲�	����?H��������'��@�jڿ9>�Ĵ��ʊQ*KFS��ea,�z������S<��2@!:�
j�Ytʍ�sc�O6wT�8҈�=�����{��8��w�}�V�2b�ب�L�"룐�,T�D0sb��zz�a(��.�sF���0�O(�	����a*k�p˵;K��_�#m�p����%�>Ҍ����6l؀]�v�RK.@�	���^ȅ�{�8_g֬Y�����&�Ju,�����'�Pۉp Ο�Ce^�Ч�9O�8?����ޡ�q��Ӓ�Qۅu��8':k��D=v7kN!P�J%C�6mb�e/HL*���7sRKe3��Y'��(�?�>�����T,���� �($S��,G���0�
Ź�|O�f d	'�?�"��_Ob�V*g0�&��Ϝ�_���p���~\<a��P��J���\��s���`�ԩ�6m��p���25�J������J�ta��J2��aZi�[� �<����{��r���`���l�[6`F��d_��-i
��G��3O�dP�rr�0u�g�����#�����CKKr�V������{0g��~��={6�� 
_��לƲ�0�B�Gɘ� +c#�nҫ)�Qt
�BTL�Bl��^�}w���ߢ�M
��(����AX����F��Ə���?�#Y�h���_<����
��u�~l!NuO��-r�*ʭepp[�n��/��H$�Wǎ�թ�\�w�u�~?���Ĩs;�r|E����� ���̙x�n������R�H��5�� z��T*����X���<��f����z��o�rV�L7ӛpk`�4f2��P+�4���F�{t��%е�[���R�r�-hjj�������9��c�p�B�}��B��d2�3UU��x
�3EX���gnGyh�H�@��l�@״��9L��_5|5���~J7��`
,�m*�<F��p R���6Q�lW���?��0�e����V� �\C�]�C����e��?0Ps����lm^�#�3�A�Ȍ��c}���=�Hs����җ��G}###�����g?�Ypu��X�-���"�=p� ��������9S���g�٧$P)�l��L`%h�P��f	��T� +.ML�moJ�+���
������
v��?1o
���*�����9���>2sC��� Fq(��"��`km���N|��8�<��OÄ́	¼744�֫7�,��������/�; s��E}}}�E�)�[o�%.굉�����+pݜb�b�޴�����B�@+[Fe1_�� H�l`V �L@<L��Ҧ*�Ӡc`J`$8��a�#̚9���yG�4b�e��B?kH������5}��ս8֚ru4�|�0Ϙ1#�����+��k�axx�� a����ǜ �������wމISf ��:�rS'����]aY�c�����V~��	f�6	�������	n��l�ထ�6n����[���SP�����ί�gYqGl��aa�Pp��Z���F���}������w�^9r_���l�2����"R=x��R^^�q��Lm޼Y����_��{()�ƒ�q��(���Ri��[�Į�EЫ>*�QP�M�'�$s bf1$�\yؑa�4 �!�4;0��B������S�V}3���`��F��(���n��=�u���������ß����o|����׾�5a���M?��$/ �E�>�o/����֮�]�E�<�:��ZrH�"����K(X�M�^�Zx��"&��4� �ad\�F�������L���$`�ۄ�?���V�y(%Ka���n�s��(ߒ�?�'�o6��܇��	qW�x��c�쫈$T޷��$P ^vp4�g����R��@	V\}�S�b�*�L  iE�G�j>N/)�����61�$lP���<�ʹ�N.S�M�O��bbQd���(A�p�!��撏�
�ޗ�;|-Ä�(�������W��+�濵�[innơC��`��Q��9�-M��ٳ�[c�e`�h�Y��#���]�l�"�$����$lF\�ZV��0�I�[�,v�6�
�P�;�c:b˄����F�X��Ӡ(�������Cs���>i�l�H!
�� 1===b��;j����H&R�1%6 �(���u��SE�D�C¦��5b���������c
�i�d���d�b�1%%�c>	$��F��$��$"1�|O.P�ML�H�Ϡ��M�)V�p$��][����,�%S�� B$x%t����M��`�hE�#��φs3�x��J� �k�!��}���|Zd�x@������yhi��h[4��%�1�����,A�����gP��Pb�x���iX�������b��lSŬP<@(�o��EJD�
�D���1%��S�����gkºoi�J���p�����?+�Ԫ��do�j`2�q39o�3�n��	0"H��'0�b��
��*%�!v��43k�d����
=��!|�/k���I���)g�km���S+ېH���H�+�uSX�x=���]��~�6+>LbH��a�l�v ղ�!@�����]"[[�O�X���nJvc�!n���n�h�9�����F$�D�3o�2���5Č�t�F�]	���e�Xb�1�aa�C���5�UQ�rE��e����>E�f�T,�~m�q�昿�?�+���3�7ǦK�`�[�������D��:�W�a�>�`xDT~r������}'+2��$�͗Б�8f�Xn?Yq�{xu�d��|�no^\���rP�(0�T�kn������}<�z1m�a�
Q�#�|��TBWC����K���KM��**K���q���'y�-k�܉�o���p��ĵ�Y��"3������v�n�d�`f�0CVj��+�u��N�VةϝvS�eN'����ἀ�^t��V:�s��8\/E�z�"�u��%o�ʦ^�������N�ZD`��NW/Y������k��`�	�����B�Ǎ��D�j	92r≎+ ��d3���긏���t}F�3�J�M6]
���	��:����͹. �����q��3�����
	3�`�A���zi��Ӷ���f��n��t��k��wh��U��~��e~�Su���/�>��z��,���F�N�5ı�wlv�0m�A�T͓ܠ\c�e��X�M�e��d��U�j�Xr3R�fȶ�e	W�/�[V�j^͉ɫ5��}{9��d�SU�,�(��`G�+���Xr�{9���-���v�_���ӧA-�V�<
��U�����z�M�q�&h��K@�@\�QU�����f�.�h�꒶���Z���ŗ	
}��fd�H�-EqYb�Ĥke�b�zI *�@t�M�% �t���3E쨧��O�߸��pDTLF= 8-����Ǔ]���?�2�%�m��R٩��Ldd�b	��T �!.�&�c��R���2�"�F>q*%=� b���b_-����.��Xܜ�:zز����5�-�"���z�\١.�z����4ؙ��a��M%&� 9[ٿL	L�2����Y<u�<Ҁ��m�t��<S��qkq�� 1�WZ��zYU�\D����.D �N�oM�܍����x�E�= �C�a�j��U��r}e�Z z0d�zE0r����L�^4	�5t��N��v�39�K�+Ki[/MT�ws��N[@��"�[P�r_��$��}���i��fk)���e�V�[_�1[z�NG���%f&+�N�1RĒy���]+�֨���J0 %�d�ntLUڡ�b܅.ƃ|Н>,����O�أp�{�;����֍��hZ%��&i��+S�+-��CG�ME%�Q���ȮG
��W+ǧ�f��IT�R'��$�O��?�&Z�_�宴/J������so�@=a�"���r�-�=k&��&��*'��}-BQ�Q���Ng����������&����M�윬����E��o�q�x^�	�v뙛&f�ˎ�҉����~����f���^aw��s=�WH�0 ����'�R5���8/�e� �C�����J)�)v:;�Ap=��:˭PLGY<|@!("r�"L~*{���sv��ny*~���:fHE��t��\�Q���S�4�>�BQCp+u3���H
M�!��" �.�3/��$d�D�{Ve-��!>'ʂ7�R�""�N3F��(9:�Hl|��e�����${԰�!��NH4ݮ'Q�]uR������[r��-�)��[i �¢�����d�i��+�t13�i�]��t�1�("r1īC�)s�In�2C��T8��a��LCދ"J�p	Q w��O��MgLKw�v ��&\թw)�y�[5bOn�U(Fy ��(�4��$]m"���b�Ʌ���cTF��V6YG�]~�͸f*#����""�.9Ə���Ԡ=(˔I9�N����{C^˰���WVS����;m��G(��*�<-�(��p#�]H��kY�#(6Q��(�TQb6���D<Rw�.��I�~v�9v����kKrx�����h=d�\A�423u�"\�۬G{���fQ�Q>���~$X��I���p&P��C�g�H�F<ڮJ����)�#J�o�$���L����R�(p��r��m���z���l=�v�El�ퟏ�.���p��;G�=������&�趙�F��mU��tB|��r�����Va‡�`��<f���Y2����&�ɹ����u[�ܜq]�#�${��\4[��|�L����X�yݖX'M���V¡��Z���~����>�v�J@�R�hȜ�QN#hDx�~���S.K~�$��OF��H�{/���ȏ�!h����S��@1u�3�i�L>E�#�H�ά��WH���9Ч��~"�����T>��<�D2���S(��T4[c�b�"wRM����vtH��~%�[�D��Uo����idɒh�I�Lj��Y�ODt��6L�o��N�9��?��^"�_P�MeQ��s�a��J��-�$��&J2��j́�b
s�MXv��ZQ��8fKSya<A��{fvu}?�~��z2��"KF�*A@��"�%s���f�)�5���<�� ]���/�IC~�	8r/?p�&T����0���:݌��K�,���ò(a���-bG?��(��RAgOr��gZ_�;3��n��^��Yb��H!�����3Y�I��Єi�O���+�`w@��y�x;�c�Xa�a��x��*�����cO�
��k�+�\�����8���������I[��f�Gd�S4]҉3j�`���y�������|*v��w�m2���Q��#q��C�x�~$��^�aH�c��0��M��j�H�o����R�x#*Q	����"5���YVh ��ޖ��I5�o`d;x��p[3���&]٦K)I��WÌ� [��O�	��J���h뙆�-ܦ~l,�'�$��d-n$F�ⲥ8��4}Z�9�~Y�%#*^9N��U��H �M�^������X�-�`�ѥt|4�U���R3p(�i,,ya4K�ܤ��T�[q��[R��
�V�$��EU}v��qŶT&�=�]C5bպ|2�Dʼj���M����$����+>؇���jε�rƓ�����`�$�I��X�:3#���dO=���GN}l�>& <~��SvG�A��P�r��>U�%�+Ἣ�t�M��
��>Y���~���T6�ALۮ�e5���Φkؚ�'�k�_�<���#?�t�`T4.��Ay1�c3R��3|r)#�/$;4ME4����CCMC��8�5���-W�+)<�J/ΐ/z��L%G�[��~Bt?�d���2s���3z�0W�nf�^�gxVe~�B4���i��_���2�{
\�ȂO7��π�)��!s�l��|��\9{���\Bb��Ǔ^��$�1rL0#͊���|㇧�u`�lnb*�b�_Xi/��W? �ɟ��դ��Q0(��.��ߌ�Y��+����"�T� �G$�_�����(��?���;�8"�^YY!th@�� ���o�.���;@���w>��ddX�RN�|xb���Ce�����)}"�Z��[���&�wx8���t᾿8�^�u7�Ry^�����Ւ%K�q�F�`b���IL󋵫(ʊ�&$��S?��-z��7,�M�f�K�}�����ja�L]������y}�,��d���_��=�"�����;g�]�`^z��&M��իW�W^�q������}��u�ҋθb���81ԃ�is��.;��[3f�&ḫ��t ٿ��a�_��0T���|����GĢ`���Xw�5q�Z ,/ ���%�(⭷ފ'N��^Y�?h�����3R9�,�٤b����iW#PYw�q!�$�y^D�F<�����N^�������* ��9��}�D�y1I֙wAIg��|��Çg,L̨�z�>� �}�Ylݺ����� �������r��%A�}H-J&�B��6" ���+�2Qpɡ]0�����������$�������ʸ�������^��1W���O��{7y�Ռ�=*V�v��M|��p�u�aӦMhiiAdd/�
莖��?Q1���^w�(v�o����]�U�k@�j�����'pD�y�~.�Tt�����<Y�%��)Y  m�|>�����/�CQ�����X�{�ʕ�o�C���F��;Ώ!L��_��W3Pv|�ҥK�x�bqq^�o2*Ƕ����4DWռky:�p]-@�r"�Փ)T���[�d���ȳ��e�Ć�#�G>"*�Γ��c:����/$���6a۱e���V���P>/�̫l3�׽e0����j�cɘa/3䩧��}��'~��qH������`O!��{ёX����Q�wg�O�0f".�_"�'�B�W�fb_I%��W�z/���Y!�=��L%a�/c�`$"��\����(5}����#����q��A,�U]�s����\/+��'0:::��}c���y�Ν;��ى;�MMM�B-?�c-�;���|3�o��!���9⌋���c=g�m��<��C���'��|A
�|�39�����Sܒ���c%MzxLڗ�!X�Ӯ�L���y�'	+������m��^�X2�P�����Rb�Z�[�l)��}6)(1lmm����E�6}�t��B���3-�j=n����(1*�/Dέ+u8A!�@�<V�0/jƹp&���y.�������=���b���DL����_W�� 4u�Ykl�'08R娴 ��ɁJΡ�l�����K���~�m��~1,	���V��LG����(�9�`��1�uK���aC'��v�?��%�F��܀�X�{��W�O��8|�E�r�N�X���r��*V5�����(����2��xy�D>��+<H�?HS6@�b������F0o)��Zk��7��zWW�w���W��e�������U�V����?Et}(�3^���{�?�)�f4��Ť�h��
��O?�@� �����&F[�Dno�ɞ��QZ�`�J��)J���Əo�����RJ����.��vG�|��$�!Z��CK�)�{�^�Ϗ�	�%�?BZhT���|¡��vv h�"F�<3cjK�T_[�%+c�&tM΄�\r�!z��֭[�K)��B���5E���Du$�
<���ϕ��<)���2R�5���m��Z*���s1ip�0m�項�>zwG(�����F�wM���_�� ( ^QCyz�_�:܏�s�GI���˿s�E!/O�9�J}VGʭ�RAʦ$E�c ��2B���P�$ :)�kD8L�%��;фCgk��hau�@Xt5�H�~�}oL��5R��Q�N9D�����O�	$Y�t��	E�`��E�o��R�]�<���p�]� ^�Z�V�yoϓsb���gw��=vƫ�[@
���6�y��C��&E@ƙ�0Ǽ���b�    IEND�B`�PK   �X�Xd���Z �d /   images/57fbf569-4147-4eab-87dd-5f8b4e7be3fc.pngL{x�[�v��mۍm6��ƶm۶�Ickb5fc��s�9��3�<��o����]3{"�$�������|��U� ���eCC%*�N,�?�N�R*��oh�p�k{IM'�������*�@!������������)�����������)���y�%/�����{�������:��v��9K�d�,l1(�=B �:(n��-4�NGC�󊮋�J��0�����=�I7��L]��t��#⊮��1 �+�w{fT ���?)���#�1/"XD�e�$�#�0;�#8E���8I<x�h�$��d>d�6q0�0��'-g�>vE�kv�n�<��x*��_����_�6���� ��¾�A�S�Y��:"��_^��}���ĸ�#�4�(�}��P�U��%4�<*6�oz7��V& ��������Z���;
_�/a�x��+��WC�#0A�A�����?�
-xDG�@Q��OO�D���^�v�2#����riADG���[ �M�����G'���G �k�O%��Q�BN�`wr�v�Ir̎�?���z�����$��m`}�qp��v��_�����VL���Ȩ����	|x���������9t4;*������ýE�13����>��D�Q�Ҟ�f�{�����M�	���C�����T2!V�}�\* e���d J?�<��c8��A<��fǫy�F�J�<�o ��ޱ�g��|(����>���Q��n�4��9�z2�.��'�Y��' ��b�� Ўa"�9����l��q��)��l2���Jdju�9�Q����ic�6�l� @���T��SH܇���3����L�@d�7o����͵F���-�\*���2�}������uHa�a��xuF��?ⷺ��ާ�hz�LR��V#*��sfo~d�����ۤ�{F:�zӡ���C��n�w�� �ɺ^B����R �j~��l�78���z����L�e6#�C�DO��\�u?��s�����.r�_?	���G�F�7t��I�Q���-;ӂy����x��HJa���W��K}#�]
?G#mT�����t���y�X0�;xC���e_X�-AXuk���ֹ�D�G�/�cC�,�<��_���\R~�����'F�t7�.�&��h��V#9^�{v�*#"��~%LW|�R�j�8��,$X��uá`�b�H\f�kJ@�(����6�S�@��'��a��I��q&1���c$�_�k�@0�'��YSblU5��)#��ԉM$����$�6\t�����M�T��Cd�KJ��r��;1>f���k��e<���F4c���>���ť��ϗ�kE��E�ޓq�C��>q�=ٯ����݅1��6�'9�>]�`0��l��DRvv?��*���i����gC9�^r���=��u��`�4U�:J _�ܢ\&	�U���cѹQ��,�����K#@��N��M&/��_���?Os*nҹq�W˖k��k�Δ��
j�l"�y�c�<������<ޝ��ld�U�4�ʜJ�h8���V��?J���7a��ē���N�P쀁���X��a���OF�ُ�jY܂#Ç�� ���a$�X�/'�8%�M�S���Ҕ/���Z������߈vfP}��K_*h`ٯ=9�}�zß�w?��q�wSfS�8�7CQVf:t��B�f�|�"�H�X���	?�Hx�«�H�b~'��T��.)z�Ml��v����b/yP�kZ>[����b�h�~�̈́8&
�d�����ƣ�+��b�Y��?������؃���9i���i)6#{W^���`P��4��RO��r�7���m=�fqQ����f��������o���
�L�t��p=���M6�^PN�{}�L�f,���բٳ�\~Б��Ν�+#p�e#_M��v�~6 ��r��$�l���zv�(3�\+[�"F+���J� !H>~��i�}����p��]�����a��U�&��G�Z��B���G��⛜�h�r��-[(���ՙ4�c�;Uݣ4�-��_����^�06I�W�r@�
#��kzg�w�$��>x�������}?Ż����KQ�_�?�_8yj�0��3��>-o���ޟ��(�{�0GA�~��/<(�䫆�c�>�|��q�auw�A[�,��f�%|�@�p685�:d�r��L���{�k���j.���:ITm�����zvg����E%rz8x��:��J"�J&�����N�a�a �F��H������޷�5��%c(z1.�yc��Xrh����r����sh�5��C���g��B$WX�`�"�#����ѾO� �����<�N��c�Jd�m��2����e�vM�~ϧ���ꐲe����$r��R� �����\85H�o�w
�塴���F�P�
H]�T�N'rkv^H���kÞ��~܆�*��v�h\��=;�����7�RA1�l�����BѺ�p�D8I�W1\@�o���D���V�xs"�� �"\
�WT�\HUR ��d_�'meVsx�9�E��Am��}�$����W��jL�?M�*�t�$����M��􀌨�#��o�*	3�s�b,����61��[U)�,�x��5TV����*J���c��}�ΤK��n�Q4��蹜h<(��[��u��ȏ�� �˞���D|�1hI�캯<�`��������xvѣ�$r�B2��Λ Lb��`���o����a�bK��Ͼh�Q�H�䆦�1�:)d�T��l�]�m`c��ľa0I�c�I0��3��>d�G(W<f+1̘�V2Ǔ�1[t ğ�~��E��8=�O�$j��n8�w�V�PZZ	[lFI�d�Ó�څɢ���������ʏjɢ!I�ƽ,&��/"���&�? �u^V��E10�1�d�����"�+T����9vu	�!p�X�1�\'Ӳܔ�!�6�^²����@���*�a¹�w�Z��b)��x+�;7��#2Z�j(�@�̙(bCqiJ��Vn�4�5�Y���Rfы��oP�2��Uڵi��!�&��|U;-X!��X�K�6�?-m�/P:C5��z͕=2���{_HF�쥼���9<��n;�D������Pu�`�5&�暛Y��Cݢ�$�߉�A�KOU�>�p8�B�L��R��"N?%��y9|��S⫭V�ʆ.rb�g�#Lt���E	+"��b7�'��PO��u�� vFIz�b(k��q�֍�w�	b͞�1I(��Τ^	U��L��]e�Ȳ4O�.������RI�'��x����jf�X}/�v��@�(M�dExD����vb̼,VK�$z���%E
�uP�h�t��-�Κ����ӫ��ȢU��I�,�a���w��щ5=��d��l ��n��j���U T{r�{;d]|^��?r�5;��QC������L�M�L֎�h�DՀp�B���o�Pǀ�e�T�IѾ�Q�#7���0z�#S6��q03�U��ß*I�y0P���e\�9_O�6%^ͷ��bF�ud=���{I��lz�A99)��&DEC?5��'7J�p�����C�.rn�vw�H�U�ι�ExwG�Y�q�(�˕��ix�p���b^��߷���~�90h�)�	�<������&)l�)DF߭���`;�P�*mQ/1�u �%A�´�|m�@�̃ 캧�~���I	�0۠��ڬ�}�Qw�;��
U܏�U8���5`��Y�r53�nF:Z�#�b~���_A;��uE��e�ʓ�j �v:�����;��Ո�.�,Hx��"���Q�W���V��,֩r��l|���Q�Q5�����ܾ�Y>���܆�<��b|\Y0��F��o[�
��?D<������z-���Yy���&Ų�9�R�d�L�A�p�E��V�W��V鬌�tX0'͇=4��F��6��*?��3��X~T~�%�{n�$���2쩗���\
��<�.sFf�ґ �D��(�U7iP���<.ٌH#���ș���	�^�5_PY~%��[W�=ݯ�D=�Ư�Z�`:n�Ow�$�r�Ѧ�^��iu�����&4�*+�8J�(3O+h�Ms�_�W� [C≺z
�'���0v$Ef�nl��� ��W~L�bS#<	r)��͆�w�JJO���3ϜC��uq�!��	<��g�6}KP�JzA��1]>� �|�#^��a��bX)Z�nTe�/�O���*����iQ�q$B�LdNC�Ø����=�W�.`b6�\]~���y֢+k���l���4? 3oeR�::��#G���C�ʛB*��FOf$��:���])�b툭2@4�F�+X��~���}cf�:��I_^����N>���1�
I�,�b��pP�7a̵�ݿ4�U!��}���A׮|L]ko�5KA��+��R�ao���[u��;ۗ^o���*� ���A�Eg��*���O
�z���f���VԉN��f���4e�z������ .������r��{e
O2������e?�Y��	�1�pr�q�*���Wɉ��?sɌ��n��f:�/���V��D�n��ǰ!rPk��D׮�hS77�����F/����H�`���}�T&�\�r��Y��_�>z�e�_��m�Ō�����>�F�yk,2.������xV�K���E�J���n��l��mE���~��!�',s'$'���N}@��ȃ����`Xz�zt2+H�ra��%:V�R��d���  �����*��(_�'���ڤ���8��U��eM#�����7�Y, �G��0E} ��t98r�Z8���5�,R+�V��W���Ӡ	ȋ�,e��J�����N��:����iiV��nX�L��G�y)�D;��~�YZ�g�EH��y$4U�u!:���L��Q�A�/�p�����>��hṄr�٘�0��C�>�6�B�M��5-)8�W��%�z�d�b[��k����*�G�U�G���œX�F��ev'�ȉ�t:V�lASoJ�32/��4�D���+�{=}v��DoUl��n�~� >7��]�����\:+	�>/3��~D�M<&o��M���u#*�8��Q��ƛ�ފx�o��@�n��u�"��hs���O�+o�Ђv��b�^%RuK���C����$Z�_]�D�/����B1��]U͙�WW����e����" s+#j�S�P߆Eg�^'�OT�gQOC��'KB�RU�5��,꣔Y���)m�cX��+�WT�.�����6��:�6��^�j&���殙�1�l��9�G
+:���H#5"{ѓ�.��A+M-B�{��R�iHZ^�.�x��X�h��!��N[^�-�p8�~��Ȑ�q�dڡ�o����-���G�d�}^�鏑k
�4Y�4�$1X|�*"F�Q��A��^�"�ݴ�e�8����
^�ij7��~ыz5�D�4\���Y�H!�䧭�r/X	6��F�&+)aY��GS���$���[`14tnT�Y���6}әh��s4C�I��1[�*�+��,���a�D9R��1�\�	�e��b�c���xK ?���F.UG��(.��#�a�3��0Y�dWU��W}jM5odӹyP��*���l@������.X+���\�O3T�hX=]8O��x��"`��4^���&{	�t���rr��Z�ăk(��w�Zr��9pӽ��7��-�L�W#^�SA�[��sm��zV)貈�,>��#ͧHe���a`��q�m�f�G�-4஭S0���齟�f�C�d����D[C�K#����Ꚏ�9A�̾��7���U� ���7djI��^5�������aɆ�X�&ɻ/���пjJ6�# _6�V�,%�q�*��Nt�cج��Z�F7��
��t
]����J���0d�`��y>�T�&9��r2\�/�5�$���f�f����V���&׀Ff�@ �l�Qo����M&h'd͒�Q�`�����.�eP�����^�e<�?�3ѭ�
<�Sc�S�H�?&ݜ�J��j�|�yl��3ثv3�
3'VF^&��wŨH.D��~����l��ʧ�@Ά�S�5x�O�d�dS��� �ԣ�ո3!�3�1ƈ6�P���=k��WL{?��2Hd/UOl���3&)K��9s��J�a����;4���o�[;�b՟/��{֪�>`�$Yۻ�2ApԞE�?��~P.
��T|~��
{��.�����)nq�Ky@Mς��i~�~���Ma�<�ٺ0Oc�G�F����`7�+̊t���
��[r���sHW��\.>��(�b:� <���Ij��	I�:�I�/�&�"���wm�q���9�d��bPt��aƊ�*W�3[^��rt��&N4������CO�Ȱ�o��R*Ů��e����;��<��=�����fE_���zv���aVoȭ�cőXY$�H�M�6�5����������8i�'�A��k(b�����7vj�f��?Z<���i9�L���C�d�M[�8���7�?��At�>��]���Fү�	I�g�������k�k�Q? L�'�۞��N��պ�AE0uf�õC��A�W�J�:�����I7���Ӡr9أ0��a�K���$��������i�=؆8蒹$�Kc(v����ԋ&6���T��M�m0zB��\������%�'(�H��8u��O!��Av��i�oy����[ʨ���!�0�u��)b?��]߬���\�Zt�W�����wwl=a]��p�cN�N�����N���ӓt)<��H@!�N��$�LY��s��_޾L���߬m��z���^���,�:���L$,ԯ����u��І .����9X�fޕ���^O#3�"��~Us�76��4��Z����q��r߾
C'`���@ь,ځ09ơ8���vK���G'���hݏpC(h~�GHy�r��d��<:�(�-��0�X�S)F3u���p-gv�ߡ��d�64�1*�B��{��7�i;Zn�hu,��wKI�WM�G�wX�w����,��Z�Y-�%tw�F�y@y��<�V��~lG�`ZVpV�z40���+*���ך)\��b�,��K��n7Uȫb����S����N�$�#܏8s�4���R
f���@z����Z�˝�#�A�8?[�������&�~������/5?ʥ��� 7� ���T�F��#�e��RFJ��M�V��9�.�C���M�o8�k�P묭tm��y�����J%K����Z�f�K�EE�H�cW5`N*�9ìL�$�y
��}��i�b�
�{J���Uy%�ҟ]�(���j1�tɵ�j9��ȿC�nMKբX+'�&v���+����9�k�DK̀a�m�Ken+�̌��`;OmA�f���ʏ��fHQ�jd�?�.I����L��Ö���{�gjH�Ŏ���<o�b���i����zj��Ϊ�[4�'�u�;0�!>�1U@�&m"w{ ],���	sL��g��
MG��FH��|q������R�z���z�p�-���7��x�n��*{|��_�n6����ŽXh����ӈIf���,�.����MV���1Y�x��!Z��%P,�1����p	S���CDÔCd}䯫n`*h\,¥pqp���4e|�����v�
{�^D]�;���*�� �
�?i+�~� ��K\�t�-N4�%��KptTc���j� &�������̜[�7K�6�9Z!�a�&�? �Єu�̧ǖ�'�gv����5N1f�Yo�P��:��o
0�L�=2�t�n�~�cab�d�_䘋�Ӓ���%���A�Z��OO�("��d�ȵj�w2�K�xy��ޛ���]����}�.<�X*��x�m�$�I��[��E�`���P�|�H��?�ÿg�/�X��BT{q�n�z$�V���d�!KR�G�Z��ZKx�;��M���� x �k3�Wp'jI��tN�)�<.֌"�Vz���?���N�s��H�1H2� im���d5{���X__ól���&�
�T��q"����.ђL�N�w���9L�Di�.��=��uZ��X�l����Ϻ� �6h��"���s�Ti��mM��wKJ��	�ةW�j���T��䉺���~ծ��o�k��8�>��$d�)���Ђ�	I��+�i��[~�jM	���� ^��[���b���m��R�f��r�~Xk*�|z\Rl=u�ӷ[ن��X�W���Z���j09�/l�3]��,J�!p��#�:�{K�v�D�֜"�i@�����H��`��?��% \��tP�U��e*����a+��s�yyv� F�4�u�~/����
�p���~����c�g�i�+������d ͵����7rDO8{�"�e5�ѱ���c�!�[���/7>�G1b�V���$r6^��/*��`'�=0��&�j2����,}͝�f�0Џ�.q~^)�l^��>h>a�r�48×lW���7M��]���{��p�f��fr�EG�^�qyC.�~x�cn~M�&��DDf���ʳ��h,���p4�u�j_31���$���T鲯�9��?b���}��6�]"��t�b7;]�Y�z�9�i=)�Lk�ҏ/	���fZ�ֱ�x*���j��.�5��Yg$�Th��!`�g�r��2-���J���Y���N�� !�/��Y��C��'I��8�c�N�����> ��s����[ $��2��bό�tפ�n���?�i�o�Wʄ��<��=\d%���+��XQI�^To�i{-H+d�us�Zd�߃Q�P����|�vra�Rw�T%��J������k��/O�MB�(�f�����EjH�s;�'�0�{��o�~�B�F��v�AqKQH[�7���A�C��"�ȏ]F����N>���Ix�����s��v���ry0�_�j�U`�[	m~.�T]�\nD�j����:�����
=�6���_�V����BY�÷�Q0i.�:�7�*X�H1>�� ��^,�ћ�`0���v�W�{����z�X�����qs�O��鈊S�C'�@�WK�F��� 5	�Q�����k~`θ�J����{�u3�z5���"m�C�*�Ķ�?��U��
 /�8���.��!�b��1=�ňf�>ȳ��r6�'��TC}�f*����Z�SƷ�Q�!��������5�Y���Q�f&�B����qlw��m����L�_C��Xg�� C��f~�B,�~@κ�9��X10|�@ܙ`o&U&P<p��ͭb�ms�8Կ��6����ǟ ��%&��i�q��P-����@�M[�Ӣ�O0��[>ӻ��|��ٕ�
��Sy�T@�E6�l�����=&^>Y�x�g�o�8?`�&9��� �·ri~�����х�������T�&n_�W�2�0��d�6��m������ ��--ob@��Id��x�w�í�V���qg��ݭ<������[s�\
OVٱ؃>
�Ee�wkyU@��S\
�=$%$�c%7K����j�4�(��d��^�s�a����w6:����$;��qt�&}�~'���u�g�5ȥ|OT
ʓ!�C�B������_�=t�.������"��r�)�v1]5�P+����0�h&����������T4���$�z�D!?�)ڐ\uL^׏�y�V�����E��u�V������_�=���ůӦ?���>~u��7U�������ٝ�7-�5���m�
�W�~���\����c�t��1�>�"z�_����_,���ҨV�Ϟt��K<�v9���n�$�F�܉�%�h)r���^����~��x�_)K�!�T)���[.;w�E],�o�ȟ�h1�2�\}�y�Ђ���RP��3`�xsrk9KV!r��r�@*��?v-b�W���C�ն��d��Iࣇ�K�b�ne�<�>>Q}��<qq#��V�����e�z�VӔorK1�Q6�f����pI�����*Oy���%mc���|�ܵ��������t;͔�$�`T0s<f�b���"�BU�́Q8X/����^�[�(�K��f�-˨j{L�+�9�N������d1�N�w����2
��~��<�Jvu���i�����A�h7��	y��@K��_�f+��;q������5�Xއk�3���7�h|�/Z��+��D,������f��PB���������^̂�J,�	�n
!���>�9���E4�y���	^N�v��N��a��a��j]+���Xl}��2��F����t�����, 3ʬNa�����[B�0��t�"(m"ŻF.��S��{������h��%�gM�R@i�p�-Wk�m��ם`�~9x(�y����ƔZg����0aw�1��O���F�4����nn�48P:.�Sw9��$��4c��/��[ʬ�r����C�G'�{n�CtZF�����q���
aΪ�F
���щ^��M��	�����v	D�^7E��t6=h�pdm��6���G}��N=&��8�uz��g�8�c܌��9���'��OˑN�y��o��S���Cc)�u�Ra/��m�樳���1^��zg�O��/Rd�[��bo�I�n������*dB���{W[
�7]hU�ɜRb�ě�`�_���Á%%����M��M�m?h���=G��
>��� ꓂	�a-�Vf�b�����3�SP���nf�3�����d��p
������c�の|u	f���k��i�tMu:�m����z v:T>GA�~�`5�m?�}T����Ϡ�ɷ�"�
r��9��\�l�CK���"�<�W�9Ғ~(�8R����;����C���mO���M2!�kݢb̓��w�m��Кo3���z�3s��h'-O��Ԛt��ڶ,��/�ױV�k�^��.�<2�>jwׁ�0ئ�w�I���)K�+�#;GAx�.킾��M�t�2��u�Ӛ*�\-�U r�*����ߐ��#�i���߸W���NSk]��۾^цz<���Ԍ��o;�Q��E��Ӥt�
!��d%x�ڎ��^h
`�8�N[z�����΄�	�8�'-��Jvۓ�?�5��u��y�(ѩv���s�3�>���{9X���^�����&��o>!�'Aݽ�t���̒�����)?}�O������c�Ǘ�v7:��q�o�Z�k������n��I�f'vU�SA-Z�OW�/`�)��6I��_�vGJT�W���S�z,�ॾD���o��r\Un2?H����h�
wr�D��Y�-��8�+��B>����a]t�֙�ׁfq�d3���ǲb�X}7��8b�}0t�YQG[��k�rX��ӑ�'o�=�l�^[��s����)�>��,R[�%���d!������fA���N:��t<��]J��6���gԭxz����Y�l��(������U��}�P=�z`brU�`�D`Mx�R#�s}�9�@N�T�q���}ά������W��G�Z�z��G%��cZ�F ���g��V��*��^�����
ƴ�2G~���ͮ1!ߧ�n�x�Xo�<Y[�gq��a+K3l/��t(�q?F�J��B���ИT�)i(���s�
C/�w�{��������Z�]�y��f"�D@�$�m�4����y�S�A��ʹC1o_���4�̼�	�~�u�K��G��%*JZ���6B]n����O�˥%��pfמ�nyBN�4�TQb���8�˪V�n;�h�Q�"Q�+/u��*��X��^�J���&���w�Je���o��Gp�ڬT��#��Wۺ/�*8+�x��S�|�l+!��3p���h$�̥5�)�'(ƚ����  ��2��մ� %�۬b��n(���VEd��g��׬�) 6���= ��y㾦�W���0Xk����׫�Ǿ�*�W���J˞A�|�f�;��T�5n�6����0���끜�"�ܽb,>�WH�e������ђ�pyS��{��Xk���b����\	Š���8~zEN�-m��C�?j�f5"h�A�~a��0i�ΘRhil2�+�R:���ٮ6���M��u�B��Yƍ��L'�ַ2�If�eD^n�k�J��OA�o��{�6���&v�PK�j	*�c�!�
�!����z�4��.:�X�PY����� �J��+�P_���)��J�y�@��������pJѻ��0DY$�Z[���#^���T7�L�����,��y�D���$�s���).ϩ~+������(�wJ������R���z�/��]='���"ra{$M�Ғ�I��Vy���`
�5>�x:[�k��V�K��,�$��E���vJ4J���vfG��M�}f�sa]�]�o;m��' }Tu����ַ��F���?Ӆ&�.�M�|*����3X��~��ţ�����i�0"{��Ļ���<�idS�7=��k[V�t��o�jKxn�v��gs�@0��Ժ������XA�S�}=Tρe�\����N=����*��	�Y��+-�I%ͲVz�<@5ﾹ�B�@��>�H���5�73^�Z/�1����S�'��Y��y�&����!�t�E�_���*vb�O���b�e�kH�.[��yxoM�{ހ�'9;�t�&p[�G�OZ.*����2о�5�U�-�y�g��Wf���=��]��!�5�DQ��?���)LR�Y����ׁ������a��.m9o0g���'
&�em�:~ŜI-�� c�d;B�����f����6�J�ŗi��+��&ٶG��h$aO4dc&U��A�`���Y�|"#�M��F��)&wno�L���_�>+ڹ����A:�N�)w�V�ݖ^����h���r�G���WC��\��޻FX7c�������ٖ�С��� �ZP��1�	zi��i���������h9��wu$�r�_��6���r�`I;�jI��2�&��h����=�Z�>�y�t�t`9����vV�����fv����=����7��Y���z2�O
��<��dN�}�}��$Zd�t��Ρ��'C�-���x$~��~�(�"gb��@h�M��߃�H#v��@�)}����VER)D�I�m�-�b����9�����a�Q��o畲Cxi׷���\f���������@"�)<�Ȃ�����W>�G[k��۪O�{+ʑ��U�tM�����[���(�IZ� �=��i��ؔC\owW%ʷ�f0�{��aԙ� 5ך!ث��uo�B���a/�Qz���*�z{�5�)z�Z��񉞯��ԍ�N%O��N��Wk�y�G�>����R��P��O�����ӨФj<.�FsRo%��Y��M*B%���0P�u��M���$�_7�����b��g�W�l���Ci��D+��q���B�^��
���?�2ppp�����:,��M!?h����Q;�'�̓u�&��4�в�ַ�kԘy��-�)x:��i���5(uYQ�X�k2�v`%�ay#6��u�Q�	��ud|c؋��9�NU��H���P T�%���ӽ��1����DӥS�pB�v�3Z�w�Ad�,�?Zl#���B��������.sS�$:��ʜJƫ�5��#��Q�Z�Ҁ=����'�I�`�$�%���3E�Yw�ݱ
C���^*�`�%li|��B�笹�(�۾�=})�%����1��N�ˮK��Ѹ��g���~sT���{���<ܛ��\W���  ��3�,h�;/Rbv�W�9�$Kc�����G�H������mT,>���,֩�^�ɰ3xW���j�Y���T;��c�]v�E��l�]��}
R���8��ҥ~�È7Ж�	2w7֧�g���.S/9	Y��#//�y���N)�o�M�Sl���G ���x5�~**�.�6�D������_�+FP�v��w��aFJ����E��!z�(S���5SI�>�44zۮ3/�,�b�DTsh��a��������zy�.��uW���̏$uB�B)jR��ƹ���Օ�\n�]��V���$�E��:����#�4�9������� ��(�f3�k�]Η:vp���67�j��!�[K3o�oB��x��[��x�p��$�Cd_q�����ս��$V�^n�ߵwk���H��y �d*����^-��J�w�����.�I�3��Ov��A�\U���	�S���u?y�;�uPGԔ���w|T��=��@*7�Ԯj���4����pz�a�8��4a.^̬IѾ����^=��ڋk�%	R>5��_"9�W��|�*��Ʊ�D��^D�ܿ�$���6E��>�J �R�h�I9����D��|O��J���߯��G���k{��;s�7ᮇ9e�F$�Q��}oM���]g
�1sv6�O]�t �/��d�	k����K��z+��5��3�)����s�w1ۏz"�ږߓ�Qs�w�>k�#z��m���w˝��G�f{��C\t�s���P֞�U\�8R>�{J<��`�NI�Ԧ�����л�)˥=bW*�mIܨ��:��<������z�֙�f4���64��Ub�$�"��:����h�+�9��N -�H��}3��
��FQV�T.���M�%�x���Ә�,�dt��ЦN����x�2�[/އ��7+(�z��b�����|yny�����q�Tg����tυ����Ͷ��-x�Z��[�T�^�P��,�-W����J=�N��F@���b���s��p�ߨNƸ���s`(�q�+��V"݈f���h����%x@�Q�iŞ�2n9���Ѽh���Q������mF:z	$@���ڄ�W8 ,v�c���"v#Àð���ϞV3�^&�h�Zڃ���k`�����;B�#k�E���bB �,�;ܙ)?�J��B=m��3ݔ
嬠9�_�:�{��̰����Gqy.Rz��bD W��zC*E�z��Q`Q����$�{.�
���8�>�&��=I�n�Vُ�֩�/%�
cYԳZ�l��^*��dC!ƀC��q���_넞eUr��բ�ͳ�-/G}��B	2�/�H��3T��?��3<��?�F��!�����9-���m~�-'ғ���t�'�vL \�,��t�;=���,E)���y�^�Z��Q$�T��ԉ�.`�CHi.�sE�g� ��~A*n�*4LY�BB��s��q}�H�*�
k*�&�m�L1s����fGu�"M����"�yҰ������<	k4�dq��o�E�ZtE�{']k�O���?ό�d0���4����!H��#c� ��TbQ�������c�ʎ���9ź�sȬ�򲕏�<̜�ZBh�-�����d�c�Qǟ�2)>���UQ�d��ۮV�Q
CN���t�}ݘ���?�o�*�{=G6���i8�رn\�Ͱ�T����Pq��T�������If�F�a�$2%�ןv�Hƥ8�SzX�y�����#���khn3
��;��w��f�:�Zw��
�?�[�}�l�4[~�#G���;��l��QE���8��Y䱑7����Z^�|������.2P�^��d����q��S��q���T�z�c�a�:ֈ�{�dI^nѵz>mb1�w{�8���t��\~�M�Q+/$rJ\`Z�"'��w�p<T9qY�` O���rma��	9&	 �)v&�Ą6.��خȭz�b�����I9zg����1�h��=ɒq6�7Z#w�` �.s0nE�t�ƃ$A�D۵H������@U��y���y��T���G�`$�2
�/���1���z�����V^/���k� ��q���ǭ�Ǭ�t4`�y���~MM��"�>�U�%������]6�7	�x�;��^�\7��*)���h�it�8�V�(=bt��kJ�.d� ���ǘ�{;���^�����|���]	�Fw?O#���F�H8v�����W���=Xt��6�vU>���:�E�m��|�M���$+L��GΊ~��?z�����`�гR�������9S�. +���P�UZK��8W���s\����c�*�q�+�����`_v����O�'�2C6,�l�.A���5j��v�:�{۬���$b��H���5'r�-z��LC�p)��ԱD����U�s{g��#�J��KL�E��h'1��v����}�oȐ����k����w@v�4x�
��� ���i���'ԟeа+�P:3j�#BB"��v}�$��xHsS�aw�f��)ھ�Hb�'�ɅI ����̢ޕ�&v4$��s�F*/#�!'af��I��_μ</Wb����b��EJ��o.�7}��N S�B�Y/����L�O����?�<�{�F��Kew�z�~?��s��,L�(�׈�u��L��尖j!��quĕ�0ZH*U�*L���deE�,�he$����/��͕��V���V�r�~�%f�.R��g��^���J�$ͮ��O���p��$e�6P�⃔ﴥ�?��98���6��Llu��db�6gbOl�Ķ��Ķ=����^��~�Uu�ݵ��������v�Sg�֟�c�+�~ꑿ�]�pR~~�c�Q��G����n�۞�%�W��Hn'!A��/�'ؿd|�ƺ���\L�{c��Ѵ�F�{�\4o��,�t)��Lg:�U�;ß����t��gU*�?WGOӪy�N�R���*%�(d�����S)�	`$|:iD�?=�?�L�Z�U'������W���>�ܰ�6�{^�I�_�a�֋�H'F��g�E�SѴ ,�N.��h�Jo����l�߱��S�#��a ⸇��UK��-��I$�=|3�5��׍R��L^n��h�)z�}�D-��fj��iJ�x��Y]�/���q�
�W��;��):���g�p\+�\u/G.�������R�&n~EB_:l�4�c�1L���U���W#��O����!�������D���Y�>M����Oڈ�H��c�f�S��o �>��Z���9+����#����Ym��Kw��-���rY+F:�^��F�`Um��ߴi/�)��%t���饓�Џ*r�s

����3���@:�}?��Sfo��c�P��1K�.!�n�]Xj��4�:��9��ȹ�P3�nZc���M�3Ǌ�a�0���v ���=s]M4b��h8Y$ƚ7�@&{��e8PW7J�i^�l@�<_�I��_��"1�[���\����񎨲i"zx�mt�f��au�+�8�|�w3�Rt�8���t��@A��#t�0c �u����)����T��h�h�ΔDK$c6����PQ�9��%����HucE�RְЩ���$W��Y���L��O�X�=�.�pR⑉���,�º#7M6]AHX����(��� ?�l��G����[ԉ�i��^<�����SF���}/T��	�[C�&J����B��&jr��i� ���vVy�wfU��$d��q����@<��͖��eB)��@W��f� ��U� W��� �pr��U��9�S��f�>^���UC�C-%�6�����>g?���?�����ҵ?ݒ��z(a�+��ؔ��U[��>���jWO4�R"��zGɩ�w���s��%0cv���,�9���N&W��{��Ȼ��y�!SE��h�sF�v���,��D�s�g�J����P� ��ٓ�~QǯTA_������?���9�؉�s� �E��v�S4�#k���6���c�����K,E����c2�c�gd���������yֺM� Y�a�0��%��(��Np}��.i՛��p��f��S$ձ�3m� �:��kq�ת��)ǓO~�F�'h�I$mOz���­�V.箝{v��Þ�E�8a�����t}}X��[��k
�Τ d�E�q������Ҹ��pr�܏"�D�3Yz[����#�e�_��v��y�$��ꈉ�K���{�,���d	��4���L@��+Sn�s���|�KRP��������66.���{ȃ�܂Z��r�'����r-"GxqtQ0�4�6���;�g_3����p�7�P8�x/-��&L�t��x|�~��(az�h���}�435|�k;'N�+}E}$�uL�J��lIC�����!j���)ţ�8]��)˩0����r�`q��U�-�}%�_Ծ�ʡH��`����kO*ذ̾z[n����Mga M�v_ R��1�$�!B�س�v!<H����z�k'�FMQ�9���&}���1QWV� Cym\�	�+Gsnjw�����F����v�A7��2�z�K,��L���K���2���1)iL�����G'�� �h��
,5�p�� ��D$	�϶c4q���I�d���s	�<�2��#S�"5��~kozȤO���-�ؐ��U�~uM�R�1�=��rB��R�������w�|diJ��f�#��5α���wE!���r���A{� ֡���7Z�<���+��w���#m�/_|qdu�}��Jd�.Q�sT�+~{�4d���x�e9pJ��˻��_Y��NM4ֆ��g���9��N����O�M��mڿ�!�1��������C�`�X �=!�h�v���A��&:�����=�>�(MNչ�X..Jq	עX|i���м�z�4�:��$DF�ޖ
�H7-���d��q����n�yY���H�p��۟`<���8��R�ʑSwK��T5���i���À�����b��S��n >!��O1��U��s�"8�zs� �9(uF�N=F1{�F�i�J����g�ٝѷ���P��'�[�B�u7��4�V�t{>�Fu8e�7l@z�R���M�w�m�@u����tM���λȱ���������tR�s�g�giW��y�[M�U^8��&��^� ]�j)���,����*;z�k_zlj�%�Ζ��NA`Tɺ�ug�T
�[ߏ0�3���ؽc0{��\�.`�,��u�L�:+ʟ7x
<�T�R�X��3��!����qj2S����4iW����zO����4<od"���?ގ)�}����_�ZRZ��´�zhy����g�mĹ�j�����f$���������A�%�Լc�I������?dt��H�9������k^8����Ȏb�ޜj��0�-NY���u�yQ(�պ0�\�Μc�	���(\�~[w��*�k�C�d�֨��D$&�n�9�-�m9�/�U�yY���v{x�I�o��C�ـ��eՔ��c���?��J�of��|bM�f��J|�C�Zb�fuQ�;Yl��Z��_ޥZ�Xj���c�.���쮮Пo�����i�
����3��8�pB
ޑvܫ�t�ǿ]цo�tڍg3����!2�̰	�����-h�\p��E�3�E�1e�6;-"5��.z62�ߤ	i0��2 �V*��^��FU��h�$d�֟
���'G�<�;OMG��r�|��s��H��d|Ya�Aʠ>��
�V�����ŭ�R�:㾱_��^�m�=	)~�ШC�CVJ|�w����IG�"U�s�=�:c�;�&k��%dT�V�q1��vz��qX��$���l �6Ͱ$߲�la�_Ȧ�~'FuqI�v݀�$U���*>z\µ{i��\t���f	���������J��+Z��VGfkR-"A�zHCm0MH�z���ҿ��j��+uמgz׸�<�]�hNe�rs�s�/�8�1�:���:m�y!E�� ��z����tr�&�L��-�~:���[.vкTQ~��gS�ѫH�`΢O�q�29��~;2�u�x2�<��-gBF�`Ӑ"��}T_W� eװimv����b�˗~�=`�Tg���fFpO�D���X��e.����9~�B�ik��
G��A?=�[���u�V���M���t�$=�QT'�}MS��}�9�,�:�p��b�e<�+�>y����T���Wx�E��9�6K���s)�^��ݣF��2nq��M�霞N������Û(Np�88��i�ovV�;Iz�@ު�xҨ9�%i��!�͘�ա�)���FA���%����e,XG5Z��;�(&����{-�)|�L���0K�$X����e�� �|��i�o?1��8ľ5T�M�������*X�%el����>_4]��!���D`���J�.!%��o�����ሱ~ZOS��9����K�n��t���=�W�JP��lA�k��bJ�NXLRv.�<sD�z���z�C�k��^ݖ��w�f��Oya��9���E�v�ʹ`�`BhI�EXPp�3�T��&%�NR��v.ݜPZV��,����X����||�y���B�n�։�� �dMy{�(�^���ד��_H@�]�mb%��}�];� ��}mEX*��Q��D'?L^���t�Ɨ�j��Id��_[�t��`W��1H�;�Ap�>W$��!e�^�sS���O��/�ÕR��0m������gǽ32��e�f�?;�}OLY�q���	��=����(�^���v@װE�m��	�-
V��\��Vw��&K����N4��_p��R`n�U��S_I7Nt؉	�������8$���!����7�#�y��f��C�qL���]�0hk�����Dc��vZD%����&���E�K�ؑJ������Zw����W�{�f�GaЍ�88�>��t
b�-���ղ���|���f��Tfa�Ur��ՊT��W�+O'�'�ݟ��5��7�Sðer*�N4�^�x�����' �r�as���X|*5�B�K�z�E��q��Eo�b׽t�cj[[[���v����z����ih-W@��;d�/s�o��s�k=��G��ґ��j[��Z�7�:a3U�Z�xqƻ?M�IZ)��`�Ꮞ�
j�(|��f?�Q�6�-���;XOU�����DB��G�^���N~�N��4��<�RT��,\3��9i�Е����72���]b���=�)H:��6~V��?�=<�9�ɿ
�-^��6�\�����`;����o���Q�@�<��B��x���f�Ja�W�������I:��)��t�����I��li�n���?�m�Te%���&,P$��3��"��ۖ2���m`�ҋ[�x���ν�6w�y7��Ja��cs_?A��7]f��(�s�{�-;vʴ�kր�O�O���|���o�R���e���S�F�2�7��b�^< ��o���}��Ĉ}*;��)PRM���/җ�����v�1������.���&��k�FX����FC�)1Oh$aJ��a�_��ix@�'=�����E����=�����l��"Q��~�����q��v�)����q6$`t;��������.�3��|g��$�{�	�g9�(��!$�J�ဿef�\���i���&�*_rl�w]�9���-�6�I>(�љ옎F9s8�Ay�>��~'kO�iL
����ʔ�u��/"
���;�"a�e;+x�Q��-�{���V�̉W�z�Q�u\��AW�{:�B�oC� ���iN���3)�k��ɼg8�͋�������.Y0�s�ϱ���#��c�Q�G]4��eR0	FQx���W� +kGcUL�����t�9	��i�W>��ع�������|D0�R4ȹ'Y�?�W������B��4#t��A��0�Ce���H�J�D�����n�bϱ'��H�F�_tN�`������Y��fȒҤD#Ét�d�����$�B�r8��)�j�k���B��}>q'E��5����Y7�zj��3��X́��l]�71��- %��Ĳ��uՌ�<�?���r���π1n�ND2��5hr.%e�2���[�$W�N�՘��{�zwj�е=,�ȝ�}n�<�uJ���/���Ӡfv�� Ik1	��i����E��J~�]�#�{���iI�L���k��$ɾ0�'o��'e�����3o�	�}~Z.%��%��B��"�F#,�v��k�n��H��@�d�
��M�-f��rӉ�e�C�����O�NN4��w�~�£�?�{�6�+��$��Z�*[O���0����C��}��?¬�*�B�@�dh�u��-*���8I!/<ӏ��H �ˈ��~�N0C8A[}�z϶+��O6(u����A���,����5�V�P���smVf/�����b�K�J�n�Κp8%6qR�Z��|:OA�A�4�"��h�o3���Yk��&Yy-��~<6 ����KF�j�|�r������n�:3>��b��)�w��Q9Jj�t�W����/d@����{bZ�?�4�1���$�I���d��E�vw���Nh#Ɨ�We-�}���݁�C62>R�SE�Tͻ��`{c��EѺ�p��*� ��R�Gv�BwA�&�Vf��k5	��5�����r�$�����bj�{a�q��/E7(Л� �i��8.��h�O����.g+���Sۥ���>� b8m���`�L<���V�6;�����{6_����ksx�)!ܨ��ϒ5�硶����<�2�����@<O�l�"�(�|�N������D-y���3�5��ޘ��˗!�6O���9r��$8��IQ���2� Q8rřft��5k���!���Q��cE�/�S֨�m����k����#�������Bvo$S+k̒�@�3{��F�U�A�p�"�s7qT
�$Fs$&�ǩ�4W΋�V�:�Ry���n��o��Qi�����z#��Q)��y��O�g�r̄���땗ULp�n�b7��WP)q��-`HI&$��j[J���Ƕ�~����Ǽ�\�ٷ�/O�=�it^���F��N=iuo��qF��m-~������M���M)ت�z�,�7�?����!�3 �����+j�I���y�o�>}|�+^���;.��h�I������n�z����*{�Cƽ�L7���uz߲)��t:��fj��K[O�s�02�C�p��"�O�P�Dݷ��3�Z��:{����-���f�10�[��R����F=Y|�jr�iEB���F-��óy��kA�� �?@���Cݯ�e��a�U>�^���+����/弓��W�U� �`ab�OFq�0S#\�R����*�L��A��Gl�bM4"�RJM"��XxP�c%9L�1{R�v���Ք�i��-&*�1��&Ė*���70@��}�O?>�V:ǣ�Hӛ/�O�]]�3O�N�����V(�Q�^^od���,��e�Y�4H�|���}�o*ʧ��	ہ����#%��M ��caH�m{�����Q�d�\��� 3Q]D�~�q+-Xj�T<y������~J���s"�?c�r��U?Sn�3��X�t�6�����^'��拃U�͗���,�Vq�db0�A$���9�F�x��+�=�gA�G��><E0q�R��1��ĥ�
_��>��PTG/���
�#�
)9���s[9V�}7��V�c��)B�H�@ t0��f�K��;�򥥹p���M7]03�g��5Lm֗�j�,��B5�0�4�gEg
H��c��^�f�c�>�i�`��6HU�*�a@�Gj7�E�3r��zS�<��ug/�K3���檄�!�>E?�?��O��E᮹Hz��t���g{tM��Y�z1e�H�r!�*t$F�m�-ޥ7�Ԑ�(VO��Î�}��[���2�*<T�^R� ãe|P�����K�����0�5�e^܎D�a}*-+	L�Z�,�
�=��J��i���?[Jv=̉:k=��KgdA{Iܮ�D����q��Y�t!^<ŒH ���I�IJJxЂ��}��Mo��~0�o���h���������M������`I�	<	`R�֣D xYH?�W�xBhR���`��Y!Ba*�-��k�CA܇7.�g�!�T��ր�g�ۨ�4�E�.0�X�0d37N�:^ļ��E8��'��P�[
��� �~a�on�,v(��k�ttCSW��,y�*/ڵ@I,jG��K&�0n�*��.
|�R���Y����7��'4"i�>����� ��ۋ;�7].�4:bW�;M{шC�d^ƏX S�vo�wf�X��ׁ��3���h����)�����8U�y�PB��Q�Ah?��j�����V]ʉ%+�
}$o��u/S~� �AkPF�3���2�]s/�����7ћ�EA�3�>��A�IH�`褪l��t��bM'�[m����K"������D�+/����y)��1�*�&���Ks�!��E_�`���tn&
c߀����o�kur�E��)Hr$�K�{G�����c�e���Qi�,��]�)#M_�n��P���5���(Eh�n|�][V[-�_B�¿�h�3�2��C�<��A��$QvSwh�H��C�'e����}K�� |SI8;�{J����<��~������j����w��XS�[�#1o� �?g�F�BC$^�o���$Ʒ�c7y�7�u�1�X2��B
Z�I�:;����	�
YR�-�ɔ"�J[q4� ��:.��Tzwj���>⡂����%඲�dd��H��J�9�N͉�]�,Q=��f�����%��Pe#�/��I�y�PCٹ0��jA�`4C��ް(,�D��lu�Gh�V��p�G»ߵ/�4c���������d�Fr��e��&�H!��15�U���:<�5��z̾? �i��-Y��B;\���BF�.�J��D;�zM99�!�Psu��a���_,	�B\��n;������M�/d�)�6Z(L���VƏ[�rV�b�>��)k ;�2�!Ӌ�h;Y��4����e�䄍�eD��j�tY7<��.�|m�8JGTe O!��JQSԟ���ۻV�kl��o{}���J?A���8<j��S92����m�Lo�U����<�'������6{NzL�C�䊛������8'&���u%�`q�	[DagWل��	�L��6sQu-d0�T/
ޢpd����=z� b��'�x�����`.Bp�B����&�?֌��@,��%C��Ic${� FE���O��(�d<�E������s�M�1��-4� ��	ϔ�A`s��]E�T�|��=f��]~fA�>h�u5B0��b-H����a��H�t^�{<҅u	K~	K!�����@37B��O���%G��bgTB'�&`��j_m4
B�9�%z�%��h�ؕˊ���M�c�����d�?�� z=1��/�<�6҆�JF�)���S+\F%w!$9���{�o��t��
e�;�*�
���`��L��yvM�K��+��O����
�KS�CE����6��olb��{9Q`�[$�H1��C��cp֋�&��GZe��6�} P�C��C>�:�>����#��hu�Ч	�V.��~�����YX#9S+��wqh+4�>���!�y�B
	m_ָ��B1�h�jeB�e���*Nx��qiD)IiB�4&5
�r�L�6����B̈rE����6H�Y3��4��JDH䊋���\�0ehT碍��`4� ��.v�#h�U��k�K;���(�7C$�+�A�gB�/��_��c�2���Rͧ�S�����xVpDۘO�#�X�"�����|�^�|3�c��J�&`�8��Kϐ�#��%�������J1D��u�����f�"�Wޟ���xS7<v�%�y�������e���`,�P�t鄽���P���D� ޤݏ$���/	����܇�|�=C����������v1�EFV�~n�A�>�]�}1��"1�b	Tn�to�V�Q1�*Gܣ�Ƣ�*�D�e�·R����p#|�PΟ��JQH[����.n�C�($�*Ҕ_-w�l���.���1M�����BԻY�h9mi��c�����ݑ��9���C',��<��:e���GrVr�~3�|Λ{���X�q� sU���8�&����<���~3����$)�5\�=���?����qʆ�UM�0��4�VϾ��$����R����ǟ��~a�W`�ehKR=�P�tN�d=)�R(�حd����B�v�������n�Α�f�=��H�zr��hSG܊��mú
G6u;��JA\��{!@��ʪW��i�Y���d��\���ࡇ����);�i/g�e����-)pd]�\������:w���?��u�Xo�jOa���3.�%Ԕ��n�"��y9���W/�mm7+$CL���1��y�a������L��9�Z��s&���*�wK����8�0���msΚ ]������2�n��9�H9�b7�쳺�r; ��-���� �?�F��B^0)B\��ю�	�`e_�w�C��y"{��`0Iu�ܟ�t��Vt��j��#�:�`�Hl�+��ʞ���(Ҡ�8h������^׭�&�/p)����l�V5�G#!mO����)�t��h�C���'���0,6d�M����h�v�;���-���'��]��l'��Z��:o 枏��}b��>��������ڶ�y�����;n$�Y���=pOKp_��8��/�t��f{Lz�+��+�]��X��z��e��S��0ʘ>�RH˾m�����Ρ��)�l�����&v����*a���r� '��S�'�0pIjإ�y�t�6JwI��[�ǲ�_�Z�"ղ�>�:���u��8��D>�%���T:�R��J��[����E	���J�[pd�d,����]~��Hd[���e�M�:�ݏx6Y0]gI�뗧c+��O���W.���2��"��H,#��C��*J�*:�-2�M�5?<�1ls0x�6h�1h�T�
X�X�JLV,� o�dJ�2 ���6)>b�u�5���&�Vȯ�Z�ܴ��}�z�ڳյ�~�IA�u���ک�����O�_Rߤ	��#�Щ4(�"�l���d���$�t�FQ���5,�SE@���Z��f/�J�Ib��ݳ'�4f�>���f��|a����I�LS�׺�-V�6��$h@i�"�.
%e���f*ޱ�}N�.!fB�� >����)�v�������87g+�6Y�b��7.J�i3+Rtm�C�����Oed0e9�U��Y�,��b���|�ׄ��%�咢�!�T�f����"��*�ί����C���v[h�"!S��顺j��Ìu�3��W��B6{/��MS���;+���2)m���YC��V {� @%Θ ���E�$괽�����xϘ�Nҵg�*��z~"({�^{2E����4p�%��q��^�o�[~�0i.#����š�/ަ
���k�Le3����;Li3yg�Վg>��y�+��օ��B{w�(E���_�O��n�[�駶f�*N��^�ܘg\���T�rr�����bl�/$`j��;�L�lQ��y8��(���B���d�^.f�5B�"�hH;�.hO����AX׈�l��Yv�^��c���]-_E��`�KP�$��ilw�D�AŮ�[�-/~\��ћo��He�P�9���t�JÛ�R��P�ѭjP$mj@;O0^����=�=ڲG %)c���S����v\pҊ��q3;/��'DR>����d�x'<%ă`��	�#� �H�4�<,H��!��c�р����j��߽[<����.�JBN��SJ8W�/H�S���̪�]A�lM���ꋿM�K�$�0c�Ն��x����� m�k}L�6߻ l�-� <!�D�r��0�>3��W��B/�u*�I�y��*�]V�&�$�E���&r�d��� '"�1Nbc+�ek��He�B��eVx��}��Aj���lz_�Q��[���k��}�9�y�b�C��jJ~u�A�t�p�V���W�=�j���Q�]��Ҵem��y�[�Ԯ�3M��yUl6���k��J���|=�@�	�V��d+��uZ	�f|_r:����z�4��/]�:5�g;��1�@~#�E��pn!RYEn���~ӵ��v҆�������j���P���Z��c���q����
�ZS��X�Գr��ʀ��<%�k([;���z��)$_A�>���x�~�`e�ا�����\����oY�4��m:��^C���~CJK$�}�RT��1�2-�S�s=�(H%���uZ��6�%q�Ud���"�ٓ�Q�E��UߦV>}e챤D���{�`��9�E(��]X����~א����c��mq9�����E�)qi��ׁ|�C:A|��<�)A+��Z(~�.P���m"�~�:�S��#R�P��5�o��b�\b&�ߙ\1��,�G�B��Cw=�0/#�07#���i��Gz:I�F��C�t���^s�c�T/�E	f�0�����w��dA�tC�e2���(������]&\���"�7
���M���g#_G� ��V{/�ԩ�0~I��=�����?��c���Z�$�2d37���L4�j�&�&�ޞ�ԮxL�b�
B�MEr�L��¡����v��:�j�(AޫI+6UO\_��w�3���(�sY�B�P���Q	͏��\ߌ��u>���- ���0t8�J�$i�5@�����m��jA��(]��Z�c�a�-�ULy^��h{����� �/�ޜ��T-#\�_y���c`w4��_m(%`Z9ZJG��C���R��&�W�N�����o��)�#B�����5�t��t�~�\�8}�����n<�z��	y*9��lo�)���h�
4Z"��J?���*��F}/'=���gO��L����-�!��Ŵ}<��C+@Y1~���L �J��Э�l��xK;���l �����й���c��C��*�l��϶��n96��0z�Fi��7��[���'�@z�J)Y&
���{S̟����Z�+ET�/x��y;N���x<�N9�����߷ܟލ(ʓ�[$ H,�P��L��B#qܽ�����b$�+M*�$ �F��bّ�Xq=3,�!�{��ĳ�M���-���~���6�(�^%�H`o�$ Jr��l~��r4��Bbv�kDr����?�'ꖤ�#����ab�6�{���@��٢����k���:0L^P��ĭ���B��a��])��B԰>.��K������������жp�t� �v������[�Qt����yO^�:c�|��נ�֯����?���y����>g�F��\�	"5Y*K����Ͳ�U�Z��w���7`�
q��k��K2C~�7��'�o�od��&����1�
O���:�Y��R��h�Ra�$�#w��N���S�L�)���ᛆ���-ֶ�+�$�_ޗ�\���ޜl�Ju��yd���o�׋�n+[��4��7��`6���V�/�Nb�y^L�d��Q=c71�&����5s��@���wekX�jz'��Ee/�������t��B��Ka�@�F-&��x�ړ�:���o5P����ݩ�����I��� 1P��Z)ayo���Ā��f{dT��E�GBk�+;^�7X���m-%�Rw��7k�<�)��J�/�I�h��F<|��������'2�ه� ^�K.�w2�|�[�M6���OFb��$�-��*q���h5��]�n��DyŽ��H�[�DWx�O�J�=8��~0�f�{�k���t,���\_��&\�=�m��N�y�_O�9��/��%Bt-�1�z@4��%	�ΓfJ�-Ω���̾8��V�Yǎ�?=��~� �X��[ntQ�k9:5�I��=���*�*�d�����u��X-���� Ϙ������n�db"��)�������O�{��B�C��Fg&���$�
��R�r��ұ���@����.�8[�;�zj���>��~��k@�|����r��E�21�����b���__B�h�6�P�#�h�p�)�`a���{�1�W�u�����[I�CC��{߸�Iɂ�T�\�Otܿ�zi�����L9������V�*��/�5P5�cT����~��U�d8��s^��B+N��i�ޑ=�Z4��	G�o�ll���Ռ�fT�nG1�u}����{�3�$MTzˋi�g��@�JNX�Ku*����[/A6�qZ(��g�*��I.;���=9ܡ>�;��%��O�Rx�����<ƆHl Y�Y�7,~)��ju糒��V�g��������<
=|���Y�Ga)7�1���x3����՛��؟^�m�YS�{N�>�9�C~�x���bT���� �%�n��q���ҁ5��nr8�}�z1�����U،���3]8�4��)��©xi�G�����W���13�;�P�Ǌtu�_�k_����t���������_PP��O�ӳd9Ck�UI�	6U~3:����*V�vs����K���F����55���̟ٙ�"')]s��q���v.�
�(��A�lӼ���K��b�']���E��ږn�\.�h��6���U�E��;���z��4����fi���a��ښ�����g D�O�$��ï�]�0RA �X�*��`�s.9r�N�t\�=}�h�����w1*�^W�f��<w{|��Λ]�,�\�b��-C�^����@���1�O�fCD�����g_´��]�9�ܼ���qm�ez��=�_#B�r�3�A~�|)�4�Qǩ��x���Onj1Gk�J�z_�Aj)<ı���zy�="M��C���z�U`]����&]�4(��ȭ�B�1�hb��X&������Sԍ�L$r��̯Ș�
)g;~O����!�r�>�����j����X���&bH����i*F�������K)�ˍb��"���H��HB��Yb��o�0�* ��?���x��s[}�%7O	�|'�0J�&f�D�A4|�w�	$Ī 85O��w�,�[�MGTo�f�B���)���hCe�:M�L��?7y!4Z̹�A4_��T}�l�V�lH�>!(�7�Z���~f7�2���4~����F��BxP�y[�󍱍��T�JX�/c�j���*n�Y
@���P�獥��E./N�[עM���d��0���LhK�}[�8�3�V�x$Y���g��C�hJ����(I�������@z+T��gb�8��"=]�i�d��l�i���V��B{�x���6�=-�]��='�=��MY� �Q��2N���'���n�dok�5)�:�zfM�]�+|W��AS�)d����b.L7֣��Sk���	����c�z?��^?&�J��>����)�+/d���ҴRex�B?�'-܇�t��)���d߼[�u�>=��D����f,�7<��	�x������W���%� 7�$�� Ɛ�^g�N����z�V�;C���-�IA�l�^Y��㪔��K0C��r�@+Ғ��S��R�/Z�A�!P98<�����p�]-��kKH���� (������
�_��<��<p�L^�أQ�b�C���%�V/�!���|�����R���?���!m,��ء��S��}a��ɂ���}��:��˕6Y\HP��c��G�t3a�娠�����z����Z:��s6�����F �����Ô�q %6��H���d��è�S �Y��]��	�~�����W�w�v	$v��O���� g��0�4uL�yl�/����RR�!x�jP�+�jW�z��Xv���֓Ja:i!�t���Y����S�D=p[�a��J��3�9wl,����q�e�B�R�JI���B��09"$�6�ڌv�aȵ���S<G���?MזGvd5
1��6ʹ������6�yF��B�������i�IWUB%���C7�/��a��l��.	s9Vqͧ�ݚy�����lt��;��u��s��H^'��� �3ϭ��lͨh�����ni��YS��B�z�^�'��\�D ���Y�%܃���{�n��m ~PΞ;��ED �ã���,z�hF����+i<�\۞4����A&01�i�rE;�� �Pl����5^�	����Ҏ�7�ݿ�'�3�1��д���ٗ�z�Ed�@炕|A=�b�>�;`����1����Rko�<rhs��5�₴���l��ެ��D.����e��;�gM����	R�o�f���v��r૓���߮"���7�֧0�
ɂn�=��K�$v�ϕQ'\���l��+3�dC��jNͯ��ӟ~����x$��c�wb.��c�w �����V|p@�7%L��{�o�����ե��3N �<��eIk�Zrc�R�x�ӻaer}|h^#���Ś�oW�gK��{-ǰ����a�E �'j��ͥI%b[�}r�S��w��^a���x��vo/�f���Z��{��=_6<����2�R�?:�!�����=��}�-�0#=?#cx���}O���n��V֩Yf�8K�J�޲�p-��8��px&^�{���o��-s]��x:�BPѩi�y��Kr���Ec)��
���%���m��M�6!5o��R���Y�-Ծ̮��@�Ya�ފޠbS�K}<�A�5�8��+�d��G����@E6��W6c���+�פ�$V���;C�����[_���ud��R�d;7`����09�}Jq8��讂����j���{�\f�<U}CrR�]�OLU���L�,hxM_����x�\�_�5�Nk~�ݽ 2���b�հ���J��s�����iO�,�.:�?�m�x���4�c�0u��փ������%�?ʛA�r{���Ұi���2�.�&]���J�$��7�0#��|Lci]�B���������������۾e�Vs�����ɂ�ߍ�?���x���LYm]8����/���N�R�u��m��^��#S�'��M�H�1,Z�d}���&���h ]���	�[�Rq��״P7V��҆EBY_y��S������$FU�Gb[��d i:�!��oK��I�[��2�C�#F�MF��_4�uT[M��C���S���C�Ž����݊S�@)���Z
%��;��{��k�5$s�����39��+}�x���F��I�����j�@]�p-���B��(.,�J��G^��b��<I�WL��B�s0w10�pI�#���g�x���a($0�i�p�y�p�Q��ki��*Fčl�>[�< ~�l��am"]6���Z2t-�0>�aK�ZF�l���&����bCT|�*Sv��&R4���z{j*��Y%V}�OPBd��~�9�3�D�Vm�떹�n����t ^*�d�S)�WP�E��@��>d��^�"�;���}W�&�'�:'�LJ���/E]w62��e�G*!�p�]��=�z�"ڔ}/f�˘΢�f!,�Ex,AuN��>F��[㼒J��ć�)4�J:�<�sTo���d�jfz�����ɷ��[��s�1ifќ͗>
=��DVա��ݫ%�Q�h+WC�;��⡖�g@�W>r2L���q4 v!���É�o1"�{`���k�D\*�e�w^\����������N��KbN�����j�����n5}�/e1�yÑb��x��arh���h)�)Xb�Y��dR��(�S*>nHv#I<m;� �W���O�΢��j6|���z�^��8`��"ށ܋�6�.��J��(�(q׹Β�e��WΟ�\��)�7.��\��ߋ@49���i����6e��M킵āJ�C�ՃI������<�ݳ����f�*h�@�S��I/!������e�{�k�?G��i?�.�  v�#�z8���1��
�/����"=��}�`�k6i7:ō��E5N�Tb١<�8�����c����cC����ٌ**]܀�8��S~��"�򮚋i�;�8�7��q���e׫���5l���:[	�_t���6�	u���)-d��Q�c��5ʍ�:~`���l5dp�2Z{pmo*�|�._՗{B��p�i�eG��G��[
�� &幭����.s�G����k�hS�zk���b�`� ��yl�,��K��3�!Ճ��[��c��Կ����}�c�xY�Ɣ�~aRtAG��0Z�����얕U����Q�٢�S�l"��2W��hn$X a��=�3�ҍ�)��nf��DN|Y]�UzВ�z�U�J1��mNT�M�!!��s1^�E,G��LR����NliIˍ��6/������*�1�0�h�{�{#g���M5ដ��a=H�q���eD�&J�VCa�)��E��j����>5�­;�6���L,u�R@����p����N�c��aX)��g�tq,��E��m��e�mx{����+������Ϳۖ��t�Φ(�WN�T��?n����;R�$�x�N?�}��eH�/Рڹ0SBt��jR+puM�S<�e�[gŻ3���r��k��3�Ծf��V��צ�"S���.���k����.b$�^\K���>V��0�|1?���^�z���.7eZr��nl�v�����F
$y�}�]���mqe^I9l�_9�;Y}�I�X�h{�����َ�ĭT~YPG���ě"�.~en{c��]�`
6gU�|��0�2T�	W�b�|�C���N����aР;�|m���.���ɷ��j��ao�e�����}V]덳�+�Ph�k6ʠ�+eA���-ߖ�#��>��,O���p F��'j�ۙ�o��B��!Q~��rW�� _I�C�����O�A�#e�&����Y��e���vm���M���>y�&5�~l#Ӛ����BP�S'
L)�����&G�Co[Ǣ�M(���l���u�l^�����5�1Z}Kt;\8������r�'$�+8�G�����|^&XX�H'?�GI��3N�t�z ���{�u��N��f�4��q�a:�t��.���\�)���`*���呀��ٚ ��oz��>ɾt�k������l��IdQq�Z��F)�a6������P�������m]�1Z�8��B��m�vқ�۔S	�{���}b���}��O��]%s.\)muI�}VN�#���3V�p�0�'�~&�ѽ(��g�����L��������U�KH�}����#c���矻���q.2��S�����[�Ou���w�����?纏��2�}��}^�P��9*r@�.Zp�"��� **0U�;�i]�H�`����˭x�8�f(���E,~�1/:|�ϰ�L���l}�eW���un�������
�&�@ѵ�dQ1W-�3��~� �ؓJG>��r��r���8��'U�j���fX^���a׏��^/w��a��Ϲ�R����\W9^�P�B}�J9���z�=�cn���mu���ua��v����x���x�~ ^}�l��?@|�E�Lsb|
k�r9����m}*�^�ǖ��/}wf�O�fh���}�i,pN�pE��FW:*Z�Ȏ�?0��3������R����+��*�P���x�u@Mt��GSw�Ż�X��ezK�1{��L�����I��x/db����K>n�e�_w����A�Z�7��n�.�	��Ov>�˧�K������n�_*�gU�����f�����
��ns��5��]���s=�v����P��y��V
T=4�Ϋ$53���� ��(��R)u6�h�Qy�nݼm��}����_�P��x�����Ͷ�T'��*�W��:NKWo�v	2��b�D����f��F�U)m�/ϼ�n�H''~5.��y�M��0S�?�m���c�g�
������̜��{��._l�v+�Rc��da�RԀ�a�������va �비�͟J!S�����[�"K��mo�F���	G��tc�±͢�ޯ�m4(A6ҙ���C�}krHè����^ �C��8��a*v.���ڐ���W��MK�W�w7����*�$�O�5�9P]w��=0��᪑D�;�8LY�Ӛ��S�sV�BÆ@zҙt���lI�G��mૼ���BK�Kp,B��Ê����4���)GO%��^��-���
�e���YۉE(\,u�m�`�N;jA�p.�����%��_����'��V�1�?��͉;�e_�P��I1��I�J��#�F�h
�I�AT�� x׏��Lj�������-��RD28+��/<C�<�Hz����l6�_\�!���'���Wq���U�v,��:�bL��Q)�#�\$�`f4��V��Q�s"� Y	0f]{�}Xj��9�M��k�0�L��2	� "kޥP2㟖�J��#zr,?l5�{9�A���z`��5qS�w�7hhX�%t"�|NU�,��B�Љg�^*��j.�C��\���vs�?_Shq������t�0�v���0������WP@YjS�x���0�^R(�R/̾��c�x� q~ַ�!����|�F���������E^����
�B������D�]%��R�����㒽+K����.�T{~�}ޏ;-��HL�<�_�4}W�'���1�4�\��p��)�	�s����&�h_}rT�^b	b��ŒZ����\M��=��������?�G�J��õAK�w��~+��8q楊����F�~뭀�`���Z����3�s��.�[�S��Y6Ӧ�������nA�9=O���av	�z�-t������e�Yn�w���;2O������\�@�Oh�/k�H���-����mH�Peb
/���y��섾��!��H6txEi�TA���r��g�f�W�}��ibiAl@m�����r��A�Z#G����������L�VF�iZjQ�HF�=τw����>�㋓�a�Ӹ�d�s���K'� l�jɨ�����s$��D�]��ڣ�p���M�:�&���d-�̦yy��Q/�w8���k�SX&��J�W�[�vaZ�'i8)�Y��N�ɩ��Y����:/�0������%$��m�=�DgF�y���$avY�~R:@C6ZF���J�OOX�@ِ�	���F�EF�&nlP���X���~8�!��P�%*�L���~	p::ߵ�Loa}�M�s���g��F
�ި��~1�?~�&����P��uvk����X����d�: v�b݁�S@W
�.|M2V����3N=��:�����h�?!�T���}� vm�z>.�q��R�J]��z���o,�,��j���W�d�����!�n�>pTZ�zl����Y���y���lu�"K�o4������3ѕ�|�[ vQ6�Z�va� �r��2O��,:���4�#$�@���$�̂����� ������?)��:���L<�\��9����W�ѕ�J(�k�]!����B����s�|��Nc%��0mG/�B_�q��u4����޿���h@j�� �WK��po:��G��9���w�R�N5l�4�8Tӑ9���F3���p���L�Ml�	�T���˚�� S���PǺL[JrH����㕘;{��w�O^�т���&�8�W�7S�D1��:~e�+>�t��d.�f~��H��a{p5!�%]b��ѽ1T�3�K����	�"i���b�δ輘����5iu��%��_�/m�o�/Х�(�>tٲ��	7� ��򩅤�|���/i�W>�f�kO�a֗�%<4��,��gv�W��!�5{y��j���pnɂ^�S��=c��u��!��i��{nv��9�|1n�;,���)1�Y<s���C��2l�Es��	���r:�	//��ְQ���m췵Y��g�Ǵ��T��Ƽл<LJ�A;��J���������A���u�>�f�οf��l`�{�ێc�ߘ��{}Yhism55zV�n.�7��|�u~��BQ%V����8#FQ�DN}�Ш'$��c���}f�u,L�xs�Ä�\��|bWn"tZ�W}ُ�'���b}ty�[3�j��q҄�n��^��vv�]�Q�e�ܺ�����T�?>��s�@e�i؂Ug[����&�Q@{��V��ߘ��b��G�Ž���n/���"�m�$K��W�Ü��&��KU��b��J�67��&��G�? �K:V�Ύ+�5�Bi���M=5D^!;�4���q�pHi5җqq�3n�����aQ����7k�ݝ�Ŀ�8_�K���y�[�*�T�
4���Y���%�0v�o��s��ɭ��IY ����2��ᚌ|q�9��o?�����]W@~Ea��D?�A	�t*Ȉ����Lr�)r�ºe ��x����o��V��S..�W~!�I?���wk{�=-���5��u�!�n>���h�]~n�\�p!Y�NǕ�Ax�m������r�0��lk�>��3Ԫ=� ���`��	�Ö�7�Ti��Ĳ�?n�8�w�>�2���;#Ж�m�d���c����8�n}ͻ{9�'��h�(��p:����Й���t��Şfc�!��S�x� ���3a�R���R��A�~᤭G������s˥j�[�����U,uD4w
e����,Z��������u�
���ڲ�H�V/wR:s����9����k�5jQHkuq#���O�]��.��Ωc���b�?-��V�����;H�����G��fŕ��u��ɼ�ߗ0�
6�Bj�$�3�dњ���F��ʟǣ6�N��?m!�Q�q)_�6FBz\�߆pI�cXaTM�=��@]l�fF��d�8����F
؄6���,\�J��YW�Q��O����m+��z�6�J��U��k��
|��T3ɛd%r���<ڂף�o��e����r{���B6{jJ߳��W��_�g����_���[�����B�W̎�9U�Sn�����i�t�(݉C�r�\�МΞOΟ�t?�o�ꍙ爉������lff��G_�٩Q>ܡEt�7�]�ZK�.�<}rcR�U�p�k��|՞����·Gg��O�u�|R.G�[�j�RY+:�Y�����H��͊��o�ɗ(�F:2����7Mt��QRR	�x�oA'��/l�ܔf���`uD��m�*�a}+��W���;3��v�>�9��9��"j�5w�WW]�
�J��Vx��Y��س��m%͛qujǤ�E`:?O��E��4��-{��>�\:�'U�����u�5�h
��~mP�=��h�v���!M���c4�+���	�R�)p�f��1MH�S�\ֿ�>O*�_�[��m*����hX��5�*��a ��=zv�ξHk;�B��㙩VVH'�E����u.�'I#���]�o��q��땀s
�ue�`q3+�����vs����9���	�mϴs���q��N
�!g�B�}�j8������ڽ����4�&s�R}�L���:�u�:f7D	2�sղ���^]��=��j[g��!���O�����*;�G�҂�}�Jۊ��1}��:��%Aa7�17��|��7Կ���SeЃ��4ء`�c�I�1�=����iW�^O��^����%.�����W)b	��o�8�t�Ed�k��$��n�l���Eb�����!g'.>B9/��^�3{S�˾���{���S��Dሉ^���@����mQH�_=��s�J�c�����ۛN5Ń�
"i�O�ؔ�������������H!oTa��/h�kv3��!r|{W�|����_���n�/~bs�q��Ω�z�ʺGj��D�5��І� :r���^��Y���O��Z�+<��s��J"��,��m�NL�zY4�Oc��j!��^��,��N׻��`-z"u$;�\B�]�ԋ��t��K�O�±�mnP���O��0n�=�M2�{v�.A7qRx4�Q�����GIF�i6���P�^_0R>l�ݙT�i	:l�������;��9j\\q�L�<�E�OҨ&rU\Y'I�н �K7����;C8/��®F��bK���@@UC�b'�\6 QN4O�`udс�S�=��۲h���2�e�C�!���ק���L��<cr���4c��;g��lz�8�53�EO������4qZ.�I���{ ������*�qFu��)r$��e�~ O���Cu�\����������n��s�=���!�9Ͽۿ��8��U��r��R'�,�P%��gN�Y��µK�TM 5LkNXj�=�.o����H��s��I�y����	�Ux��z�}+ٿ�`%�WuR����q�g
�����rf�#�F�ͱ��x���CH����|�@�)�Nƫ'���q��~�ȴ^8� ���_�L�"b�su'�N�p�wT����/���b;�5�c�X��B"qok�9��I4��C�jP���r5��h�8xt @�/�K:���j��sUw|w�7; vۤ�$��A��I/�:���>�*z1 b��D��Y�jc�s���8�����9,笕��@�!��G��ߝ��0�OH7C������
b��`������0�H�9J��5�^Ȥ*=�����wZ���i#�����K�p�⪄��Jlv�����������������d�2��0f��w}�ܴb��{�B�s�j�ھ��l;�o�[S�4;�P�������/)�nNe��lQh)�U$�t�ޕ��vS�#�̫���j��G���Y�f&�YZsbQ܇Z��ĥ�Vw�^�Ah��F��q3��Ĵ�`���U�a��@��E�s�lkc-��	�p�����vKT�ܟ�|G8y�R���d}��������4ʑÚ*�kܯ��6=G4W���zɳs���|�.t�������X��d��R4-j֙���k.�dW�F���^*����Q�o����x#r�Sv;��8O���l�^��"=��;�^`�9�w�im��u�P�9�@@�u�׈�@�Ǡ_����C��0UM_,Ζ*�檳�����{ʍ �UNie�H��2�NS�C%F��fLp`NxB�{q��|�ѱ4� �:��TL\�f}ΖѠNX��i^a�/��=�X���E*�� ���R���|*��<e�������=
g��6i�,����r?���y=�bLׇx�'���}�����xYB��W���.�H�ٹ�:���i��ŵ�Ž��3-�Q�1_�N�Ѿ	c����B�j)ڃj����?�;�S]����u�
�~���E�h	�){��f�Z�n�����R�" .I�!���n��9��&�ר��\�X��q��h� �O�롢�x�[�f&)ճ_��h�rJe��V�$=�7~̎V\�U�e��*^NZ(�X��g��<� :����k���ة�n0
m�C��u��q%=z������S	�c�'���.�7�	|�\�`����i�m\&��>
�'f��]�3���"�[����A��2�����?�Uo/�����z��X{|f�>��6�{�r�{��v\����l�?U��M>L$Js��!�D����I��ҳٕ��݀Ggzq�3���f�B�1�(���j��*` ;��6���G�S�7�M�6>���$-���?���9]����h���m�H�C��L����*��ƃT�=%h�3��l�KD���j��+XQ+!|�u�tV�R^��UoN�TRaIԉ-%o0g�{�Ic���_O#��b��
�@�aӉ�b�jn T���k�O�?7�c.}�\6H���P�-���ڙ؊4?ɐ�ډ�T�8f�nDV{��a�v�$W|�͸Y~��r���YDp�.7uuN�3�*v���V^�t���S3�^�ُ����)_��M�DrÌ�Q��M4�u��u�k�`Lк+_!:��;:��3�v09��u�sRq��Vfh��ϢWЗ�H��k_J���O�5_��9��٣4�J��OQ�C��1Z��ff��Rg;[�+&�z"���K/g���������n�����w�B��w�R�i	�W7���p�2�����:\��Ϩ6���^.M]�Cm��s'�C/3�P���EJ,�J�]�JI�Uw����^JM뇰)����c�i�}hP׮i����]����g�����YW��vYe��6'^hUkT�MN� IK�t̷�=������v_��h(��qR̊8�����v��棘�)ux��nn�Q�&Dz�s7l�U��4ѐ��(N�Sus�}_'�ڝ(J����Ņ�>�%C�� D ����� @[�V�Z��Yn�G�+b�wNъ���>��4T������'�P@�Wq�#��@�Ć��mK�K�nL�C)�./1��ˀ�0����D��+�l���V���՞J��[H"��0�X���3A���J�2���%2�����X\�4�n��Yq c^�O��T��*���h�[kBn��Z��C
��V�*��E��r�%�����Ut�\T<r��"��N*ƫ���d�����2}6���&����^�L��~]��W~r�
;���t~t�Ź�7Z�n��X=��M����X����/�"1Ο ��P��A5LoXw<У��B\a��үy�P���I�+�����@e�z��-��y!��N��ۍ$Pu|�X!����s�G�;+�ȋ����բ��畏>6���.rw�|c>@>�J�Ɛ��d��BD�;5��GZ��� vR���P����>��^���Ӱs8���@Q_h��|�K�m+�[����}���b�/<S���T����A<f%n�_5��kwk�H]v̘+_�n��j�^_~�ĿaK-e�g� Pc��F�l����l�Y2|@u��q���<㗊y�>�3|4�ߦk�>@�dz1j��U���Ӭ���A�[R5��%�O+H��-�H]�vYS=26v�1g��P�[5�xM%�\^n^�}w��n��?`�\*�����]���hT�w�xk��	�w�-R��Y�m��q��n�]H�s;��U	���*Q���j�ʤ���c�sވW$���t�h��|[��p)
��R�2Z�/�A��ű����	�
�?v޿RL±�r�,�( /J�C,�&G#���gƞ��ƾ��|���a^2�j)�g�Cyv)�{Y#	��Ӏ�OJd���
}�XA�������J��-��F��>Xϴ����}y�zKuD��d�
ڸ� {wm�~�e�*a��h�[�7+��hWf�bxܴ0�����MG�����Ϧ@:ؼ��=zjx�D:whZW����64�Qn)BGOpA��?��܇XAΥkA��D�����ѧ�43���!�Ѻ�*+p%�)���]Z�kx�a*�R�� eǍ��ʷ]����ϏU�z3fơ����!����(�YO����`�Ci���$G�3�b�<���N�2��]7����C_O,�t���������%2�����pP��а�ˉ[�ְ��qB�9FU��Q��I�ShV�,��E\� Έ����-���Z��-PTp\�����G��#6�~����IWQ�{���uy�[��������?�Κ������h��d,�	���^���zFV/ei�^�ݧ6�-	�؋��xG��B⢳X�9���}�κ��O����n��:U�g1��X_�RR���bCI���F�_jr��O�R��;=�BX+!��b�N��v�5�֟tJj�q������`��@仌-g!�k���6�C��UW�	!IT) ��{cFm�!U�ʉ��� �_y��" Q���t�s \Ȁ@@�$�3��d{de!����|�Ԫ�(��;\�2��"{�H�d'�b:��	�Ȕ���Q2����[$a���A�)	�1���tx�E���=Փo������<E0����,�?���>R��n�p�CS��T��}����aZj|]����=Y2�߾확���3�
K�"�,b�7ծ�+����Ӥ��Y�]�xV+�+F+Sk\E�b�v�,-3�I%�z����a3*1��/'zn�
�h4�F�� 8�*�5��.ۭ�����	9��$se��G���;��1(D�iQ����00]�hξ���J%�?�5軁y �.e�LR�B���ϼJ�����]{�R���p ~�=�e��½��TÛ$5*�x>��AGG2蛦m�FY�wQ��̣�5՗F�����8ϒ{a�(��rlR}3����f��Js��}Y2�:�#^��Y�s������c�s��rw���f��4�	<�)**+MyI?��Ք�F��'욿��,h3�O��y�����xI1�� ?p�6�e55���<1��?�+U�<>&&&�x{˹�p��8�1����V������8*f%�#ebl�$҈�l?�~�#�RG�K����3�``���>������]�DRo:��%1���ަ��5�[��������b�d\��c�1��լ����pf��A��B���k3I��2Y��}~�s{J�i��JK�g_��pN�/�$8�8��g!�_Z_W��k�DI��w�HM6��2����&�p�J��L�A� ��
r�6Z��iJ;GԤMG�DW�@W�I����TCEE���V�ؘ2��ǟ������n	DL��o�r4���_^��͉����~K4v�DI-�����a�z��W�U���݀
�GN�TU	�o,�ۯz�9p�����̡<5��$>�����8�����Dґi��k��I>��?�ԋ�k��X�Bo����}%��
�~�Sd�ؼ)7�;(����.,y���
�!�b���EVZ��Y>�r��zW�B�/O��j���2�[hJ��*���}7prb�w^���# xz~�rݒV��1N������iQ�^��]0���>/e��k�U�B�K�� %7�O����|-9A�^{Դ+��&D�6Q��R�����*�aN]�vz���/&s�����gD�������M��~އ�ʨ���c��P�aT�t��t\�����ém �׵��ޭ�jr7��v�����G�08��i�PY}��ˤ�2�ۙ')��_HHH��
c�J���H9O����_�Fo���#����=Q�&}Şh��Qk��յB{�����,�|ʵ��r�I8��%P�/iH+�3���Qi��2��9m�tq��s�@��$�BS"��E 7N���:W'�82H���E��w���ۅA��g�.���T��i��k��M�R�����M}eS 3�<q&�QKmGhOϧ���Յ:��`(Xhu6�ILl�����y�EbRĎ�l����k�wW���!��C�p7Q���nLR��퇠�z\v�&��'���xr�~����/�1�å/o�^�M��z����C��/P�i�*��"nO��k� w!f`'�~N��8�WbZ"���/p
����_�&f$ .xI���Ҁ	R*�z�y���$�W�Й3
(����V�}}�`�}s<��3�ʟ�8E'���yxx���B���8�/F��q�����T�W�"s��	�&ʝT���npe�U@}���[nW���/�+.�]g��Iu?��n,�j\B�����ޭ�:H��>qad놊��_J2l��S�|�g� �C}��\5񕒊_(��i{����iJ���r��1�/����w���6�����Yw�J�󆅪Fl�0'�tͩox�<�p�a�"XR�ߌjvv���|qZ�u�b-��7�ec���OG>�^s�#|��l\�=�K1����'P�;{����싾m�)��ҏ�L���7�,�p�4hs�)�w_��2�yT���:��bg+��TN���6je��p=�9d��ݐ}�L�e���ƛ�q��m�[�'vH��e��J?���o��'4�l��@���M��k��o������5�lb�����`jZ�\��#�Y�*-�ؗz�{�������a৛������
�s�u3PT��!�^�sV��S��|xb(8�����uF���z�׳����Vy�0[��,*�0�KU���k�'�����@FK���/Bz�9��,�x7�1�|�����D�}T��f��/p�u< V��BG�C���.��*�����\�~������H�R�����Ǹ�|v�l��[a�+�vԓ�y"��~�[9+��x�=rD����[����eȶӆ2�����F�R���\����FN�q���C��_��`��?�g�\�Pc0,��dMo�|�SoF�s��o6|/��=�ӢX�2pU~�Cg�!A�h-�="�/�E
�&��^���i�BLL
rRyh���z��qx�T��j�"M6�r�P�t|E&X\&H���j�Xh���9l��a��EQ,p@jt�c����ݓ�"��E�]�'��My$˦cb���؂�?p��yc+�b���M6D�̱S������U|��kͭ�f�����`Ouw���xFώ��[��'��1�"�I͠Z���!��Ih���p2-UJ�M�����	�3~�@Zx
.{��&@�;&-�OѩB�O���b���&�`���ϯ9shMv�gɇ�������-Ҍ�R���Dx�P�9���h����vͨ�˱����A(�S�Ѡc8���Nޖ��n=�'���� �@}�U�F�<�x.Ϫ��K9(Ȕ0��hpE�F�哛xg��DX��Q�\�g���[2u�E�d	/`}Az���&xL��H��@Z¤E�A��=�8�a{���^�;���G����l�+`/�*ܶ	+�+�����J�T��\��nUZ���=��<M����!�}I�o ��
4@�82DS�K��G���X�	>}����H��#J	2���D[�oH�Z˔R��l��j�|.@�����&����i�0X'wR��S�n�Ř���#J�0��7)j�;�F�?rA��JJ_����	�J��������h���w'���Rq�~�n���r����T ����"�CǁK�^�چr�Z�v�(�x��poS�{���qv%��� 
��;�
��p��?k�y�1}zJ�>��ĶEO�\gg���{�+v&"Rݢ�gRZ���
;�}�Jl!�z���"w���A��F:�?��භ���lp��l��"�Q��޿�賮�vuM���Ц���<�<B�:�ȏf\=�ɫ���㨱/z��Xk^��`��L�<���ᡭ���`:K��|�L�+�<��ּ��ޱl>�5㕕Zܩ���6�:f�S��\հa-�T&�Q�IO.��c�M'IE/>z����5�D^��KU %H-<��,��~�▁p�����0���`����&�6 �f��q���Ϗ��Pٱ���e��A8XO���u�,��%�C���?�ڊ�j��c�	f���d<<�j,�Τ�(�g�%�\�` ʴ5��.�� 	��]A�����Gȹ�A5�D��Bx�\�A)$͏��!���6Ŀ�Jm�v$����kL��Ԏ8t+ǐ��w'�_����z��د������� JEzxH#�/�ِ�ڭ�}��8�{���+71�͛��A�,�x��H��{D�FK�9o��햨Ԫ=`���Rcc�-��_�m�$��2)�O���gQ����PH�
��+<6� @��z�~
)�W�Z��էZj�ɬ��vX�!ݭ�%<�Vv`�kJi�/�����W@�ɗ��E���75�/���-�!ôھ��Ԫ��:%�T�eg%I�8�oZ]��0�dU�Kr���m��Q�B	�嬰&�g���5k�,⟁���b�q7�\K)���3���F��5�p���Z61�5�ҭ�N����o"������J>���(�x�H:8 �I�������qg����՟�۟��	��u:�7\8m+���X�z@�>���&߆��c_^��r�-����"�]��}8�ȏpP�5"m��񝵩���(P��,�e���L��"�p�W{�JeO����������6ר}�K:NpSyN�(�5c�������o�>����Ue'm�+ܙΟ]&$Uq�#	t_�M|,�Oe$2an��n�jy�-�	T�����k?o�.��[�M�%Q��Hz��d���E@#�^XG���Nj�g��R��w�y��߳ ������⼝�����D4f��#��T rzN��v��@��yU�����{,1Ax�<P���f��qN�;��I���?�q��H���ߒ���
� 6 ��\�e
��W�4 ��`��]L�.�|�"�Ɓ��v=�d���ҙ�	�g��p�ނ'�.�w����Gmt�y�r&���3E�̅vq!O*�89)��tGF1ubhh����vѠ�)b��;>��e՟�>���l�9����(c��~�
����+vD71��a^���wy��a�םg�j �1��� &D�\u�M�w�������m�Y�ˬ�'�?{S�llDd/��+�'ܩ#;��>����2͋
���C_���z3S ǵ�uu? ���
�4b������Ҋ?�N��լc�uե\�����^�����&BF��V�2���r4 ��4���pִ��ESR&+A��D+˛���Y��_)��-�����$��x�2��H����ްH�E�)��r���)�P�e��F4�eh���,���ޞ�;ǊᲬ�G��^d����$:OS=�}����o�B�Q�l� y �����|�a�G��{3n��%�9��Ů���6m{a��[��X8�r�x��&8�_P:ۨ^v��gMӂ���}�jݹ���T�ݭ��������4�x��:�$%L_��D�&�}�j�32��Q��p=h5�3��owT����>��/�_�J���b�;B�F�by����7������%[AtBDMU�`.�Sk%o2��I����R�7'���ݎ��"^aP0YsZ7l�M��_���%���I�f��e��]i�ͧU�$�ͧ7�ǥ�/��{Usx�{1��P�׌>!Ӣ�B�f|^)څ	�~��ۢ!Z��o�&<��U&_-uK�8]!Q֞��R���ι`��t-�I��u:fd��6q�s?��H���[��>�:�ms��������m���-Ag��ؔVԫ��)�l^[����L1�悉Xo,a���#���N��O�@��t�7.���F����Z+a�G�#�q�٨�L
�z�]ٻ"&^����X�	c=����%�W�Q�?��4�&1��,sL��r?�P�������g��CY,u/��U�5_O�ڴ�u�l�g������5	�lk��mb���W�}8mES����j�VQYIJP
Kr��21o�wL����tYi���qb�CL����8JyH��:Y��R3� ʖ�`�i7��~�^����Q<b3�<��kYE�h�	�=˗F2-β��I�:�^�~{�f}��<���i�H@�����=��P@�[9�%	�}������d�/a��Q3.	�mBl�z�p��b�������.k_qq��6t��Ņ���&GE�'OV�������P>i�~dD�����4[�*�S�D��2��LR��a˩�ʛ6�A�H�?Q�cQ�b�q�+2�o�Qh�*ueXVa��2nû��_�B��0�ws099�k�Gt*���T���Y4� ���DJ��2b�D��G,�1U��yRr�U�8�(>�u��D^����+���޷	鐒����KR��[�sD@�N����FA���|����ŧY�3{�qŽ����IY'��y�C�!~2{;��3G��ۉg� T6��c�j6���S)�㘧�;�a��^R��u�,Iǽ�C����mZV�<�Ř�L�G�u� Xeͅx�Ow���v\5��^�qU�~S��1G���A��J�_ߥ�"��P��.Ӿq�^�`<���c���5�R
8���	������&��?��{�;}��P�K/M���ͷ����CK�o8ȍ�6������Jr�h#�z5���Dd2[�ђ�>&4ñ �7�Qhv0�eaz�a1��~}$��܉°����Ypܻ�rN��[9(aY�gPG��͔ +��4���r��,N��9|%,/ ����׵��2���!A�˓�F�*M����PTIQA��c�V9��(��Ū"h�ip��R����\����L��v��&u��K���K�=�}����BG]�^���wsvxs�TӶ����Dh�#����	H�^��r�W�~5s�k݂��d�6��ڷ�V��D��]��_�0��^?
8�5Ċ��St��NZ0X2�,�GI�u���;����ak��b��0P�՛�$�)'�y�\��_A�[��oKK	���W}p���J N�⁻֢I�3��Mx�� "��st�,ۻw�@�3�=���,��	�;��wsZ3HP�8���Zo纆�j9x�}�{���T��ų�,?��&{�4���y7���n��6c����h-aH�7�4�]��Kj�͉^^I�4�S������	�1L,sT�xL�>d�F���Y�'����J$b��،�F70[պ�r_��
(c�����2�X��Ԇ�.�o�Ћj��ω#>>7ç	y����R���>�0;o�P�UWw-w�wQ��ۧ�q��}�j/����p��tM�IsI����Т��$�K�?a)Ҳ���{~�oԼ�tKDw�PK"~�[k���=�K����we'��&X�MG�\�5�_�@�˗�&��E�>�Ŀ0�$A8��9@4�B��9m<�~o��9@[��L�}1!o8Q�[�M�w�!��T�l/� �����p��#��8JRs���o�;"�\��	��g��c�a��m���J�����p񨺚�u��Q ���/(2э}{�;2����^�3w�����u %{�Q���%=�)g'�h����f���a@�p�q,�YwOͰT@�&��s�eag��b��9W��#���'�O�##Q��Ձ�*�G��p�o���N�*��p�î=>T/� ]��ݳ9�n��?0ͨ���O'7���}1BC��
��K�4L��V��Xۆk �M�Ҏ�~��v�
�"�����M�6S���?exS1:M�a%��^�!Ȱ��ي�Η�Ib�c;����˫�n�;
,���5��8|d��X̢S�7P����f����L럞:MJ��W�i�ϻ���F�������zB�d��u�)Er�}��mT\C����
�E�dE��M�jUď'kmE`�%MD]oQ��"�$��f��m��Jd�Lёe[i� �����E����m���+]ղ�wTw����=%�)�í��O���������Dǉ�������M�"՛su���n�T��C��ȓN� ���n�?E�O�GW0E���hh;�-���++�||{��E���Ba�V�~����Mp�6�s�Bї��%��貫&��q3(au����\�yŗ3�7(� 7V"�ۀ��f��I�~�M����,��>�	�ϔ$�9�u
\��`�ܖ�b��Lo�E7ܒ�����_��9ңL='4e�o�LX��)�w/���l�PhԂ�fkNܓ>{ġd�$�qzj��<�?�Y�5?9�X��M+�a��F^�Bdhs�mP����� w��/��4��D���I�l���L�#fΉDD'�� ��X)y��>���%��kݭ����+J<T���9�D-8+�d�����V�������w��n��Df�����]��ח?L]
I���1 ?��$߬^X{+Vh�c��H^R�8���A,h��K��5�� ����y�	n6�JJʫ��%�;�B�vTC�京����e���p?��"3
����Y����f����V���x� u>@��-Y�֕�����z2m�y�.���Z�
74k��I�7����� ��ԁ9Z�]���eԚ_�����U�B���V2i�?�ԣK���x���8Ǆ/�h�K\8��T��?L�&.�|�.��#�[���}��R*+�ťϽ�;l"]wb��#��[�{��4�'�@��=����ݐ���n�m��^@��EN�W��	�/��v�D�Q�F+;Jt792�g�.��{)��њp$EsJ���qb�=z'%�((�}n��8����Ѳ���ă�-�>���}Oь[k"k�+�����IBExV��GND�ql˳�� �0K��)4q�܉�YKQ�×�{�a{B�٭�\�g���Õ��8u�gA���i�S���������(�y�xݕ�m�Y�W�|�$G��ʻ_@�������2��+D�^��E[�[�؄�{٬�д�u{�:��gB��X;W�C����T�k}����>X���
DW_���	�­�$���l�J���
����5%�&���%��~Z�����c�?;Y�ԭy����V��蹰�Y��98|��Z�&՛��VZ���S5s�zm�Bg�J�2�B�'��A�WT[�D�'M/��r�g֎��"A�K�k�sl+$bi8n� 툉V�'iE��C���S�J����bwC�߽4+���H�unO�R�C�/IZ_��d1�\꩟N�΃��i���wX��������U�h~K35_e��ut��/1O�͡�8O~љ\�s\h�0)6��,}���4��'ҏ3@�?�E(pa!�(��'�s�Q��χ�ua�ݯ��n�N�tw+*+�Zc������}O�t�S����']����C��%�ӫ�/ME�͊#�b��*g�|��o��#�'�ఱ� e��۱�4bO~�4;G�F��O���t�^Y��P�Ln� ��i�堹�6a|Y��-�Ʋ4��sw�ɋ�e�7��'L�%B�k&Q�>ol� $�0���z��陿z�-!�2�&��L���B��W�� ��W���o	�""uV�1�A7;���8��b'.�=����8b�sz���m6侮oom��=)���f[�e�e`sw�S9 ��Ê��М���u����1[�]�ւ�@Z0TL�2��١�$��f3K��0��ؾ;���G��$8zc���`��9V�OG	1a�~k/�L�8��jYK��Y��k����?�C�7�A�/W�OztHȡ��������6q2�״�r����g�t@(>r��G,χ�Ys�h>7*�I�}�D�ު�!R��s���{��:W�
3���h�����n�E�1����tJ0Ӫy(�5ƽ��.XV��$�1Z�"�����srf���6Z��>��;�:ev}[-�J��(gޖz]�����k��ܰ/���)~<л{���5HBA���EN���Ǽ�y ��	�ռJZS�N{���_EFO	�Uu5v�s/s��C��?��t�=Q�����0��yc����;;n\h��#8�E��`�u+���m�W��NM�~b��f���~��ܑ������%ߌ��dJ���h
*�˳e��٩r�č2�v޸�Q�Je����*쫐�䲇PzWWT�{�sG�I�P��e3?F��� �!�:���&YU��%���<s	����9dܑ(�!:{)����Wpb��8��s�-�m��E\e�C��#4{����_���rn�$m^�Q�Y���4?Q���*g�����)�XO�ھ�}����['����q,\M�no_>w�LS� ������Y��٬�i擙F��_	"7�sq "J����{�G_�����'���"Ia�i��z�y�Y�VX&,!�����P����B<���H��,+���ѴјE.�]��p���MŗEt�p�gA��^�aKk�U&�g�e��b�gv��,���+�D"rd��h�����w�.�/���$��>+g���߯����y�~��w�����x�$��;k�����i���?��'��	ߤ@ϛ$g���Dp��e4��)88�i��pY[B��B����f��MԄA�Ч{:���h��88���`��^������Q�L�����7�G���r�f8���}�xR74��Q�ϕ�R��j��P�K��[°�;�EM�뗖l�������B�Ҹ� �ʿ�j��4J!���2�Y!�ɵȺ��̽F[�<7٭gr8*a���*;�y^9�a2	�ry����/j�ܟ�6�5�v~=F�2�٧��3-�!V�cˈ��m��n}f�2�Ի�(Ki2��k(�5�a��*���=_�.���Hl19�cэ�:T�|�k~(?��YOЅ�a�r��y�<IA�eϹq���g��}�舃����:�kSu�TK�{�+��v��f�h�����BOp+�k��t�c��<Rܗ
n��Ow�onin�|4}�C8[��JOC�x�7ir=t{4�O�sV	: ֟���[�?��j��z/����ɓ���������J��W)����a��.�ֻa\�>1ųQ����2��\L.��l��#?�MNuG8.f
�:"2B�X\����ϗY�-�����:��Wՙ���V!\���&f��iI�#j�}5��^l	�/�O����M���,^ٜ��pN	;�6�E����&9���ύ(���c�a �j���>+�KvZJ��b2%&>�f�1SĹ���	�І����
x��=8�7���Kﯓ�� ��E���i���,~�D��P� я�*�s�'0�g>ƅ�c�/����}(o$����� �8�4���]��>�U"�-�ԟ���ۙ����ӎ ՛��3V%�g����<J]N�T�B�h�Ui�F�<�`]e2���R7�%�|V���W��˖���iԼ��ׇ\��qok�Ik�(w�Wdll�)�$%_z&Q�t��Jiӛ� �;g�S��(��#L���	��/�{Գ������ӥB��������u8������-���^�LB�ʝ�b��n5Ds�d}})X�E8�
e��ʰ�g�Z�|���G�SS�ۭ����e��=5]M��9�(?�(0¾�\����.��wa����^_�ؕ^�a�q��4%=�w�eM�}Y[��z�:?oul�󅃛ڂ�S9�#c�P~�.��|]�c�O�Hy9��ן,����.}��7$���1��~��Vi,-{��w[��#gW�W��n=�GIy,�+l�D�ou��j��|�e��G�o��~^�m�+�N����!�q6ێ�642HuKC�z�����f���w���9dȿ���:H�W�Hzh
���[�s@���Gz䰲,����^��3(����e�t��9�ߋ|���c	HK{��20ң������d�����.�D�V��h�?�!�z�rD�z�y�C���@�k������%��K!���ˏ��Q��o����$K1�I^�m�1W��)�U��T�;Sd���mrPKNq;W��*��:C���u��-����R�FIJ�~HIq�#��h,�Fl|��Ҝ�k��İ��o�M�ܸ����V�c>�~AR�P;K@ Y��N�?���;��?,+$��`5��+����4m�^�j2�N8d/��om�����Dn("U8ً�T�ٽ���h�j���l���DR!�H�{��:������ �~���
�P6�5�����شn	�0N	d��*�t����Dm�K8&N�k��k���*Q�g�G�3�<�_fj3C�b�� ���Fi-[i�WM��_<��b�k�ڃ�����Ş\�����V	���1�x��׸C�4�b�mqUu+X��3�	n�3pܶ�4;f���N�����Z�؞�z\&�s��1N�ע������j�ӽ~[4�5s=�Ӥ0�a��H;u	��m�c͢��t��>3�~�����fؒB��'�M��B���+��]-C�G���1{�|jcw�:����O��W�a̩�.}�]m]���,�!d��n$"�w�]�:2n�u�/l��XҾ��R�l��i��1	V�(�7��W	��T��]��Tg�٠�����y[�Kdw:�����[\oa�8.OA} ��t�9�;S����l�6!�_g���@��ęܜ�.��g #c�~��u���B
�k��o����"	!�mڿ��R�*2%[Th�|MzAqQ�xH˃V|})���X�1o�S���c�L��nI����_��Tgu�#�Uq>i���6�������C�f���g����(%%�7y⟬]�m	��Ӈ[�R
{�C&Usp����a���]�hsɦ����Y�Q&/�[W潽1�!�ı;�Ǣd󝒛JǄ�ђ{�Q�j~i��s�L���xd����U0�Ԅ��X���� ���I�qH��9�[)����J�oɯbtz�l��8'X�M��Z�����$5������>6�ZT���"�w�R������7J��):��MK�<���|Ӗ񮪨:�>YW�@-��&�����&�������W���8��d�M��7߿�O.�qr�����\�B�o��� wwa�ut���T��� Y��J9O�q'�������BB����j �v���#TQ9jln~{[$�;��MD��Ԅrۏy>�r4�%��W���g3�'7M���k�F���a�Ҩ�p/-6����Øl��J&�$/��(����_�O�Շ�צi" �\-&�{���f���R\�����Є�sba����Un���o��O;Y�/��U�>*K�otk]�XS���5��{�j+�~]J�T?^��j�C�|�Nt���@�n�1��/�}fyg��~�X��!�ƫ�U|������1|,K�	�VWǋW7)}�BM$�a;p''������1���Qt�����,<W��S�%�����$��]��o�X��>`��q����1��������M(��9]h><��;�k��E�Un�8�4��*(cD�d���w�[�U�V`�
���ei�k����5�+�z	�o�YL-�"R��q���M>*��am�	:u��ő
�b��И>?�W�Z����wM�_S�}d��F}D(p�/��פjo�=���|�tu�>r�L.��-������֭^M�) ��af"]���H�]�U X���z�O׸��hj���)RN�h�!?�m4޾���.�iW$Cw�'�1ُ{j+*���)n"�K>�b�� #���_���^Z:$89ſ�+M�Ro�H�+	M�V���:�;��ם��]^3�d�6t���v�7S��  �]'�Z��񇞦�#��t�7�rbD(R 5+1M��ύ�Z�M��z���Rv��Y�lW�":`Iqߔ޶�-���7��#�t���yG-��a��S�J1Q�E�>�ɩ�5����+�Hsag�ļB��t@O���w?�r�:�0��\w��;�I�X�rj��	B������� �`VO��:ѻB�!�i��. �9gR�,��`�s2<A!�帥��X�q���*��%ȯ��$�y�Z��m� �	喅@����L�U�bF�5�T�"r�t7F����g�y����^��mvW�1}U+D��S9���[gs��=cAP�����l���R�����U���p��D�4U�[w]�{�:���@c� I�KZՐ�ǌ���f]��󵅃Q��ë2t"�^w��$�Z�ى ��B�a~�ۺ�!Z�\~��&��f�yE��Y`������+lZI!��@/���ҵ�s8���;�0���_gB�10v!Us_cڢ�����7�d�R�t�(TZ׮�j�����O�Y��-.a��N�J
�e��Pc�Ӑ���Y�1�r��2�Ul�0�Il%�;#����m��~�=7R,�9{���to؂�P���Z���F�;����fa��+o��� �x�H�>5���c��;�]62��)����o`kި�zy�6�ͽC������1΄�P������`�w/!ӾO�(vɥC����ᨪ���(�V������欘���
���$�������I˭�}Do���Y5$**J�'��n����
��~WN��7������͉����>�txѬ�}�g�k/����}�
�'P�}QɏnR�V�)����y��(���փ����?;��ԍW^�;W1�&N�谏��Ou�]�E2��0�U���a�Sh�~�=o}z͹�/A�	�竣r>��g87t��9R�����$> ��ۗ󟺫E�뉳����,���g��㼡~�֜Y'3hĎ������9GnC�a����Q(�1�>�చ����/RN_A�㥙/=��pqoEv&�I�/B�U�uM�C�i��1����� ��E
UE�N��f0��}�%|rw�s*��h�4� ~mB�o/D�ۨ���n�H����(:��c�WH�@NI�����H"B�23�?���eF�-�f�ė�H|*�"<���_ʧsӐ1bl��C�O���f	��f�,��@��},�����3���]/3�ݮ���3��87 ]]>o⭓���.�{GȽj�@;���KP��U�܍�r���;Hk�3���t�,���?'#���lg�'՞���bޣ���8o��G,�;�G�gϣRBA���'.3��tiY�QVۅB�U�P�t[^�2-����}���;g�ez���-T̙�נP|e�"f.���r������ZQUr�����G+^x�4:t΄?�T>��7�����#z?������u�%m�E��Q�zo߶qh��ܘ,/!�bߔ0����}ZD\�mp�G�aD���BY7x<���-}���P���hv�LY�E��X���{=��Ӭ�!G	S��I�F��,��F1!diA�Y���u�����d��3��*�j�&��E�oF�eç��^K@_V��S��z��v}UF��Q6D�'����X�SU�"&2����ӱ �O���n�s�Ry�qk�������ݜ�VS����Gs�/��
�����^Ɏd�~#crlI��I�2˳�.�!��o��a^'$�|��pWj������nj��"�o�"��f��C�m�>������{����į��˫ PB�0P���Go� ,������H�bX��6ϖ�#��1	k��$��3�}��X;�� F�~�����{4)��C��iV���KA��8|/�@��=�^K��2����6-�GG�E�o`A�Xi��#�����AAd��.&��ks�'�y��&D���T��&�Sx*�Sح�S[��7�@�p���ׂ>S-45����6`%d�#.�t&�N�?��Tq:L�#e��*?d��p�S�h�B��\�ۥac3��Z�/\86����yFݢ��"!Ud;��=��M�3ٛ���2� �N�bVl�Io�h:�3fE6�c��������SZ����G��9lEc	̑�g��|�"�z��"y���
��e6d.(�������xO�p-j.b��7K��o,��e{K�ɲV�B��_�KM�.���u��
_����dѾJ~�y�w��׮��JJ���56f��dE�O�"�D����������4�5��?�0k��y�N<�Y���1�?�"���^�.	�.���` �ҳ�dQ�{s�Վ�H�e�p3�	Qu��^�i5ݩ�,$�M�����c=����v��(�?��&e3���Dc�c�K{4|'$�=������.<{N��2N�Nv|Ý��
~�����l#�``3H�y����O99��^'�Yǳ������G�\�K�̞��UZSC$�s�O����_��+$�%W8�;���I�pځH�����ڙ�|��شq������h��yOw�8.�`��6G�JVԘRBw�p��5<��L(�$�U���b�h��׎K��M��
e;<��z�Б���.XDJʮ�kI��xl��U �mlR���|~���V�~�gߣy��#�5�4U�Tk3�}"�~�*떃x�i,5cJ�+�%ͅܛ�b\
X�T2���8��C:��Z����� ��ڸb&���P]�p��evR�Wo9':b��%AT̿8m �4϶6��m5[j̢��>g_�sUtHO�#���jݫ��RG3�a
�C�]P��5��C��-t�����v�H�B��@����E���|"O7���m��oߨ*D8}ⶦebR�����n���C��͞:�z�cS{��s ���k	��>��g���Z��W�[��a�%6��V~�l����	PtI(	��9*B�������Z�i�܄���)C���w�f��}����@�uܻM��Whü˺�!�O���F'"�q�Y���+z���6�+�����N&����FB��S����|*.�VM��������˹�&��@�藑���>�_;ޝq#*ۜ�QA�M�';�0q�%h��{pE/>*)�q�.�ȟӡ.l_�먨��aK/C�359�t����}Vɿ��edEGZ��J����ޢ��apj{�����WX���a��y,|�do[�o����a9�	��@3�h�ʌԈ�������^t����k�97G��ZX�>].P����w
�8��o�UU!�����n%q����W��6K���׃�z=��jqZ��Wۑ�J��!��7nP��ȷ��C?H_Љ Ц7t�'p�,��A���>�4λ� ���rqz�������l�����3����I:����{Gӹ�z���0l73���{k�K�
>g���e�pQq������}���1|�dk��e"wc��j3��Σ����6=�O�M���s� ̕�\�h>^A���{�T���|����0;��$��˘�2[��=k��釯��w�����`�$%م�I�#/��mNݤ����,/U�ɯ9Yӳ���V�ؽ�F�P�^��� �s{}�.S0�����.]Nƭ��mv�z�������J�#�_^g��ӑQ�� S(��K񥐓2-^q���Z�$�H��9���M_�"#'pL��#L�u�v��������'b�6,��A�hK�:�G���^�m+ꟲp�)����g -ms���%k:��*��p���H)7��s��y�����'M��p����;O�z�<;���X��o� �4.rM�M*��wp&10���9�SF�,}�5��������c��8�9�J:�7c^��gN����>��r*5�����D��-�˟\Vv֌5�-�t�����u�X�Ks��鳙$���ڥԑ�I~�g-�Ĝ�H�}����(���P�ֱ�eã/>%��3��,m�w����k~n7����q�ۅ�ŸS����}'7�F~�q`�W�a��:�"vs,�p��͎H�-w�|���iV&I�#U�	no���W���Pj�������q ���x,F&1�}殳a�.T�0�#����ym��B���D���X���/�7�E/.L���&�Kl� =o��ښ�#cT��
����M�{b�<X^�1Q �yD�2�1�_�h�7��3_%Ic)�;�0�Ԗ�&%ir8.z��GDI,�����~�������D���f浠��R��rh˻ E7�����έz:|�5���54&�I"�1���@� � �����Y��i*8G��N�탫��p�Ό�=�̭`G eM��n+���MYI��R�^gYi?��6�+aO�$�|�C�c٬�b�{%��6�h���A~c*����e��?���c��μ���"�YO#�!Jhk��QxP:M���2I�7���q.s�3��y�[�AT�K�;fL��-�����S���qB�@��$!��A��k�f����������N|���Vt���P��u�:��p���:��~(�F�H�(���~�&%���ѤIb���|�!�/*́�/�Y���qU�} �.�؁F9Ȓ2Y*���|wa�Ǡ���oz���p�VR���)����$EN���Z34i���/�ew���׮~��yJ�REt��m�ɜ��{�pq"H�D�%/\�t"�r[ݺJH�c&���(`�}ښ�i{�����i���F~	+H
�H���:ux9a�}�S7^!���8�t����˘��C�b���z��PW�����Uf�8�>��Ǫ�-�o�}����&T��r�l5d�l�Iԗ��ث?�Ŏ*����'��ps�Fޏ��-z�����@����f}O6��D�|š�+���9�m
�D^�r���֗0�j��U0K��ۮ����M���S�ȃC�<[�?�U��������r$⎋o��Qq�3����ԒS��
LN����R�@N��E9�aWO_)���D�1�TUS��Ti�l��,#�&ދ�Ds�uZ�2!x�8K���T����#!A��M�	A�U bOfAQ��0�^I��1>����������[�Z��b�ג▫�e�}Q`�d�.k�yb����>R|vF2�N�WMį�U?&$ ��@�=�%G�f�8��`><0K���p�	�\�3�f�ǂ�ݔ�	�u>r|Y�|�ޝ�*N���Z �o��:�m�y��|-�wK�D��B@\9,�w�$�` ��	���)C��j��E�ş�e�l�$�>�.�<�<�$|�s/�E�WP�?}���&Je�B�v����b>�>��Z~�
��!5�	����c���(�G6;����$�F#��̭��J�犕���b��Z�������[�Wq�aE������wZ8T��oπ#�1���Ƅ��K��1Y������H�����<�∥�%.�&L� �
Z0b�S{�ƪo��w��w�}�b�
�r�$i�?�uH����
������O��(Y�L~�3���^�%&�]f�A:bt%I]2��a(o�m2>��t7��z��䔥�@�|V� "�m����f��:`�z�#��?���@�o�	���\��`�T�z���N��򉽫'�G��o����䲤'�QPNϔ��3L���o�Oxŋ|���*jx�R����z�q���Vs���w���8C��|��D=����ʅ�E�7#v���&�co-����O��98��ay
S'���U�Jw��M��_>e`��)蛪�أ]�'F\g����p�
��"�8�|�;�ǒ�<rP��q���#���;�6l�s��g���a�1J=���ǯ�!�m\H��=�d�^}7+D:Jp2ICHdr6u}X�!ȭ���E�	�8����u^�:UNb�-u�2g2��.@����G�\n����E|�a�#^'� +��̈z�����\ǂ3qf�;s$H��7���U�=�zS��Y��E�>C QS?n?)��H��k�B�ќ̻��="bhX
)��̩�m�?�>ea�`Y�xY��<�������3B�1����|�'�o^��Hf}�`��O2�V*�!�%�W��������*}~'ؤ�i�ˆ�zR*�r-�����=SH�4US��$(�[*���YԘz:y�*�.c����o�9�.���⭬�.~!4����}w+�LW��kb���|�@62�;A��W0s��>�q�7.�H^��9`�rΝ�y]���B��6�4T4��mCM� LP�~���L�
���L�˗���^�^G,���bX������#����\������\2�����(�=I�sx�P�>��x;�^��k�v�i��#�G�+���b���n�h�[�%���*���j�8�+��m��e��_�})�W���v:Ѫi/���fPQ�ݝ�<�9�����^9d�yƱ��ћ�e���I�ʶu�!mz:���z�
Jz	�����*�]�e_��S��s��Q�z�M��[�*[��b�",͓"��Ig�r�JEz�׎x��l�� ���Fc^�{X�۴��dӝ�����6ol�����8r�q��[�HK�7�gLzj�U�Yqh��Mp�������%�7;�֔]�ކ�b����_#?����8)���6|w�=^�r�p���ew~qc���m���c ����j�GR[�_��S��UH_N�;4֍�����H��TH�
��Gm�dB�X����
0*q�Pfs�� �����`ń7��7�	�%�{A�j.��kOL��q���F{js����mP��hΨ�	j���T_mIm~}�s�����en�����IX��<�*��ݧW�G#��L#��^q��>���<�^qj���.��J���q2��e�T9�c����ܧ�bϻS���{��ק����|��[��w`�_S9ȫ`t�h$�;�F�9N���6�x]U%��hu����
��^qf}���<��
>N�<�����
G� `��8�:;�S1���,)ڊ/]H�W��$�@�8m]06/���d=�_$��y卟�[�,�F�%��F; OE����j�����]�H�Ǖ�M#�U%�`s�\��.Fw{Mt�;d?G�A􌕬r*�*����gpw����f.�������c8}����������,�g�YQC?��.W��Dpo���ºɽ�����_���;�#Vt1���{�J���]�xM�5��tD,�Ƣd��N�%��2���J��e����5p$>u��4��5*|�]�?�?���-�������Cԏ�Q��-=�<��Xl�5���V� ��2X5*��~^�y�Q���sw_�7�y���ZWT�
�^@�Z��v��%��{8@�I���s"�������6��Q���~���z�(���>E�CԨ��li֑��h@Z��6�ԋ�L
���ѓ8@��F�R)C��ѧ��H7��yZd�O�!76ʜA����[_M�x�.�A ο��7>�#	�� �!#�Z�K���Q�)��r�>�&�n�qv�Y�ƄT4~7!�3l������}�diI�uBdۚ�"n9%����4� ��[���;o�0��2��Z]���h6�	��FM�B��n1��	���N�c��6ja؍����M�g����T�(�ô/ٞiG[�4m�*5[9�̷�ފ�&-�{ڿ�#��m_(�,�	)¶n+�8:�''bu��������wx8�p��D�(���y<}fI+e*�#�CUuk�� ��潹i�KV��/w �dY_�U�e�d�J�f�(��h��qǑ�w��+$M�,��aNN�'lg7�*��S��4�}r�
h�	2��W�`���r�D	�+=��H�^�T�t������� u�����j�]9Q>�2�O���t�l�����|E�v�)�n�]\�{V�]W{'9��Ǯg��b���w�ʯEs�� %�.�&���fv
ޟ���sX�����C�i<��2�R��L�q>��y�V�i9��h�	Y�v�]�Q��z��q�Ŝ��2$��ط2ॠӕO�^�3o�(��W��Ed�ڪV����v�A^#�t�Tx��4��W���T��	
��N[1;�N8��fo����2��Óg�: �i�J��租���V�6_Q����*C����zǫ�� �1g�k+��`n|UC^4_?G�F��2^;J����~*���QP�s�'����*N�?]o����l67��k�@�hv2z긳�k�i�1
�t��S����{���s���P])��K�T��
n��b<�iG����k5��t4�`�O$E#�>y�����x*�
��a�����ǭZ�-�G̜3id��"�-�N9 ��E�w��G�x|��o�u�!��~���We4���f`#��>�����P�P�VL!>�c�s,v�`�y�ǉ�b��6��p�G99�����r���sL�3�zSUvR�$�f$y�ʽ^��$Qeq5oz��aA����]ڪ淊�����nw%6|pH�K��k,����J��gÿ�2gp�!�����p�4��?=���P���u�;�U0AX�������(�"��Us�E�p|������r��\f��SF�S�7���(m��J����	Gzi�S$����Ƿk�b1��E�0"l��`࿾SR½H��f�k
&�e�V����3��Ee�E|p�1�G�k��:����荀���8�Z������9�wG�˲�p��O����S�SF��l���+��E��ǎi�Bj�;ڪgp;HMM;��k�����z���/�,�8N��:����͐����):J"^�N�̌����}ӣ[wIӂ���-al�a�ѵw��JS�Eۚ�TǤ-ґ#Lg�N�-(�����}��P�F��&��~#�Ŧ;���j�k�l�9	v/2����<�;��&�^��CE3T�*�a~�����zM�X�0�Q�����ٱd>hf�n�{���u����q�����V �k]����
e��tu����Z�wb�݌��`�`ɵ�˝�e���̤v:�"�n3�!dx怕�]���d{���E��zE��)fS7����@{v��x�W+f���T������*��<���;L��1v��	/�~d��3>�
K�u��%�no!�I�4}TT��6JI3�4:t����ݍtw*��Ѝ���tw7�Hww7��w���?�aւu�sξ{?�y��w���YY~�
d�a�������6�e�^��27�;�o<������T.��+�@
�f'DW����Y��raG�ܵ��z���Rs��Nh���}� �n��n]Gw�3s���n+avs�r�R;�N������Yv��c؏�� ��0Zf�Țd�p��t�OC�}��zř�I��/��qډě���Q��Q�(}n�z��"H7	��d���]G�h6Ù��j@�Oj����=�8S��7 ����y�ם4B9��PO�����هIq��u'�w���h���?��e {'9�M��@u��+�c��A��\<u�f��ҡU5��E�|��3��I��%�f( �����(�ٍ&���(K��<y,E�4ڗ_a�N�~0q�Ø�G;�F��Y}�/y�Я���xu�L�8�߂C���E�&��IQ��c}�}.���W"|�k�l�LE.=�]�X�OhtL����A��j� �䁯�B��{�=3Yo}-�N�oo~����_.S�1,�n�}��;��ym���f��E���M6����2>/.	C��s�
@C@o�tg��79���ݪ�j���h?�A�a>��_�uv�ϓǹ��!����r��󸀀rj9�C��F^��Ѯk��X���TH����?h�9�MX��s:&�F}P�����掺ѹ�1F柭WK���n�~����x�n�ڞ�Z�o�����T[�G��h��oG����v�GҧIgAc y�9m#��N�����S�0M[U�f�b����Q����������c�ǘ�S���M�J�����ù1˪��l(�ؘ� �}}bcn3<�NO��<��� ����!�� ;����¾�M
x�+E�~H�7���Fs��5��u:N�²E�m��1��_>!���-k_O]QVb��l.���C{�މk�_���6��zp-*�\Z��@��ؿ�)I_IzR;x��6
=uW����f < R�.Xu��ԓ��A?gU-T�W�Bؗ��̪��v�l�ݻx�M�f.&!�U!aBTE��s�[9���k?5��ϯ�<��Wg�^1����"�A;�=璮p�c�������C��߼%N$Ԁ��QZ�v\�`Q��n>�g<;��:�DsGn�=��QG,�%�|hA��s��~�ی���F�1���ӝ�����T!���Z��B�f�-�_�˳��&�n�Q��DSϭ��'�0S]����bGΜ���H���P�C����8]�X�r�6���՘JǞ�8�%%%)��!{��T�
S�;l��)'�}[��6�+k2���L�e��h<���BRd�ܴ����z����R+Ŕ`{G�2nbגsDP���[��߭�:)g#+{�bf��[E˯Nޓ���6�
h�L�k*E/�0��h����7AF�b�-+wU���h������M��ri�W�q~�zӭ�����L�?��39H�qm�+y��v�KT�����j��/�w~�\������L�K��ر����I�y�z�e�1mܮ��ᴨ'&F�-�J���W�����d�����5ѓ9Y�V��#� ��[	Ҙ��b�Ս���MĜ	=�:�V{3���չ����qۿljM�+��4��1��	���E��0���V��/o�q<U\������5F�� /�]����{ᔝ�d)�$��d獫1=BQ����\���Ӂ�+�=�v�!u�rG 9"*u�d���1�s�K�#{e8hb��)^������Q���h�D|bY ���o}���Z������Rm��`Lmp���c�~�ٺ�ëĨ� ���H�F}:�'.1S�M('Q�v������3�U�x dDDw����)?�f)!J�VVVc�����_V5��8F��(m���!�/Gƌj6a8����C�޷��6 �Z��[/}���u��������\���R00�.��2�yr;;a|&)�v��@k$-g(��g`RO̪���@# �g�DԪ~��Po,)@tzv�)@�Qzl�bo��fOJ�檡РVshO\�]uu5G�����|��ZW~d*ͤm�۶�S<ڏ��ʷX"��]�12*.�3�d5�;YtZy�l�J���eU�^W�9�Q�.�ئ��������B^Z�Т߃�3�7v�6F���}��M�8�y~Ꮞ�X��^�G��8������4�`<)��V=6)uu�+/!`���A$$��yČh�0J�?#o\� �F���bu���,�.�t��;J��wق�^^ܤ0�Wa�)߾^�;�Z��f��h=�J>3�;9�}we������w��.�8�v�͓���]����tRkAŌ����Y��r�Ww�jG�?�h#���ӕKke��3�Z
�����މ�!������l�xu;{��� �E�#�P��!&c��6|��ɟ�Ds&�I�c/�4ȍԯ����ƦK��Ϝ��F	��'�6!u�h�������Yn9��2~�LZQQ��ٹ�pC�˻���YM�|�P����hQ���x���V ���/F">DM1���+��^8��i��=� =Z��渽^0��Q9D�CL������� �[h��m��0�㱡Z�HA�[�u-*��2.O����>Rw �mC�t����j�JOnE�5�.ߝo������������_%i�����K�*�����o��_=�7�0��D7e���&9(9��1��t��d�]���tv{�-�,����TqW{�U�l�4:c�����{�SيkJ�.S6<�tI��bɐaT81WD������p�O�_�g`��l��?�F���z�U����H~�M��p� ��5���X����Oc~	q��,8t�����B�:����*�O���H����[�jL�&|�n��}��1�Eڏh���Z"���D���c����&���]*kg֮�h?���(P1U��bܔ���t�e4�����^������~�@��-�Xۏ���G�5�Gt���-{ڰ�^KQ��u��H��ߢ��M�,vq�qY���E����v�R�t�8���2G�NX=�~e1�V���#�N�\���Z�A̓y渴;c�Ƨ3o��+��{��HϗɥX�_��س��yN�����'G����o]
���31c���v7��.��T��J��D�Y���G��PE�$:{#gv��GXh}�9m�:�|�r3Y��}s����@\Y����g�� ���	����̌ٯ��]{<���]��I9O���u�	 H���;˵�c�w�S��\~9��[?GQ�Pvn	�����A���e6���L��jL�r����B���7�}%񹶐���m=X�ކ���?�N*�tP?��D�M��-���&�r��U	B�dƕ��j�K�a)G� �U��Ԍ{����SK���\G�� d�I�o<���2�
�>�!�`q���rnB4�bS�@z����mX[�N�Z��V��`��<~m6y���!Q�+�,���i��#e������t�$�g�:G�?��Yl�gv=��fc�u�=�ĩ7�e��E�]�4i�$���.�c�������yה��ͥ�m����zɛ9r�k����C!�vno�%c��u
�>�q7K�ע��a�U�d?�I�������V����|Ή��w��a�9ﵫP����8 ˤ!�)��鉙�4�&|п��*�=_�HV��F������]%�j���޾D�"��X���ؕ�&3�H;���I3ƅ��h2:	W��/��Ɔ��1�+Ԁ������K@��C�p�/_w����~㭇t���(��u� s�}V�t�&5gˮ)�,��b�i��2B~��zT8=l����K�m)�j���q���ob����֖H�v�$D��]�T]� +��|"���RA�.�0_[i�-�V�G�$Į\��Z�*^��.�*�+Sw,���
����N[>�Ru��*��PWY}�QN;)!S����Z���W�k͜�v�gάŽ�顈���[��*5���tsD�A�s|���=ۚ�Ā��ԉ�y�]/�a��E�����R���yբ�F�j��'��Vפ-�dJ�	��4�=s
�����aDke�}�C�}����,�\�7�=Y��%�C%Bt�}C�w�A�\�lmS�esyL6֑K�w����"���+��d\:z�*aʢ.��K���p�eR�-j<Ȳ�}�nǇȈ`S[���ґ�]6�ym+�`��jØ�m�
X�v�����&U���	����r���#Q�����X���w�����>;�4�EIUaM4屲���j�+~~��x��O��/����9TP��T���〨!�A'�R�,z?O& !���ȁ����5��w�є��S�@��K㑛������&=$��~�(i*�J@�N�ґ��^h�`�-�K�o/�����z�Y�D^M&TfJ����8��d�J�.v�\S$ V%�0����k��P
?�tL��b�n�O����m��\���(ɮ�>C�Y�_�k���&�������"��/��3�rR���.������p����Oc��#��Fw��j�u���bM�e��h�T����y�	O̩�1b~��|����?/�E�ԣ���oT�A�/��g���H	��|��P��%c^���H�ߊV{$�"~N�)bm�;{�"¤�o%�#�tI2:��v��v�7��zl�����Aq����[�>
���	��{M90�?	��դq��¦N��r�c�"�|���a��_WaG(���k4��r���������ø��Vc�>o�m&g��t�q��4�L�!�`�Ҙ1:C�^+�י�m}�7�ͣN�ƨC�vb���w��tF���ɧx3}>���HN_s��ۈ˾�P|�����/*1cw0����|hμ�O)�eI@dQ�|�Ǳ�(^:9
��������,�����M�~v���
�q	�룔����|�9=_;Q�|�A%�`5�����M��	�P��`��.cg���N�G�����L
��q#�����ϩ�'D������������Jpw pA�<]ڈ�6�v��]���e�;P�p6����veA?L���6�e<��.��]ߙ�R��L���g/����o)	������*�%�oht��\m�z���Z<���O��d���(��� ���v�_�2�=���pr�Sj���px3m䯂?`!����) Dz�ں�Fq�u�yY����Si%���JD�UZD�Y+y�K���=��VU�	�X(d�z]g}�zd%����|j��X�H\B����b�׊�������`w*�(��i\|��ҵ��0o&[p����Н��s��ʢ�F4*P�$'+��A�pZ�;��tU���j]��ӭ��N��O�0�F�R��#-/5i��,�񖐋G���cP�QW>=.		Z�"j�*Z���(P%!�g�U�}��93(ͨ���o��(V?�t�#��O�	�L�R����sT\}nm8u��3L�`+�o�"��=�� l�H��u��伵C���qe�.��e���e����Xp�	6�&��h�b9��1��(�A�8��g�����1�(>��,$;��B�����az�_�������^�~��� !
��L��b[ի	�"���oو.�I�k�F��";+�-�j���Y�������ㇷ��t�+rw$�(�Y�F���{[�;�_��[�|��`h�>��ӿ��[�/��
?B:芭��D��TήC��x������\����s�z�$B�聘FTЍ��������c���a��G,��4� ~�pU �?7�*��K�2�u��"a�eD���P.D�E�,0b�X-b��/'���C�� /qE����4�Ѭ��";�!���yECC(�ސ��t��&sj�d�f%UhÜt�{�x�h���棫�}׎I}��'GG��)����䇋��Z,��aEHG�����!�����^�?�éۅ�߼>Uw�����"��y�\���W�c�>΁�c=����?�=���"&2LU��t�^Z�[ !@';���l5�#��nU��\n�!3�= `"H�bY�[l��.m�92�à�m֎�Me�&��j���+���F�םj��;��5$�.gJ�K����Rdr��ry�kR��ș��b/���=~ {f��\��19�� |
�2��7�J���~�?��G���H;�l#��Ϲ��+�ݕ��b>9�12�*-�Q�4p@z����U=@|oyi�����������I�;��Vw�7JG
�����e���L�'뭥�_,/M��Z�vq��l��-��{J��^�0A$��Oo�}ɼ�Xu����x�n(CH�?��x����V�zu@ 6 � `G��m��龐���U���m����\��L�����-<*ӹ��n����y� !dxg-�%�5<�"g.;�5oGĳ�/G��8�/O��"�/K��Z����O��*5�T Qi��\��0�E��R����B���b�o2���v+����v\
㍙Tw94�KHx�;��@����9�|�G����ɧ?��b����bT34<L�v1�C�^�>՘v��S��~m�(�4� �X;^���E�� �ϖ�{��6� S��Y�O�NT��D
�U$���,�z{�����o-� �:l�?EZ����oN��8��Q��&#
�Ĭ��C"RR@F���h:~�?����;x��oF�s����n+���j��6�m�������Od2^�``p�~�M5Y�u{�0�泊��R��- �\��rQ�N�|�*N�ͪ�']i�D� �8N�W��H兯��wI.�f)�{�|aax^-RRe޾=���vj0R*����p�Ǖ��ߥ`�P
aK�!��m$�����V�:�#�<�M�m5X(j{~��`0�;�]蒊Η��Z1��)����+�7��s!�,U^;Hx�12B�2��=����4ρlQ���F��(����5��Fp�Rz�� �O}�y��:�pt��z�ن�)�1��N�)^�*��q��hB��W@Ś@��d*~�B���l�7 izvW�a�L��e�'��S���?�����9�>戚�����OI '�l���ZY��ly�ѻYT��Y�n5�Zj7�ŷ��Mg��W�������^҅ �YAc�maĦx�}*�PSf�5qûJk>���5=:zt�(GY��}J�Q^�e�O�����~����d ��dʓ��%�����v�0�ZsfX���o/= �T��v���z���|}�lll�?}� ���!���`!�c4��4��#�o4�L������K�) ��7��U=�����m=������{_+��G_�Q�wH�����:��͑S-�L�z��y�0(��r(C��u�oE߷*�����>���f��SA:�4�6Ԋy�H��ݎX-9��4R�0sd�w�h�-�ceu�H��[��A�x`� %[n��WH?&C��j������� /�&�VB��U��s����y�.�C ./�p��ܐ�Y�NNB_�5}����2�����B��iq��6�T�G,..6��AzY2�A�ͽ!�-8����s����s�؅m��j��~vM:Kw_���3�욠�M�N*RSS�t㣭�pҮ�y�r��g}�Ӷ���m?c��T�<l��eDG�1�=pʕL0fo>�+n	_Qn��vf����[A��U���&�W�:0��~R���eJ�f^
� 1�U4F�S:`���tlx'�*!���������M�݊�3G�Ltb�>w��U��L(�͚��t{u/o����,p�[��/Ln3Gl��:� �j�r�C��b7���&l����`��54Kt5���Ǭ�u]�2���2���@��ۘ1�鏪K��29T6~��m����yݰ��.��m!�ĽQ.�d6}I�*#��3mMt�����GwKi0\�
�ᛇ����iLQy�1���!�������[��f? y�����V����$<ٍ8rn.����C�f��R^{�L���Hh}�V��I�6py�ʗs������6�Lf}ej����΂�2���ʩ.�Ν�7G��7���!A%�X��%q����)� �*�w�a�& �朝����Q�cɕ�C�|�ua���0w0�z��5h_l}
�lu�8mD�M��pTZE#��@��@�,H�Ioi����QYA�vkE9��Y;H�-�"���~�)׊\�����g8�e���)4�śL��ԓ �_�a˜L���JA�|<$�B4ׇ�N������v��.@�Q�BZs��.����Q��%U�o���|����'�Wvx� ���f)0����˭��`�T�����f�#yX�ob��!u�T��y{��F���ށn��祿�9}my �.�є,�`��)+�V�8mR�ٗP���
�l��.�-��p5��_N`ye����_X]��I�������Ln>>jAA�g�O���?av�v��.�^" S�z�'�}pdg�m���P3R�`����7r��.��5��J>^U˻~<K���5}��`B�9�]5L�9B5/��`.��"~B�wߣ���Ўm�5m%f|(�n)E>v�5T$a�m���vZ9��k�CH� NɱAAo��Xl���N�Q2��f�����(���G9��|��i�OB�n͋���]�_�ô��AL��'���%��ۇ��6��&{_m58��1����P9�P�U&�ʭ<�.9"yy��U��d�2MH���UC����i�3~���] J�D]�ǿ}�|��(���d���i�?������/7���v�2�y�|U�4��mօLie���hŒ��.o�W�3��<�=�W�VN.�)�*��׍s�u��H؛�|�uM2qw{䭙[�V��]�]����&�6�����,!��5��{ds�D�	0�Q���'��8`)$���%�gJ�E+g�1:�����Z��ee�yضcɧ�GCU�1���\^�$��2L��E�:o��f��.�#��Oc�.���W�&�%�y�_��
�x��@�v.�ty'�,㘔֞G��ԏ�N�0sWvx[g�M=�	�㾖fa���t����L5Ob�rǡ����
pU3�M�f��N_�̲C8<D5�q�<�A��x�M'C��U5������T�U4ǁoNU��>�|-�6n�g�ie�A���&1��)`\��űR;�~�+'g#%���c/=�L���D s��P����*-��g�/��槚/�\��P���}U\��.߄��MJ��8�V�m��J���y�� ��^� ��@�~Q�(g�:�@�Iۻqo����|���FI3�C���u�>XXfi��<���Ηh	8"�F�̂��vln�9\���� I=�x�������9�~�,S�o'k?N��FM�-��N�)�$�N��������L�MmQ\0�4�OQ�=^`�ǉ�~Nk \}P��F��C𛭙@CR�jJ����>/�~�YQ��z}Xj�)�9
�q�Ѵ,���Q.7���*o���{�J����9<Z��� ��$9��/�����HR���Q��0�Ç`�m�A;c�:��H�H�^/�����lP������@��������|W����]pVA�'J�R8a� mE�ǝ�}Zu��O���MV2+���0;=��t�O�H��Fֆ��Dh��8�<�zWhX���g?|�@!���T��,� �9V�#�04��E��y< ���Q�tf�p�m�ׅK���v6�혭\�쭓�P�tE���v�]�5���9`9X��$�������L� h..����3,�]̺)�ĦH�w��3�@��7W�l��9@+�9�����<����u�U\_>yjl�.��i��^�J�.����Ě��+�r��
��uI��&� �뱺"G��X9�63�
�-�zź8Q��~6CdMB��M��PÂ�������s��TU�>��=?l�qh/������b7�O����W8Q+��1{h�A�� cr_�*\���l��	Y��U4$���k|���r�}�O��#8<��U�['uo�<��)r<�k����,=p�̴@q�r��H}�[�0L��N#�q�pu���*x�8��8�s5�+ܸ����Z�����_�[��}���Y�&-ǅͷ��7�����Ds�N���q�[!|t��C�H���S����Xy�T~ Q A�dM�ڕ�*4e2�F������(X!��%�oRk�9���o�fLw�weh(�mz��z0��.`F���$�习0�4+�	@�f��-(���ڞn��YE�;Q��5O����i���4t�L���ȁ?t���Ó�w!�]:ՊgX�0���CG�$��E��9� Z�uLX�g��PV�HW)��dBc����s3t o�H�?�
�3/���:�bz%j��F�S�6x����o�y2Z�����e��~�è"�F|�+��|�䚥Xx �%�#��h�e�����9t�f�jU;��׫�޻���}d~�#
��bOX��`�"
��²�ZY-s0CM@��E�ù�B/Fb���o���E���?
h �:�f��M<Pe(��O	ĉL.�o�7��F�G_5��>]6\���]_�|(R���w��=�J�)X�[���-e_y�N�p��0�w����ZPﹴeӉ�'���/)^�&�;s���_/�յ ,)�H��Z�527��~�����B@����-����(P\�@���?X(���~��DZcG�i^�(����n.bռ��*\s�	Ek�����w�D���euI��uw�l}�pB��a����LIJ:@	~!��j�(��.�9������pBP���<Pٽ�m4�	Ѝ,·T��z.����5��ݓ�{��:O���՛���G~�����*+}���o��D�|��5#��U$g�T���ꮇ9>Kz��K��[��X�����֎�Z*�(*z�7Y�sqq����eF3��n7k�]ө��������+eOwDi�m��ݞ�Rt��]�x��*7lB�P����o7\�B*��"�d�e��r�m�@xO?��9�Ғ��3��-2X2�mW�ƻ���}�_GYnx�mُ?�#��Dn��!��+��`����P��Æ<��a�T=EO�$�e�`��e�@�q-�7���_��{#�X;_v��o˾r���.��j���U_�u�����|�6������n~"���:���)c(JW�~`���|?��Uā�3� �&#��Pؙ�jѤǦ�B���ۗ�3D��ٞx��卭��XNIY�SU-%UeE-~\��+i4�����o��k�+D@���ye�w0��I�X�>"��#8S�8S)&�"��;Z���R��֒#o'�m%2草f�[����߱�V7%�� 9"��������Gǈ2C���$�x�8L;|�s�Yf>�Cݜ9�Ⱥ����e4��7E�y���.�b���Z���^�e07<�e�M�*!Fr����:#i��C�}[�w~��7J��jc�E���M��7��&%H%-1�v	�B ��CG�^��QD��#X���k�f(���e��F.Z�{eW������)A-xE��d��_���Y}���	Js/ 累>ھ|Ԗ��Fj�62���HO7�(WBO����c����]6�T1�?f��$|OB��}�yh������7= ��l�"��X�F8����Z����^��j��ad�"����y[�w#�=�<��ßZ�P~o� _�Cio���j�
��b5.�R�m�`\���X�/�R($����6�_�|�t�q�-�0T���1T�1�*�J�Et' ��&�B�XwZ��`��Ci��v-x�H�@�Tu���
�r��#�F�\�wPs�s�C���@�5�fDL^���� ���|%,˩��RJ\\hb�v$/p���Άi����YP1���$F*W����_���f�+�ԭ��{�� �G��q-��Te���u�� �fT/����Ob�˒+Z��X[[sI~�@��5������ "Ъ2?��Yy����t%NWұGd&F<��A�3�����[A��^rК3�^����K����\�����	�~������o�_�[��uY>/��3V���H��[�Bb?]�2p�3��vX�ؠ�E|��|l`eh0i�r:�Ϫ)�l�M�E��*�Jc��7�Jsz��Ol���H��e��&3{vf�U�=拇 ��W�Qd}׽��XL�%�ܦ���,K��A	PhKB��1��"*6�\\O8=���_���PRY��0�֖[ �|+�a�q��� �.XԴ����;ڎb~1�����(�/A��m#|6_'!Y��ʫg�.���(�	P���T3�] ����4����!,�0݉>Wq�8&q���p� ���Q�νk���(]
کz���׮Q!�q�����4�l�5��­�$H^�i�HM���%V��о�dU��k���ߥ0A@f�c�
��Lr��Yh�iKV���l>�7%G�
d�t0�����U���`i ����;R�K[:4����ٚǴ_�����彮�(��Z�K���_�a뉹������w�P�vaqs4 �qjm��P�>?�r�JB�K�UtB[I�NE"��Y}��Bﲙ�7�ëQ�,����0>̡C�P]�����G&KVm����:��>55��d;r�%���0�e�]]�
5|� �?ST�YN�<�ZpbJa����P��� w^1T	�i��h+k9RD���R:9eu_K���L��x����p��Ώ�����2?��d�\�4����
Rq�er��������N�x��>Kǲ�[�
8+��*�	A{%���".�h�55pW��w7�vO��ྲ}X�/u���b��M�Z2�w�fΠ�k�xȹrٍ���"Ȯ�ӣ�U�9T�7.����_|�I�=��i�Ӥ�Bz�3Jϰ�������է,S-�R�SP�S(�k�z��9`�I�p���{4)��6�����K�W�l&�E�tF�Fagc9r^�mU��Ծ2�v�$i�L�l��3��1#���Mh\R�-��Ͳ0�'k!�g���
k�W�I�J���� _ B���+C������(������(�t��I,�x�� �S[:z�)�v�߽����=��-����v>ͯ:s��s��I��{�W�c*�GW4Wj��)>�����q���w~8{�^�74w�����Ĝ����Sa3��ȳ��+d���7�7:�v�����M�A/���̰I�@|u�o�!wղ���R'[4wq�����w���6�x"�� %;��%��o�'}Sj;k�~�TG��n��P@p���_<��-��t��{`��'�+�Y(Ӧ�����Rs������W/i�婃���[>>��_P��(eO�a_9I�䍙�n���6&�6m���^��m���~�3�g�-CNZ*>�֔��iUU������"��>��w6~1�	�>�����C��b�������eܘ�yV��+V�����B�ݶfW鍪Z�����}p�_�����eg-G��mC�vۖ��Q���ߖ�r����\�1�$"�a��]3�Kf��UÎwd�y]����w?*�_��G@���^~��Ÿv^Q�)�4E�����B�<=�4�r��`�Ea&��?x�%�Nd�f����o6���ݹ�ԭ�V�d�~�
{	[��@����>�O�ԹF��X(?��򡄁�+����.���c�j������|E�S'��.���h�C�ۮ�\���p���f���Ј��5K	y3��W�Z����8!>6�z��lqͦA41\Na���D�̟�|��[��*L}.�(���DR&�ޕ�����Ul~��1�%:a��^�
�w0�n���BI�8���4��r�i-�2&�D���W<ws�OWXY�l��v{#	��&'�G]\�T�k�1�����f�39�{-��Y�)[e��A��yb^^- P�[f&���$�L=Ԏ�^�g/ ��В��Ʋ�'L�\�sf�Uw�������jK��=8�+ѩN�_�*$�&s��o��	5�7Rc��- �u?Z�d�me;l����?�w�O�(VA ��:��j�0̄����#���曽)�	����~'�������q��z�GT_��1�Լ\�O��?���˖����/T�"k(am0���k�c+:I��D��<^BX�D�n: �������(��E 0F�jxb��q��V  �= P�1�z|u�S���r��1~��>Z���+�o{�^����� ���7SU�KLL���$��ܻ���a�D���e���䤻r����z���|�J:����������p��#!33��ˮl��V65�� r���Zw�+��Y.���ew
��щԙAj���G)Q�����\��{Xނ���T5H�)���ݭ��gp`Q۬���?��k�f��+^��7ě�Wk�q����@]���XJU�0˫#��33�$�Y�f��&(�yx`Smql���6ף��#.���	����M�#��7=�8�}��T�\Vg�r�G9C�������a��ߡ�l�tK��?�5 ���ŷm�?3I�V�9�ޖ7u�5�=B�Q�j5�:��i���<����	�i������|#�!����=�5\h�r�5��"���sIJBl�S�I�e��?�G���Ni͛n����r�]۾�23�]��2��XR>�TQ=�����Ԉ+3C�j0^
����Z��%�Ȭۗv��ߗ��5cX�S2#�" �wp�[̶+�;I*<�c��Q6��3ܗo�;�����+�E�W�r�����}��k~����߭1ɨ���hP����[r*%������4��
3�+.�˲r��HF$$i^������a�&�b�N�����P���H��u��6�*�:cp@�l���_L.���@���WN�=B�W2֩����̚�.���o�X���\]
R����7����*:?��5���k�|8���xj���92_A+���n�9�!L�c7��K�K	��.׿<]��E��8R����!l�Or�-���x�ϱA���h�Jl���km�E�,G ��]�naS�C�6�ߒ��!��(Vܮ#}�k,��M�0��gI{����4�Ɩ�A�Tnt�wE�� �f��o?w�|o���`0�n�_L��o�Rcb�� �K�6kuUT����0�3$�C�0�b�DB6�:F~/������pH�o���� �O��ļ�G���þ�dx�mT�^��s�����ġ<�������J�$�`�����u��-�Pc��W0M��~i/�ݴ�7���ͥ����?��ܱ�HǼ^�H[���9k��ɻ�[�H��$'���²��"�(6�D����������sO���tȑä �Y�.��Q�$.o��%-l�*(@n�[i�_m��%���-��o}ٽ~Bd�n��� �Y\{�8�cY5ʱq�%B��t���9��kWHʳG��_\�ʀ����.����s��k�	�W��������J����r�G~��O�>"�
��QN�Q� ���T�8�"q�L��e86E2#���Bp�yJ;���M���$u�4�9s<��cT�݈M��/8��G��	�c��a�f��6������Rw��ڴȣ4l߀���H/z��e2�#�+ާ"e��(7G�1%g�i���ma ��,iB�(Ep|��J� ��L]�����᫧�1���C��3��pj]��f={�o��� �F���M{��X*����L\7TWA3!��<�X��D���3|�>b���/���ɗ��-��J�NN"��:�CI����A����_e3�E���#�i0�|(����F�:'4�b�ӿ	�Tf�y����f�����P̎/�O[$�O�����^#�oaXe"�Ju�3��i���vS���:��˷M��lY~�����>Hvf�^R���ffL.ww^	�&P�3/ �06`�N�3��c�>W�"��9��,�_��-
����-i��4��%���I��ܙ��wt靝�U��:|^�鋾OI�x2t��9V$��Xl����.���44p�%�v�ۑ���Χ��0�kEO��M�^3�I�����[�s%��(o�D��*`6�iy�j�I���$J�cs4�}Vw
��.��Fw��f�9ŉc���Ilj��Oy��4�hV��$�$!)���ٝomh�i�@a���2=,$=�O�n<t�i!�F��L� ���#��6����?qI|���B�{��|����[tۗ-b��@8�1[0������i��s�����#��N��Y���۔�����Ӕ��5���'7�λ��|o*�4"E�*�����UbI|eS��M������0^��y$N�D7hq1>���*���S���o�R.��q�+��	=i�FIB���������JF�㳷@��"���iT��UH����g��#�Y+GL�+�	�.��ֈp|�D`�f3�\[z��G:FA�F�'�����׼�8�4?	���/�V�$aK��L��V���ׁ�%��s��^{ס�Us�9�v���L�PAG�����X��@ �n$Y� ��^��}P48���xL��Ʋ��+�q� �$\�?r���Ft��ì�W-��s��d�RӜ��EW�%4����P�r��5F���v A����R6�`>\,�p�q�J��L7���3T��B��%�d���uTU�7zH�I���$�i����ЇiA����NA����t�}���ܵ�z�{�����癙gf>3O�����6�!��-s4b~�g��f��՚L�����\u�-m�ï���D>@<v�?V��]u�Q�7���Ypޘj�Z9sW(GЖ}�Z$�o���|�yO���E���7QD&��v'm�x��sb��M"!�xʎU���N�{#んoE��b1�Kw�t������d a����r�;Z�A�F�J���"E�<| ���uܣ>��v29�Q������k����4��H�����3C��܁���od�
F�o�	D��¿��N�RP鱒OH>Y 	}ˡ[oB�|;NKB��
L�'ri��e�����T���}�U8�T̲��m|@�%:����D���[׉"��5Y�lŽ��j�y��U-#s
|����Kc3֣�>: ��n�{חh�>p*/�y5����8(�AkX��Գ+ࣞ� -ە���uU�Ϫs�ke�:g��I��%!>���2�ޑ"����40O�y�������[��ڱ��7��߈ ��m̹V������9�ׯ:�BU;vcJ�C��ի�ǈԔ�KZ���|�������~r��R[��%W栅�%.�2��12'�M?V��5�N�������q&PPR�[�V�p���4H��? у3aq6h�Ir�G}qk�}���%��˯����]~֬ 	��c7<�ّlIC7B�;n�X��Ѷ��>J��3���V�ʹ ���km��q�O6�?SEL^\�{?����wV�.�����!}7Dk���^/�Ѽ>H)k�!��!XE�q�a�9�f�/3�\|�unF������	��N�U
�(j�}dF�:��a���#ӏ�#O�L�����8��ē�������N���~f�p��X��6����)���@	z�
�2W����c�3{u����j���\���K����1碾��n�Ќo���߿�sg��s*�i��ڂ�K��4�-�X9ԛܚ��773�����u��	�ٹ�i�^���uW��s�O�b����+bwy�۾I���Mlp�m��b��1���?��쀶b<�M�w��G6B[�=��n�^*:{��~���jT�X�{�3('*�,�>�|���5l���mk!Q
�oq'�6�~�8���):���e�@��N�����g��&}�g�o=�{9��f�K�&��a~��{1��{EP��:��[ɠ_Q��|��/��b��ƭ�z��O�L�K�E�$�.�߹O��:�������6zk�\s �K5�[��	���⭤��j-[I�q�����C��GQ���
K<�.�9"��n�^��N�!!�7��"�w�6r�������^Bg�.o)�@#R1�r�e��mE8r��L'����p�\��MT�)b5��Q�G��s�HҰ�y������˝�җ�4���{"d�Ӻ>H�
W���m�䂃4ʟW��tGS���{��;ƽϷ�؟��#���ǯ=7�4]��z�����3?P(=����ʢ��H#�+����˥i��MU����X�x��Z�8E�޸��U],]�
{ܹt��i_�F+.���|�Õ+/&������w�'^*۝��Ǧ�f�LW�����N���3:��)fj&��C�����&��Ei�;��9J6]�/�R3v����c�}���v֛{Z�IsKK�vA��*�ݢD�_�<�	
M@���Id)�ޠ��̿��we/{��g���\��z�Y�~J��-T{0�e�y.��\�DV���/�ߓj��J�0�ř�[I�9��xd�}آ\�͞�-Zw��q�	���o9�m=�X!�A/.���m?
5��<̿oo��4�+�E"�����T6�:��6نwv�&���P�4���}�`(-[s x�N�X��r�}*23P��ơm��eV��V��W���%YUl
�aa�))�V,(�6n���&��W�S�k{�3�F���<5��0È�Dr�
͏���<���\��ܶo������I�o���xhliX��/����UTp�VR�\�-�����9���;lv3ŧ�R�\ˀ��I��T���F܄%��Ug]�GB��M��_���3Z��X1`�����<�)�K
��T�7�h�Pb~N~J���c[�E���f'��ı=��g�Pt�<��t���4����"���j��[eښ$yҳ�&M��CC�1��G�H�g�<n��� &���:Ս!R	�њ~�E/�#>11�V^�%%%5��1�c�>r�@ �"/|N�-�Y�(R�0&�����|v%�-Kdh}�y}Պ��@;�ȡ�-BK�j�Ҷb��kqj�������>mk��}/q��NvsQ˭���L��༦�K��{wy�S��Y��p(��q&���fR9iQ������a�2�jt�;���<�"I	6���н9�=����B+��6��������+)���E���SPS
D���L��!++�����ۂ-O�.����6zB�WX�/.y+j(�s��S��Ut�]FH�F^�U���_o.��{yW�)���TMC�	g����N��[C�����nط��Ǉƙr#�J�{��*8=�k��ӛ��. J��T���t?�i��i1���<K�u�<�:���FA/��5��5�$~[�1�[o�W�g�������`��pr��O	x��J�c�I����n���a긻�QR0D\�n/"J��bM�un������\E\h��E����:�X�k¸��|��;�ᕕ��b�b�|�Y�-��x�w�4�o�ST���o+�[���f���\�c4�A�G>�9�nР��$��"�)�$|�����Q[3��EZX�����=4
%w����q���+��.T�[�ַ�W"���5����?�R��V����N���5&R��H=xz��vQO{���VTT4.O��leY��`��;�،��/�>�i�&�Je�d�t<������)��gڹa���t�k��ɵ�o��빘v��X0ŊI����y����b�ϒ����<�@��:{?e�*���z� �6����Y��r�f*	WNZM-ݍ��ٚz� ��q�]��)˘Ch]CdR�+,E��7�>�o��G/G�,�
9��z%a�`r'�a�3��$���}���0����L�;���y�ڟ?W3ccy�>�m��t��tӯ!�R�� x��%h}EKZ��k���.��!���3�0��u����Ÿ����2�B��1�u��y�NaT���+$/��=���	Fۇɀ�ne���gT����]���x���+��z���������'iL锤�įV>.��ی7.�Nz�*r
:�������9���QV*ě�Z�&O?&b��;�$�udmL7~"���iq6zl)υa�7p�r��J6h��zumK���^�,y�S*��s�@�	�| o��럩�
ڨ�/ƛ�@�����4���zz>�)�=�q\'1�t/�V��c0(m9=ï���O��8��m��(��bk+��[�;o��L��1�?����S������Z[�#B`gx�B��R�̭j�H,�}��Z�^ ��_}y���f���
]
���&���sfP�9���ӿ�k�5���Bf*C����t�w:�*I�	"-vo�F\0X�H�D�_|���	T~2%�����M ���\�'��;�����^����r�H��C"dŰ��DìY����@:�),P�����>������i����T�+�V��(,����z�jz/`Vp�y=�_=��$) ����n�3A%���E��śX��o��b'-�y�$*�*\"�R=�\)^���t�v5�4�)2�M+�jx���O�IJ�\.����Dd�I�M��ڇ�i���(}{��):~�1��������zd���8{ƟuG��+�H��p���ݪ���L3�e5�K�����Ap�mI�}����	�,�7��$X�A�x��38�i��p��vE��nk�h,�a[�>*I���$��*<�c.kY�Y%������_���<��8�)J���Uw�XQ�@m�f�6Ƃ�}'���ss���8���ߞ=ր�\�S�/#Kj��g|�O}�,SG������	R�^�3]Ȍ�|��V�c�U�DoVԦ=���5�����_~���$z�x����D9 �9��6]�|A���D'F9���g�)�a��]�������$�ߤk�� �8��� ����E2
��NuC$�.
�qB���ց��!�"����7<�%Yk{���fy.�p�53��7�y�4��<*f�Ŕ�/$\������h"��Zy����rm]��y��W��:	>~���y#��}���1����o�aJ�a�1A̶����`����-5#qHQ�ax\M�oj/,\9aw�����5�х\]��<���Ҷ�D{��I��o[��e1��6y��.���Q���bQ���;���(���C�� F���fS���)�Mb�P& �D�hc����g�}�?]�E�}5([K���҇�*?h�m*�{Z�g4[@���p�'w���Ν'5x~A���f%{�j����<�*&n��Y��f��\~��d��Y�o÷��Ow�魆�6�aa�8�^�ӌ�9w��~Bg=�P�����,43U�^��9�h�*���o-@\�3�7��w�}}�3� �
�g��]�R/��6m_���&���ю��s16~�MD��^��W���i�Vo%n�CY-��ğ�(��'����/�ܩ����6���XzkO��㡣�yΚOQ���fc岵�@���ub�V1yl:��Q�y�WEEE&��t>���볊
ؽx �x���zc+K���32���5���vb��/_����W�6����1��D�O�}
� �x'AO㵒e��\]�{o<�����#`.�4� �c��W��V����Bm{\��B[��u'��?�#>8�D�a[]�u���rI{�����8����8Sm�L3��ju�R^ÀO���Op�il��Y���xNr'�1��Ehw���]��\���Y� rJ��O������%9#�4y�Wi�L�ņ����ǵ��9�x�^"��1-j�uui�Ϸ̇ḛ��l��만�,�RQ�w�j&MMą\&�D�3��}{ү��ߗu:���4<��Ѵ���w*�%���ڟޗ���`,q,B����T����{yE��l����B&柧2��M6ș(K�OJ"�6:�L��������a�f�B��<44X6�uR����'{jĦ8������W�K���R
�@�d�P `TT*���7Lhvl:�VO����?�,�ʔ�LQ��sp=l�%����Qc�*�^�j�ws�E��!*aS�]�I9T!�o�8�;���d�D�_�`"��ž�Kk�~�I�QVK�~�f|�2�@��W�+_N�2�"e�n�j�!:�v�-�oY��"�WB���s���/���N��W��J<����n
���u���R�N9�MMQIO�^���=�XIg Q(*�*m4��='\<n���JT���Ο�
���@����aUڐ��<���oت@���.KY4&G���ҳ����H���6���d��;,)o���K�y�����:u��G�CBi��������Bu�lUK^6wL�L�Pk���u.��EL/��j5��.��}q]������27�u��Kt�S��E�}\�|��@��i41Ͳ���������I�����_��ad4rx�����_G������/����@⹑�/�\�I��p�ΕA���R���^���+l������0�~�騄-c&�]�|�[�c�9aͻ�k)��RLo'��A�>��$�Mu:c���G���RNr���b`A���4Q�V�������N{YY�%�S���g�C�V�92)�yE����XEz�x�S��::�>��yez$[���ǌ`Y�"��纨$&;
qh�F(z����נ|ug ϥo���T�'��ߍ�2��|3o��n���gE�؆��jGgf|#�^��A�DQJ���p��2~��ɠ��� ��]�"�ēQQ�aj]c@B�k� p���a�r
�܄�
��xC~��3�p�a��Qw>�R-�������А�ebS����=Ü��9�r����ا�z������������2bknB�d>d���+���������W�nz�xy�A<?:FqHaD���-���a7 ۠2�D��I+un.bpv
��I��:&���?�VOu��S��B��l���I�(.{WCs�
��z-���ڪ��;��%C0���EuN��J� +�Ʊt^��}(�I++{.�~�lg4���U���o x������:�W��i���d���'���bt��D�6Kd���ĖA`[ɐ�ڷ�PwZ�춦�a���_k0�O��-���!N|���gE�E���������Q�L����4���J��11�Z����K���I�X�a;U�;g�h����]�Z�Ͽ�*�'����}[~x���H'+�=���>��\ԑ�����<,���p�Uk2�I(�'�ИWK�\Xpj�����AI��~~!�9{hnn.��*(dP�Q����Ju7�ٗ�i�2�җ&H��J����C�wb��,�_a�(�sI�ϫ�F�y�H3.��sR���<OE��A;i��%�����u�3��|�Y�J%jM�!�c����[��D>J�&�N#�D�x|��ꓤ�S�F;��[�J�`���S���jy#�@����Rx�؈o�[�5�s��k�����?<��.mݿ�y�Z�}w���k��H����r�_$�Tk���[^�4{w��y[��k���K�-8͡t+�E�c��p�o`.�ӻ���0~��Ա�w�[ �.�B��\3f�@!M
o�Cd���22��'I1D�_V�e�N�'n���hb�����p$�f���^�Y,FHa2Ҏ;�W�J�iv&l/.����ͱY}���e54��m,��6l���c��IL�3?�'�/d�vN�B�y��Bؓ�*�By�ք �]�$ذ�&l�S���"�Đ{#�U��k����:�Җ]�M܉�iFb<�o䢁+!�%m�>N8xx�\��OX}:3"öP������m�pn;�A���K ���	m���b����E�{�$���k��m$tPy�7̊=U@Ok?��Z��և#�C;�\�n=�]��^��˗ۯ~  ����S�$�q�K�T!b�������ʢ#V�.'��{Q����������	����9����+�z�XDط��q,�?��tt�������pY�HD����w�UY���*��m�#�b�� ���Ӗ꽚�����au�㻬�2�p�N��4 ��kl:JtTT��>MLMe �|pp䛓C��y�6�[�.��k��/������5I{O��BF#�M���{�&\b�%v�4�U�����SsrL�4�&=������6�-�S/!�_r�b�_m���ޑ�-q�������d��|ر�]����-��l��nU��;ؽ�{�^:��?�e%�[Y���̳2],G%�\ޮ����Jd���	EII	v�S����� �frZ�gͺc��Ni}�׏E��G`�߆�Z���i��o2��z�o
��j�������u�*���F`�G�E{|g�u��{�Y�)��H�x�|�c�n��������A0���0h9f`?LE����¥�pS6F�"8O�Jlqi��qx)��^e����l���,�c�r�������n�8�b!��¶��1��/�-�#E�ʗ�ޖ���#��dHj��0�wn�L4--�� i����9�,{���6��1$h��XG䄂�������e��� x���Md�K_��p�]�����?]��W6K	���������^{:\sJ���F�����nSvv嶺��?;]3���
[T�c7%�5<�����'.H��U��B���^��$�_���wX׋����x��|f����0&� ����Η�n�5�UU����'[�_{L��/H�4ɲ�o���OK�`|���5嚯VV;�mokNp�/O><�C��#3�%���:���5�j�D����&��2n�m�?^%���X_��:}�a��'Y|�^�*���{�A$�����K_^D�o:��B"��Uӳ�@m.Q�-Ǜ��B��V(�2clOw�m�� gz���e�&<�o��V²��>�r�SJ�r�	�|j����hF�"JA�&�����죰��"��B �a�N�f���l����x�ߧ�_g>��Q�� tJJSS'��pq$�oq)SWXK禴3�| �^1�h�{y���3��~�8����~m�
���ݼ��,z>s��lP���K&��5�
��������N"�-�b�'�]/8\�����3���t-�tj�tk�ƽ���J{I�>�`�*d4�2���賍����u�<�X��뷟��>���-�e7o"����#��@׆SgUV�2*CCUZ�28������+W��M� �P��E���ع���f�OTD1 _�km6�G�W{(�\8l�ŉ�Q
`3mA�ԛ]�-�W��7^�������������{La�xH�o���Ib8xW��MZ���`H�T��|�|�HS	 �(R�k>��4��s����x��, Ь��{�Pj�$j�����WQϾ󑔄�E��w`q��M�q��o˧���˜�N�����<E<�sœ`&��@L�%��i���;Q�q\��$[!5�_-���}�E��'�]
rL���� ��0����{���;5��ۋ�T��9b�b3甏��ݘ=� �w�G߇q�-�e��n�T"���b[Җ�Y��~j\���+�,�p��@|��w���K��w��[�T��Z��~����k���^�^���ə�T�x���P�ݫ<�O;EJ�v��hf��R�r�w{{_�u8]���=�5j�l���+�q0v�p�?�q��5ʫ��.�b�%�/o6�t�.��K��Ȩ���@�����Ho��{���+c��|��������E{�A5Ωg�qy:�"M�����w��"�M�q�z̳}]΂7ͼ=�Z7~����ك��X�,���n���yx\�쾫��o�N�K�]�$.��bAu��56g�D��F�N����2�w#���t�v���v1�}'�0�K�UUΟglsVɄ�=�觊���"����u�7�/a�6d�~＿i�V;�z�y�?�Z]X��x������R�ى���ܔ���'����<�mX�Ik�2�ry�w��Ǖ%�����v:O"�6���[���lכE��0 �	�u�hq�Z�� "{Ɨ<x� ��9C�癒�;Vz�v�h֤Y5.�ʂ����*��K��D�U� POǛ��M����8�o/�ec����KH�����o0�0�r�����'{�1s���t�@��QPP6\������~to?����>�k�*�����@;E:1��ro8nXl�d���o�`h�N9��f,���{@�=V0I-e:Ҧ�G�����)�Gׁ�pT��,�m�E��7��GXc��Ҏi<_8�΋|;�7k�_��/!��D�EW��k�V���v'!T��U�X���E[�G�k.G$�ʵ?=��f��V�ۏ�.�-�U[�����vX����:�EG�:��dZd�qA̺�D�n����.oq�ǧ�3��~%�8z�<�I{��bk�S8U���i;o���.��c�#�t! X6b�u�c�buT���{������G�@ahǑګ�V'1C�j��e�p6&(N�y�_�lT���.f���	�zv�_�l���:N8��0U�j��~j6���ŝ/�3*-��K �`M$���Z��L.T�p�}�`�j�<�ֶ�����[g��KA�V�sF����n�|s⦽j�����wtTc����uxZ��2#4p�O�ϳ_ W(�/-z��rg۱~åq�ױcѻΌ�ϗ,w}ﭢ�fT�ީ�Ű�!l}?5=��� ��d!�k�v���Ϯ��!cy�?���;�-���=�`b|Zڤ|XKF ��DJ������-�ss����P�%z(��Z�_�<m4���n8��Q���V��C�h�NۋWx��n�Zvv���nyCLVݶoך�N�y%��:u�©�~�Q&�_i� ��hf��,b�`M(��nl�:!�k�Z�k�l���*t
��>� ��Q����O��{;dPX�z��4{z��T�L�u��gO	�l������5fe�˛���<V�0�~:N8���".���2-g�#�%'����	͐-`DSבP�o.��d8�rJ��������z�2=h*{��w�H}^,�|��KVX6��8D嶒V��������v�}ZIa:4��k�w�(-VdY��B���縁yS���6���m��H=K0=��vA`{�/!��G�A����b8�#Գ�1�.mv�{rφv�����.�1D0�-[!��`�8S�|`�(l �\��yd�.!�IMNѦ^~K�D3��v��fn���e+k'ޥ���'��Z���#T f����a��m�}��T##R��vd�[��w�N��N��E]b�������	�7��o<SB����rEZ�?�I[��ƥ̥y
�hw><^����Rs|r�L2�A^.�(�hG���K�P��!qs6g�q`���sr]�Sv��~�X��.e>�#�����ܘ�	�?(85��o_�_�҃6g�72O#�3���>1o�@���l�W��n.���%�(!_3,�C�Y)�k�Q�bƣ�͒)�r��P��c�ɿ]E�X� /eT]s���l�w�
��:�i��Y�bf$�w8I�!v��<n�.^S���/���]�<����q�Oa2OAS��HZLC�Q#��Io��������:�?�(��~�K�P��F$���� �ˏT
tח�@��.<:)��N��@�mq:�gUm���R�������r���\��ύ �d��b�c��bɄz��$�j��Sd� �ʅ�%<�&��6+�|�������ǳ�I���{К��ؿ�E��z�ҩ�2�&�9�8T`k��藳�H�Y�pT��i��D��?��8vb�kX��K���@U���ư�ϟ��л��=�;��]:����إ��I>�K�"�ҴMQuR���;�Z�yN���֙��NN.�>kPGz�_Î�pj�=�[�Y�t-���*���τ�mSw���洫�Q4�|�t�$ �<��E��-{�������X�pA�	�W���"���s���[�&���u\fL���q�ܩ_Y�[w��38;E���m����~��[6Y����!���xS��0�އ}���8&2�N��`"a���RE���G�m��!��3G���1��3��nB�	�T~��ym�]�E���L�Ǖ���m�7�cԥ�n����o�9=V���Sf���yr���)�8�7R)��k����	��%:t��ك�k��)���ʖ˱g'���=�/E=1?�ڬ�TڴV���N(SǩI���@Y�r����#�|FpU�C�0��f�koJ_՗���_���%��ٗe�:G S�f�����$��ٴ��������z�p�( 3J�˅�g'$�����щ�<t@��*V1<�/.�}Vy���7*&��]�t�c7m�t��a&֨��w����Y&�0)���d4A
J��s�uf���^�6~Y7�Ut���u�6�o�*�Z�*W��v\CXKZk*{�_��(TSs�S��7��	H|�*+M�����[I@��j9�+[���/���o���]��h,ֲ\f����^��~![�e�G�����D�'�-���:㎔D>�84|��Tf>4��w���-.��6���[��K��1�g��B�Q��{/H�1V����=i�Tjl������]'�]4"���g��3~˼���o�wh�d@ ��=�;�fE�%��Ү��CS�w�����P��=�Ad�,�d�]�E6+��޻H�����,w��aЩ0���8�~ ;7)G����-hM���8L�R-w�J��pX]W���׃��;~��4�r��ŝ��t�C���E6@�G�.�!�#I$#^(��`:"Fz4Ks�~""���{P���O+222�sDNN�,}�<�,{�" ��s��5-�l��=8;|�Z7��-��u����һ�!B��Q�����VZ��׸�ʃ)V�&q��y$��"~���\�1�\����n��Xl�GKT5m��_��)��L��	�bǧ�	���[_�Z�"fX2�#�a_�D���ҹ�p������ů}	(�e�V�l�
��CK!��J��[p��#�c5U�z8/�ψb�r(s?X�縆{���K^������*Qq�𸷫i� �K�D>(�$ˀށk������d�����ɒ��'m!)�����xܮb�џ����2�����&�-��\$uC�9x�����^p��Ne�@��̔6Q�.Κ��C��{�c���H@[���om0��
��S
Ҹ�T�]�.���C�|�hy��_y��o��3�6j��k8��,��.���md�|�LM
��������1ic��)�eL�f�U�L+ƍ���s������؉P��3!�TU��aA�`5��H��Wג��_v�xtd��g��@�]�V�3���<�� >�k6 ��������F�ER�ֆA�g��N������7�9�V�3y�O�B�(,���mll䞹���t�������N�z�Ń�e�Y}b�﯈�a��Lpي�2�ǎD.�55�C�6������C�m9H�� äk���g��V��&�ZZ��3''&Ft�Li�L3Tyz]n\��M��!v^�+��<��gΒw��ƚ+B^�)=�SP���t�Ȧ��8�R�������g��S ��~�ѵ�I��f�[���f��������b燅�����w�x+v)�FI߆��g�^�����}#?��t�mW�S���+�ˀ	܁���˄%W�u�8�X7�Y�8=�P6~�q޿!(q^"U^��c��qw:/W�d��� ����w$�����7��k%�Fŉq�e$��DCP��ɏ>=��/hV�H�^���!��#������ɏ���X�n;�;�����,&E$O����7XC�Jj�hX$<Up't@��{�[�k�̀H y�Ю��U�?���2Jv=�zY���PW3f{=���C�D?�ՙ��!Pz�+��%�m0���ևx_�	 }������]�I�5ei�́�2`|�R���7y���D�{-ؽ�p��Q�v0�{��r����9g�w�"_o�0῎q�&�mXA��?�/#j>	��|�I�T��=�"ims󽔫kL�w4|��`U�����!G}u~�{{�$J������?��c;*�U��D)�D��pʨzb������(^�'�n��L�����+�w�e����[��Qͫ}��eʏ��N�a���o�i��8t���L�[�U6	�M�Jc�ۑ8.E��vFv�Z�P{ލ��ʛ$,�h�s)�����a�)��A"a�M�D�j�K$wsu��\u����� @䧥�e�{2.~�b�X�B>O� ����E?!a��Q�����)�œf�r�%�D��t5ʍ��!@+���0Ŷ�_��&������93�5yo��5.?�Jdf��Tw& �ބ3�	��ً�O�x ���^-3j���.��	�P+�])�"�=Nr<�t�{�&ӡg��H������o�Y�r���m}���:*�=m�gA��U��:y��EO^�~���u�*��z�gpʴ�D!'+����G�����[��Ϙs�"�U��iB݁�<�~;s4�U����@�N>����"�)tq=���(Tƥ��rޢ.,{�3���9E����� ��v�������A�g��F8 P��nQ
)�R7ʆ�-Z�4��Ml�zyCX��/Z�Z�-����l�,����\�ֽۺ�*)��Z�n��G̝L@����z��D���s�j�5Ա��R���I�\�M�T_�w�%1�� R����q��[\pwܫ�Y}�Y�������2�F��Ӄ����z���۳K: �w{'4�g?r-�n���3�m�� )��]�$�$�;��q�w�>sͯ6[�t��n~Um��:��_(�υۻ����>e�שmāsS:��f�����ln���O���5Ð���h��&(����<V��%~�3P�&f�L�3=k E]Ƀe�5`-t��E���ϙ?9�*�ƦkOPx6\��!�QHWۆR����ꓷG
-煖N�Ko~��<~��_��x�!�ʆ�WV7~8�

�7 D�ڹ~��:$�h�?��r	zYXP`�F� Y�t䢹�B�|�ͻ5V��>�M!FĘS�����bycl��}�ר���⭬���Y���@�o���o��>��M�{���	��������	f>��ݺ��a)��zZ�%�Bfgf��VGj�M���1�H������-����*�_��f��`|3< <�RX�&�B�.X���m�:��j}.��2�}l6���EF�b"x������]����-��][IjK�`)�ۣ��[+Ɓ_ۂ<K7��{B�*�\N)Q)v%���Q�3��P�4U���/dc�̹e7��;d�~]�ow]0j�z�h��s~����?�\��"	J��ޟcO�o��/X����/v��ݑ˅�U�z����j�j��NAvU�k��I`�� �q�.d5�X';��0�zҸ�s;�Kw�:D��YRt������X9��ZN.(+},X��V#��\�ˋ�B-Қۘ���T�"D:�5���<B˪�b��:��=�_ۛ��{&&ٛ+sN�H�L-��?33�/����k/�H�8��X�bN���Χ���7���s~�yzf,qa.8�JVԶ^�����$��^����Q��/��&�vN�|q�-�tuX=s�J6Z��Ø��.E�H#V�\�÷�̟�"^�/p��g.��``�
�%Zm�C}��w�ծ��̪é(����G�-���S��=�8&)*oV�%���PY��a�W�R�*,�&~p�(�ji�XY�$ph}�>�M!'�0K��f!ŭy����:K���x�l���ղ+�a�"5�;t�op��o�dAH*���(iጠw�fٕ��7rT@aÆ�u�a����&+@�E����#���e�ɣ)_w0]%�K�[WWaD2�����r|����\��IE~�jM�|�w��,����V)����h���_Yci�������I�TY�v)��. ��<���Md�BΩ��]2s���/��E�'Mf��/>w+��*	��_Īq�M؜�ܲ��u�a��I4ׂ*r/��4�ϑ��*e��q9ʠN,�
�+��ly�L4s:1�x���Ñ�O����챃浸�U|;=Iza�6&ح$�R�^/�<˼w�0�A��M��J�?@F}N�gTw�P�]�-��{˕W�$	}��1��)��X��5�l��u-R�}�ܒ`�����r_�m�1���``d���j��Ac�A�q-�<i�_�<���js�:K
��T��hT�*~��z� -�Z���@1�Z�.��\?בܶ�uӡ{o��1��w�4�)I�k]����$K�a�3����ǒW:��:�O�t���S��6��^�n���J�8*�>�"�;R�㙨�)��k Jc_�r#�׍=G�k�#S%(����0+�))Ãgf�ߣ������sk6�6��
��%��׌ dtf�ÒU��}��N�
�{.���t�3[�� \��S�����Aַ
�*y�d
~]�u�@����#�a��)�l��@�X��»/�a��޹��qy��b�I��ӥ#�
�{Q"yd�3�FAZ7�G��80�Z��vƣ�C �\���^r��ݎL�/��a��:�SS�+��;�$E�+�̮�L�7!x~_u�k�%�/��z�iF)ד���$���f��"�ܛ����p֛���7�5H�q��_�[G]k$Q߄pU��^,}熒*�z&�/"� %��OAx�N�{ra�|�z��l�l�}����qĚr!�g���(X����h�B�bu�h�r�{�i�+?�nU3k��'X�.ZztHkx0_q]o�����ÚI?�������:�o�=%���;y����]$��#��S%c����&$��z�������D�_/C��VJfa�-8�� ��绾$N~6����qY�0�WG_�?Na"�"��I��s���?�72Ȼ��&�<�-��L.��"���=2$4T�i�MPͳ.����/���є9��;.�C�E�8��~�Y��62���k�?T����N~8.��8B��~������'�gaR==^+Y�ׇx#�ƅ�H�Ǯ;=5T'Z�+Lgc(I"\��© ��W��G�|e�e��[���Q5�#e[��B�X��ɹ��A�Cc���*IW�}(=:V)�Ol�E����b�E9b�e%䲾�%%����������,
��ޑ�2u��1=�EZ/����[��Y��G9��L{`ě�F��C6�K*���{?I,Zya��A|���
�kX�aXa1��uP�*����|�c�l��c��q�'r���7>!�th<�~C�="�Q���'wU%=ÁX't�g�
����Y���|'/�s�F�x~I�{�˷���څ�OTV�*��t��>c�QZ!f�6/�?<}eX���D���;i�AJ���n����[����;�A������\���3{����Z�F����X�*qf翩�xz� 9ݿ�X�A���lqP4�<b�8�P���Wu-4��������nN<=)Z�����!����F� {M,3�i)TI���Vט|��:��f&L�㚾�4���X��'�f�Ypp=�H�������:�0#{	3�g�9z����:8�Z�i?�>���2�4t�%���w������_$���XV����4�MP���㳫�;T��J�Wl�!TS����٧Z�wpʓ���� �g֔�?;�[|ٓ!���>���-6u�m=��^{���h�/�/�{.�U����
m�R%�YH}����g�n���Q�܆/��]b�2�!.��I�bi�b����������?гe�kvL�e���#���=.���:��ꝅ��V��m��`��<���~�0��,��>�w|��㡓xv}!}�֛DP���1U�aRbF��4��a>�pŵ�6G��
A>8�;��K+�u���F͟���,�c ����������+�S����g��ݪ)%|{���t�K��|��Z���F |�������%� v:¡\�T�m$)���"$κ湗p�9'-y���*UtlZ!�\I-�m����N�&0ߔ�ݎ�=�	��`3���adLJcy�<p�� ��P:�`!���et���B7@x��;�O�"Mc��0BC-RiY�%�����|{�[	��W3�,��F�&s<�L]�dn ������f%dR�喯R�1}h��<Iv��	����%�QfZ�����Z�K#K���T��>��3���o��ի���=�ߗ0�����m����~7U먊�>�=��X����X���LW�zM3]�LE$[D˧y=����ԯI	wI�Ѯ�߈�f����D�]߰mm㫜}w#YJkvڷ�P ^nVш�>��;n��QK����N�'V�z�5�m���}*�8r�m�s��*g�w@?@I�z�O�WpnϮ�u�,��{�I����H$� ��0.���D@�<��
���O���&mk�����|��m�g�w�=*��؜��P ×*��Z�[��>N"1q�}���U��@$FX닥o��@�R�>%��mk���`�,_q�Hr�%X;��Q��"���).}{�OZ���e��B
��Keq�ϊr�#�?ug� ��Xh�IJ��&5���c��aW�N��\�Ķ '~�BD���r�ct���#�G�*�,M$y
�� �~���[�������Q����J��������6X
���ݶ��߯|MC��0 /�����C���b������02R��-�y{�����? �o���jh�)�8-TV�w�@�ks;�z�q6�xH��;��:bL$�d��B�eR����>�Y�K�>_���k��	財�D� k��Q����==�ÿ��|:ޟh��d�SL��o�k�/���P�Շ?-.�y��^�\�C�E=�ҼI�K���s�����r-�T
����?�f��y�r+~4���H֋xώw��y�{��s�F���ϸƁc�Q���(rA/�m0~�ɪަ���+^�	�/C�'>�KY�!���`��>�{\?����KDϩnz{}��HF��(r#O�J�|"A�_���_��� �4����z�ֲ�����;�d��Elۮ�2�¢F ���|P���e�H���1���6V�u-�Me� ��#�{�<l�eՍ����P�ϫ�
���_�o�QS�B �l��4��h�"����,�_=,.j~����I��!iD Ό��8�3&�������a����ۥ�Ʈq��% �KC�A�BPH8�L�O]�iV���‼���V�K�,ju�x����R�f2�z�wC��2�������\P����Ւ��Ve|*>��p�w�j9)��9_@�F�7�ӫL�6�/�DWh�������\LD�6X�Y�ԁ�������nf��N��x�p�	�aw$ʝͭ�v�\R���CL�~T��
s��=��S��tإ�>Z��a``PTV�g�ǃ�P'����y��/-RM��u�no�r$U0?Fi¤%pp*�%�4����raQ��!{%n�t���Y�}�v��&�U���>�k_ ��ST��ؽ/a���/@EA^n�ګ஍[�t����߿aqpp
srD����c�N���Ҹ���
I��n�!�>w��e��3*�JW��AӼ�hoz[��k3tR[́��E1@$IY�$t�K3f6b�J� ��k2�����MvЩ!	(��������2�G����>Y�����yb�����E�r��󵎦�I�o�@�X�kPt|��ͣ���_|,
[3⁚��~.Z���X	�k��[}d��w���Sa��3����*K����ì��=�ĳ�=�/8��<
:$W�ԇ<�x�ч��7�Z�'�}���&Ed�Rf��5xIG4_��h�2��m�? �KO�6��سux|�a�VE���Y\_�X�W�q�Eć�B��M�֒��ҳ}
 ���l��E��xS/�/NH�LQ/�P�A����Q�R��daN;�()_΅8��Z��zӦ��oc��"�}�a�(�Źj����&�H/��i.�?�U{8;I=j���F)�;�ʖ 
H���q�FZ,DI���9U�(��I>f�ஓw#ɢ����?)8�5hi
��V��ᢪ��1@˼t�]�@Hf���#�K6ݚ������6�=��.52\��O/�A�U�����\	��D��%�e�wGVP��/����dK�E��C��CX����Q��ƥ�Ͳn�Fhh,)/IQE��
W���_�/�T޾tz��9�{��Ę/�Z�۳u�I�j'��T-�u��;se����_��r��>R������ s�.m�^���ƍ�2O��Eq��E�O~�@k:~;�Uߥ�ݴ������6O�\�]�`�H|dN�I6�#�k���fl/}�ad��x��C�_�"�Pg�']��Oj��	w���\
n(�%��/��Ғ�_�/�;�g��Tf����v�7˒1:���:�����2L���^��i�ϊ�̪�}p�%X��O�ۗN��$
鲍�*��F�^�5�(�r��\z��D\^���|$;q���$��+v������?���
���~��aTf�%O���8���D���􈝲��s�ٛeo���:�ƫ�����u��¨.�-jCK��i����$=.=]�������.V��a��C��}N�w�*��9>��԰r�j���(*� �-�ܒ��0��n�� o��ŶY*����b߉	���}�24D��Os�!
�F��e���[$߼X�C�Ɠ��� {%	YwR�3;��yHЀ��b��Z~|<SG�\j[ND:��g��1���Zw��g��&�޼�w���lX�j|�΁�oIZ�+����sp,�j������,��(w����D]����5q(��&Fj��.ۻ)�܁,��� ��#�m�����t5nD����>���ޝ�����|�..�})d��eh'+QGo������D#���/��W�����*�m��6���ҵ#��~9��a=p���;6��3ߤ5ڒP
�%�*���n#Y�O�
>�����"��V�VĆ��}�V�}�չ�)��"l5�NOi&nr���K3���+u#��>H@X��K[̡�7��!� ��	�.,��gCG�=:i2<�U��\X������lz~�5�`.������� t.��t@���p�t�\!@A	��L+�w���Tv��(����Ѷ�E)2������)��DPDr��r%i�P���!6�(�V=��$��G>}��;���Z D�%�jh"�@1��:R�?c������L�����f#�8��%'iO�>�?$djZ���;Q��A���Q����.{��X���	{�r����0���U^#]>V�|N�qd����n�m�9q$����_&Ja�/�O*t�+�]FvtB�u����}��@{(�8��u�(��M���Uehf�54_��sAh u�3�t�=}����V����!=h����<����`��mAߋ�*a�/'��F|Mm�`P7C8�� �p�lq-.7E���=�yq�]�&&[�׍d�	\ɓ9��g�@�Re�2ܜ�9���|K<�p�QB��äh�}�W���Bza|g.�/���7���ș��(}�j7�0Vrww�g` �����Մ��t5�����	������r'��>w2n��JYڴOx�n�77@���S:]�\�1�Ng���M.�_��?�ݺ��G�9U�$[��׈	ZLE31��G�omLޟ?\�T�A��
Ȩ�K���q�siQq�Oc�
�=K݌�v�rz�l�Ku�>|  ��2,
�	o>6�}��16�ax��VTW�;��t�%��v?Tckk�j����v\�x��G���͏f׮��o� ����L�^[���\�:S{9���:�B	�~��IB1DǛ9�I>�`fT;>��E�V+�p�th�r�#���x����Eܑ�c�����W��مmj������d���t��ZL�lPo4K	M��]m�N]8Mqn�^�3_V�DQw,�.����I��<Dn\�N�����[w�Z�G|0�2=�Y�Fd#!J/��PSU�O�$"*�м�;i�� �;����(a�*�����v����z�r����CjvSJԍ��g��ǿ�Lvn��RnϘ=��l�^������g��죧�Oڬ����O
}�m��	�t���&l���i|��8�$9�<��}%��U	3���p%��xax����T.Qe�n
a,�Yr��M��}3��t�C�����}2��>n��Rn���\?˕�L1u���.����O��v��6C!/�:r��s�#�g��^�oOoC�qj�F�L���W�m�\���H^�N6c@�Q�������*���c6���`��$������̩�����[�c]n��:����$@k�|����t>-��_�����?�~C)�;�����l�y���J���W���4�}Q��D�}�Ѐ�D��:������N�n����5���ʟY����p_���|z�_���}�SQ���2�=�����A
�?�.1���-M��R����:��M���W?����6܃����8�n`�]������SaBβ��3T0�-��T������:ggٜ����:��l�Y�>� o�p\4Y��2�Q�p1�a�IEs��_:q,����:�v ]t��ˈ�m�A��B�����h�.]��$ӛIǷ�z����`��9Cc)�/����zs�ٖt��ا�/ּčg#y��. �-9{u���E65m��m����>l��/��T���ɉ�U>�x�;���Ʈ,]�,���W�����MBD�dYծ<tKE�lZ+��{�&��y�k�op�Cc���O��1V�oCh��q�uh�30�Om�5.q�$�S��r?E��U�=o7ޟ�RkZ��X?H$1
�֋��U��~��>��>;��j[���j���KU�٘vV�������V���&�4�æ��W�h�NX�`�Cb
A;�1�*��@���i�&�4'���X_�a	fW_͠<�jy��Ɔ���,j��K�["n���������Wn��\��ŴY���v�':=6A�P�x���3	G�h>�\�xe����ؽ+��;�'�T(����7����n�7 Fp:b��./�T5v�^�F�?1�O���9~ �f�;b#fѱ�2�<u��ଞd�A��9D�c�f9j�P�_�+Z�=�N�d�U�9�=/�KW'����T�;2ap��g_$�[���G����᡹#	�2����^�=*젣�N�͕Ū�O����p��T�U'h���u��o���VW�~#�Q�ے&�����ݎ�}M1U��s����Xz���y�Hx�"	V��0�Y�W.W������yxC�"dF��EkBb�����v�d�)f�@f���%	i��Rjm���ݾ"�@�������C��c�o��kbTK!���)��p���e�!�����Z0t)O�\���p��3��|�B�2��H|�p���� 9�i<�s���(���[u����P"����I	�����;>��{\:���у���Eo[��_ 釵^��αz��ڳ9l����/H�����*=N��΢�i��_����ʲL�
��ـ"�qe&"�52�p�?�:�$��[:?�t_?>�ۯ�;
R��R��Ro���7lZ��/��ĳ�]�MdL�N�Q��@�S��7�ۻn�� �����ǽz�����m�=*�R��?0���!����<`U�k� �n'D�tl*��������<%ִUt�/��z8�:����ڈ�L5tϝ����p�C�����"��3`�- �8�IW<j�t��泇Lۓc�A�d���!��Z�!���.R���ӛ����M�Ҫ��A:��-�H����-F�3�OOP�����qF�uEe�D�x�-m?t������d��,��K���yu21��(W�dI{ffm!C��i ��~�A�us����>M�Z�`tн��]G���F]��r�7M>����&�5�SOZ-X���9����R�2QlwGM�[�u���Y���T�5�wx�;7�9�\UJa3�OKb �l>#@/�g*�b�ƚ�ʮj���(�_�\5�w�``M� ��٦��8lC�O�y�����|�?��鞚�#��s������g]���
s�ǯ�
u����	�ѯ~6���%k9�f6lF�.�!xN�#5���Gz�o��N��[uR`8�j/�]n죺t9����V�L���!�fˀQ--�����d'��W�#�/����q=C����w�Zt(�:HwW'����M�޻��e%�<hahǮ?�6M��8�3蝕;���Q<�K���/���JR���~���Q5E�eձ�q �pm� ��e
/}&��]?�C��׽�1���o��X'�EW�OW�f�E�#�_���)8�+|MeG�\�7�l�z'	s��֧i�W\���=��]��h���hVI�'�kƮ�c2b[�B��.ν{� +_�nZ��.�ܐ�K되�w-�v5�K�,�%Zc�Y�h��4Ve5W8�9�e�%����\����A8L�L�ȵI�>�Lz�E�u����c�@lB��9��� 2����D��i�E節�����w,�5�`���.�#�_�u���zZ|��b�k����B�b������v�����"/FT/[���RG|�j��di�]1u-ݣ:�W�HJ�>��YM�y<J��h+M��s�����=�'#.���v��$᎘i�B�6�@o$�zҺ���Ҟ��r�r���R�(���8��5�:y�e���i�
詏����T���)b�,��Q\�
l9;ui��J�c9����c3�I<�V�Ҭ���:�� S�=��:����ᓠ���+H�U�)��zgb��Q�������z(V�ƌ�G�m
A�7}�g�<XW��d>�y)g�aq�j;0�(���%]��j�W`���e��OuH���ت{@����S\�r{Uü�F��E^���V|%r�u�?��F�+\�ʿv����f^ ����p���pW���{JƷ�C��W���cF���}ff�)�tפ_�N���Y]��(^@eJd+��>ߍ�S�s`�� �u����*���d��>�"�pu�}�#o�eؓT���w!�+Yo���4?���@�h~�Gt�{���SH:��2�o���B[��4ulz�4��#&S������K����ׅ0���t��>'k���>��6���E�g��O��7���fk.,�q�v���B/#4=T��n@�c�J�`�?�վ�#
���}5A-��D�[�AM :Ah&k��C3����m�]�A�P��@����p� �FQ�0�_`�����d� 0��_˦��+�~ب^&憗&bgI��J�:��ֈ��Lc{�����^ ���s�����^���������:Wt㵧G�j�al<Ir��^��̗�]ӫ�`C�i�f�6�lՎTe/⬹��$�f2�:6#X�S2��a��ɣa��re�D��Z�����H�ylH3&�^�z���-T%�ӟf���)!��@5��O~��JVf����c熝+1w��	��&y��i��J�n�z-kB��m
��Y�ވ&��_k�T�L�:׃7V�����=���ٔ��]�n;��F�Xb.������8�i��P00kY��@v����8r`7���[�&��\䤴�>"�l��Q����A�.�R�w�b���Lѵ�g��v���xL��8�?���]�p���b'u(V>*;��>q$�v<�ϡ1سAoJW��	�_s~��J'+��X]o�Ϣs��6��Q���L'�Xu��,^��;���l�i��lv��a������Ya@���R\{n_�-nT(�fdx�6˱�����Y�i�Gh����B�g��q�{����dEw%���V�޴�3��n��8����1'���-=9�E��*��f����[�bL�ӌv�1n����i��x�Ҍ�,(�V9z�x�8�l�E񫟞͹�9:���4[���fEbn=�?��׬�m��t�+�|[]Q���s
	Qk�(%H�Cyʤ	v�<�-i�fv�D�dfނ���\�\�K_0$z�ʥ����AP���F���@�R�����+7�k��G5�wa��~��r��XN��(��-ŷb�����J��w��a�;/=�����U�����W�9�O��B�~:|PMpփ��^�s҆��z���'6���]���to�8�uǬ���'�y	�x���!���Ӡփ�lͶ�tڙ�`7�Y���_���
���,�ZGv]��ٖ~�-y�.T'xZA{l�Ma�u���s�nE��d�iҺ?)-�xh�ͬ+}�1��(��
B�zO#!e�q�S�eY�-��G��ڒ�e{9B��Cߘ�-�|VZ��x5q׸)�����7�ؿ�	-���3�NE,���S�$(�m�d-V1�g5������C��	b�7�`�DX�7}���Θ���ho�Wܚ�w[,V/���W�
�U��FL��뮮���{����9�Xb�L�G�M��mD�O[2ɒ�1'�/��t:v��}f6�( ���[Tl�i�eg��F�J>k~kT!zbe�p	��~֊U��Rm�hs.���3u���r5N=LH&�LDp;!��V^	wݬ��m'���k��h��_���B���?�$`QA����L�9�8�7>'I�.���*1E�r����ҳu�
ΎP��#z�7�|���ն�R�mǺ�f��b^uab�4;��h�p��MH��5��G��v�q)nO!���'_��=��Q�ܵ��?����8r����B�zK��(hz�dd�7��c0��Y/���R�g���f7�����3k�����þ���O�k-�D����04�란����}���}~ߖ�� �cf���b������6��nD���7�E�
�TN,�Iʏ�f}N\�	�O�x���L_�R�:nV�!����@-_�b�I�������䩳��=�'����bg�8�t�[�f�,�Ԙ�O�:�hW�:�!���C���N�D��*L�A�����W�G�Qi��Rh/�D;z~:ndDX��N]���Qƹ�N�mX .�AeMs5<��Ed�!��e�?|bZ�/�E�U�����4��;2ឭ��
���%!��f=�H��(>lh �t��8)���]Q1^�]�#>��ۿ֟��~�� ���4[��`��?ھ4꟦\Ä���ϖ%dL��&�
' �������YA�[��S�K��&r���S�ğ�k�[�9%��~�i�~%s�4१��_�� ���ao>)�	9ݼ�k�*�U`/�0?���Cf���9�{#��N�E`Tc�_Z��V%�����J���ݜu�=�3ޮb�A�O�ֆ���>=�R�2L���
�*�̓���	� �r���~}� ���ʜ�H;�=,�m���`�Ȅ"λ=�~�:����}��ykR5/�[���v&H�+�.(g�W�n(����rE?�X(�[�Vȴ����$��/��V�-�
]�[�D�E	 �C�x��xo�!  ,���+�Q*���T�e�ֶ�a3[c4h�Nr�3A\��i)N�a,�ک~����z��|.K$H���GM���o(p�O6ܦ��q�'B	�c��8}�"���,��o`�M9{��*��R�����ǟ#����xұ�l��1�;����ء�c�K�e�����tϽUd�7��]y�Ք�>�l��[}�4M*��Ub������>�{��My�ٮ�}��R\v;���<������Px3v�1����~s8��n�4F#H{�&Y\3䍰���/l!㟮B�_���xIjq�'�����Sj�luI3Mc՞om��֨ut�ސT{�y���2k�&?����Ð'6,sb�a��`���U��ӼmN�ʞ�&��rB,�w��~������I�x����h��|��nI�dr	�2��6Ӊ�I����]��d�?.�3}Y3�c��g���?�h�"�H�R�������˺}����t	�]?DÚ�g�3� �E�;��Y��PT9�
���,O.�X���g��`�S�3�t�u��#r8�rk������{�0�;��QY}�'M�8�qxb���� ��G޿���׬̮j6�8*m*�>��w�t�@R8�����#P! �5��^;Y�*�ǲ��wO7ӆ�!�ؠ�[5?�} usZ�0-N��
SWX�Lݤ�$'h3���'Ss��f4���Y�i�A!	-,vkv��o�� 9(��.-�e�/�������f��$����u���x�F�
l���j�J��jM�b#�9�^=��M@��]���2nhX�$=*�^T�
��|�[��<��z�~N���v�M�_]���V�~g֕+j#]-?wl�ߕ��7�[Wȏ1 ��-���DMd)��~,�*N�;h#!��̬-kFV%�����M�l��m�7
�/ֈW�����6�ZE?����-�c݆�j�E��V%�_��.������ۉ�hcp�N���	�ظj2r�oen�Q���F�� HՇ�;�H��G�����V7�nM�q%���. ��"�J�-�D!/�o�Z,0���E��tƙ����e�l5p��C 8�m#<�p-zQH)��P/?Y:����[c^=�ا���6��d�4z�)�~;��M��aDpǱ[B�w�R���+��0�]9p I��n0�c�ƻ}�����C��D�����E1�A��C1��u��d�!�V��q�7��`�4�yU:C��@�����`��D�x,O�F@y����V�E�{
$\YA�}w�n���Ӹ��h�V�� �ȯ��^����s~�?�a��=RRW~��Ǥ��.��c͓�U�����ʝi������K�����s����#�H}�4�?[SJQ���5�b�uN<�{�xSy׸�O?e[w�pI���x��"�kÈj�#J���;6#�G����l�Jv��1O����Ȗ��qkq�97�F-	Z�F�m�� ��2������9��टnE�(\$W�5�Mv�gFkwʯ�T��Rkj��s۱x0@��z+�؇�a��T�o��N`l��5�^��0uG��͝x-�=��!������-
E����A4��%64\�g�`ubz�{�2�:8��p�1��
�=��sQΛ�����8w'GYT��et�6"��N�Õ����A���ϑ\Pq8旭�����f`W������Y��t�|L�	���s�k~���k{!44�KF�)�uY«������K�����=>����n��;�1��5L�G&� ��Zf�Q��e]��-�? z�ʬ̍�I�c�Ў���$S7ҟ�T2
x���{��\����( �1���@�4����W�W����޽
|��}�����TM�� V�tS�{��qXuŤ�.I�M;
m�gR{����0!F%(�nF��I�fABojC�M���9u�(�G���)�U_��[�~aqF�;��ZO�� �Gm��kp=��J��J5��-}�G��Ay��Ӣ�kl��&�"����P�6�v���#�渣���.�NHn�����B���d>}Ι->W-+��H��C�{��[�J���[l3����h���p��5{�߲���l��U}���,��Q	�C��&;������6r�����W$������fY\��enL+�]�z*;�������R���X��H������,�5-9p���B��瀵��Մ��G%c��`6
f�Y������R�Z��Q&y^��y���߼�F)�W�@��ux�?��&u&\�\=]r�Pw-C����@��R��� bÒTPgLwT�\������O>��7���I-&�[�m���2��N���p�֣�~��a��nl�N���U�����+�k�;x�vھtO�w�\k���*q=��ۘXPR���..|�b��M��S�s���X:H���du�\��'����M)������O>Y��"\R��&�m���I�P?r�'�,�n��(��R��;�)� W/�9~��{�z�˔�~\��:�����`0:���Nw["Nw�"Ƈ�qF(:��-m�-y�?f����(�o��M����\b��
=��a���g�3���ƴ�q��Ϳ�.�9��f�,�,��~�A�,jcOC
������y;_t���Ͼ�IM�cn;������O>����6+�� �V�*���t�o�h,,6��p�T�ꨉ`' W�|�9�L|�r)�v��G��C��	��::�����PL�X�3�B1�Ɛ�h}��/E�[�Ӣ�J�~�
��B��c&�	5��V��3�Hzs�j�L�B(���rp�x`]޴I��|�1,�2����-g�1
a��8�`�%�tzz����`'�P�q���}T�c�$��䊑�Q�*x�D���'�G0���d	�r��y/;.Eu#���?5�6)�)�� \O�xR�v��L��I���:d ��z��(����k.5%�=�����ʉi�����j���������j)�tG9�'���+��\�KA�.��!��3�NG�?XYp��)3�>~�򻞛��6������/[KQO�/�<2����ߟ����� `��z��Ֆp��sqr4aq�ߓD��~҆�8	;o~���Z�hX������|=�'�x8��6��古{�S�N���%��~i��_[A�H�zBF����M�7�-���9}Q1?EwQy���O�<ϫ�F�S�uz'13>�y4te�SP��ɏ�J�}:���!�z�&���N��+� ���~Ո���Qv��$��K��ꢢ�Q���g���|�ybK��jH�X輴���>"	Rɂ�]�r5E���|���c�+@		��Z���iNu� "�����[.|u�{d�9@!*�*铋�-�i����@���daOT���������/x�)���Du��`���⻠��+��g��&�cf���:�OIkS�Ғx ~"9Bv��)���9�������Ȝs��#�]�*�D?	��C����zKVxz�󫷛zD ��e���ء�'���)�)�L��p}�	�#hޣ u��f�q��o�� �������S���F��	��Z���m4E����Ӊs��G�s��E��n��ф(_���lV+�/7)k
�j$��10�ߠ�)!���#D�e[�t�(#��^ca܊������{��!�,����x�)�J�c���+��T����/�=8b�h�*倰� � �+N��
.T��.�}�&�0���(�����Q~ha�w~�3Է�1
TΝ�Tֿ�)(<�Y��D<b����Ӂ�s���G�I��,��h��=��@*�w���(��;�����<zȎ�Dݗqe@ʋ,x�UPrg�x�~���&ƭ�y����p�n��͐��M״菏,8Ƚ������ �v�j�j���:��I	�}����7Z������K*R�l�Tg �[u�:m�%>q����uPo�1���[��M���d��ȁ�3�0}>|��dI.)ʩ4�*�R:�=�V�}���S��x���0�.^7]�'�¥�[[b�#�fr**m��Q��Qxab1��	��z��l��.J�R�?�m�7��q�#ܬ�&ׂ�����DG�5oD�K�T��G�[÷�`LD�s�|����������`�	���[�2o�r_@��T<�a�j;ޯZV_ �p���(��kMc�(�G�G�Ie�o��/�!��y�ն�� �`vT-�N�Nɺ` �؏	iS�3�,F:6�~9�B���1�,�����T���Պ�/�ȿ��7��0�����4	M�SP��͓��GX���}�Ԡ�9,5���l��q����
���U-$��$H~�2�q�A?�|�𒄢�����w!�~&c5Æ�N������p-u�~"�H��qʢm�Er��h�/C�����[�|�-�Q����5 ����ҼZ	��P�V^-��3�3�A�N%*��� �N��i��.�{?�p�~������(��?�br��KI���ȱrP�S� �$wN�ݞw`�G�ˇ;LG�Հ����5�|!;��n��Ҽ���Zm�EV;'%��ʼ����+���,/ߚ�2�̲�w���Fj�>>ʱu�<�-[�v�\�T�l�"��81#I�<!����7/���k���[x�w,�Z~�]��G�\��f .���%��\K��?&��/"��Od6�)�����5V���ĩV~�BM��7�-��*f��"�	����XVli!0z�?l��T�u���G�/��k]��2�$��������<��k��S������y!u��NZ&	ZK��9V�}�&W��zl���@�����
��;��)(]��'��lf�V�S<�5�h�8�:�*o�������W�ְy���0]�4㖕�_ɠuƆ�i�`ΰ%���Q���d?8�E����?M���و�J��6V%�Γ
������fuǍ���8��(G��b���[㡒ZʌrYF�U2�2��m4/@���%ݬ?l�x_��h�^��ʡk����[��OI=9p�.`¼4�y�G�g����^OA�C_�L^
�a>����ptxq�\
�:�$�݇xm\�b�b���聁A���p>�+��#��A����-����- t*fծ�u�'Gf�)���5mE0��N��(e�ZT������ *^J��w��1���Ȃґx�e�++��jc���ik:�EA�G��͖�=|������7��J��3`�=Q��Z��D�ѳ��˗�L7�Is����p(���X46�;
�z�ݡ[\�(��K ���XT%N�(K��������/���Zӕ&H4�A�N�D�{כ#\/_z�a݂$�
�/�Bxz��!�b%<ρ/����_��8�l�x� u7�xx�;�W�:GZ��ma�}�
���D�Xo��x	��w�{�7w�S�OI�U�Z�/�D8�w�nQ/?�2��j*�.n�C��Z��(�\\t��i9+pѐ_���%��ы�PP�:�6�!7=5�E�Ꮧ֪D�@h.%6h�8uY����[���
T���0;w���f���n�&k��)n�E�i�ji�
�"���]�&�v���z�M�E;oOL�{g�N[X�o�X|şv	��
���gR�m
P����:hc]�:����<��?���uL%��Ϙ�U Mb�e
���c T� \���˺����2��P� <c�A�H�e��w����n��r
$�/�K�+�'(��}d#�s_�%�gk�xU:�P)n]�FD�aYx����NC��Rm�R��1,���nq���W�Ztq��a]�d�w�h,���\�gz��@���\���t[��z/������u���r�P��xԫ�d�wY�֭4�D�9?Z�Sȥ��:�W���l ���f����b�v�&M������5ym�L�3:�\/ �~�F:3�`)�,m��k{��n�}]>9$D;9%fj7�u��\\��\��^���{��Gvf�>_W2��ȥG�V�l���|-~��@2�
��@�ͪ]������|SX T�&�dٿ�o��D	D���\��O}��92�9кBQ�#H�؋	�Q���IF�J\-���w=�9w"�j��"E	?� �����ea�os&�Wo"�W8���%ǘJ��H��:w�m�C��Ip����P�lt�7�s�X[稀o@�IDt����J��_;�C|��|{�@�XI�D������g\�YB�e�V�D	�'�FZ���Px�%��"g5�Xݗ�����f��W W���9�x�?�}�XNǣ`�y���!��B�z����������[�bM�-�����=D"-L<�]z���(��o�������@����	�C�[��:�]�="S�т�S�i��`��	ST9W��Vo�Eߺ�H#�1��nƧtp�U�=:����Qع~*�^#�ɚ��  7��<���A*<��v|������g6j��!�_֐�LK��-�/q=VD݅[�[߻��L� HY`aX,@��D8�xm�������N��s�#Q�{���!�.;�y��0v�;��5�Ȓ8�[Bd]p~v}���Uk�J�;����֢w��D!�zz�:��1��\�3@�.Rɰγ�?)�C"�����	�D����,Olڅ��i���Ղ�`3��řJh��'��ͻ$��;�:�����j#\����(m�[q�"�Jp)�R�8ww���R�@p��K�w�9��ܜ�w��٠�Xp�)���Kb���:șY����]�F���l�eΩ��ܴN+%�`�c�̺�Rr�f3=Q���38���4NŸ�Nnƕ��'�Ǎ
�ñ�Bӵ �8i��~�䓯7L�Ik!�q�c�E���<-"Bz���@Q�&�*C�/
Ι�,TFj"��ik�-k܏sx|��ݛ՞g�/���7L����A�ƻ�^��+=N�&,鞕ӣ��OS�,�]F�����gw@�y�:�h���ޢ�P�6�2��Sc��� _��͚��d�k�W$#2a��c���#���.#[A�:�R׽���mo�i�n$Z�̀���5�����P��'�F`i6EW�D�*��@<���	;�v{8�Q�ǀP>)��;�H�L�kt{w��d}g0H�5�h���x�(kI%Or��׭2�	��x���v�d_T�����+(W�ؼ�������tj���(bD/@�b����P=�6	��0�RoT���ϝ�e�*\�D�#�����7�G�!�UIn�p�^0Q!���!ZO�S�o�ZƝNV�N����B��C3J���v��%��W�p�6�/�QI�9>�d:�m8[�?��01�SȢ�U�/(��e�3�V�e�����e-���;U���Z��Z���ŃGJ_����ۧ�;����4|�Ė,����}M�g��8�T�p�ב�P(���#h1��Ԋ��:@�'T��A�/��IO��qZV�����G(q���Ʉ� �)�E>���TE��j���6k�P��Ƌt�.����-�>\�ZZ��2V�������_t;j|^�w7E*��4����ϾyWJaV��R����Z ��^����h�g �Ť�x�EMt
6r�k�
׾�4Q���W]�!
"d*bt(�r�Sd��9�7p?t�r^HUA3���=M��)��u8��I~�؃��Rko��������b׬�����Me)��2�Y=�~��8$���0����|�#�[Q.���o��C&��+I�4�&�����_�@���e�|+nSڎ!g��[jY��� �?ˣA���914Գ���Cg��
�HQ�8�h���2��P/鯯�_��ݻXs���q�7�_���5Z�Od�!�㼥����aP��&��_,�M��q#+�)��/���>�%��uXL
���r��8j}I�d���&d!O�ٗk{}Vu��UN|�`�A)���C|�2)���V����'x�$OKkz��Z`%��K������o.��W7W8<��<�]{TY� ޗ!A��)fF�V�^��l�\���酱�C��X:]Ƒc>�\�뷰�Җ_�x����7)�^d�җ���W��l�J���rW Ո���4�~�I�<b+�3��QD>O�����"�/���{�ZUUtY�����\�+I;��d�2�R�؜zn���&���+��F��,����'�Ks�i\�q{�i���AG�^_���%z_厱��^���4D]V�z�6E��|V��0����=�|����>M���1V3�������j��m�yBDįw���t�-@�ɃkG+�H,��|��S��b 2(׷�2@F�rRJR��Ԑ��9�>�x����$��i^����Aa�}~vi�����8���w�p>�j��ryJ7l5Rlq[J�u���Ara�*-+��>V:|��-M&@��̂?��ae;���VW��{H�-a���q�VDz����gu�鑠��������Å#L��`�f�wzy�ɯ.��^�6��p���*��*�Md�J�t�`x��.�z���k���-~m"��g��C�����І�)�������.Im�j�f�c�s7v�����E�71O3�]������Da�������/�H~�p�.�d�QJ��h�*��<vC����d<��u����h&����X?��ʅ�Q�s~=�e2wN[��B��J�)�f%O���)�|C�2t�m�cp��,>Jp�j�AI���QRb���Q{��k�o�Le6z1�ș���f�]�#������q�T_�g��C�r�O˅Lq��]���Jx�D'��w���?��s�̳��ހy$D	{Zр%��8(�(�S��Z"|��ZHΉ�W��z��E����K���Qz��$���*��8l��xk��;�E�g�2��+�b7��:�����v�S��|❙'�W�u�:pl=�[ʆ�uu�}'�a9�9��h;��e��38 �{�G�?��!x({\)D�@�l�ZP�JA�f	V3����V�=���Ÿ��d��[|�?����U�D#F��I��,�߰!� nw�O�:�T��ȈԆ���D��(��Wق[�K�j�#�!�%����� #N���,�-S�{�6�\��5��,u����?	�ʅ+"o�z�$MZ�A�y�������ʫ����d;*�J,u���������WC����9��$��V���h&iɖ���d��Z�'���%f�>��'/aW����Q���t/K�)&&C�PD��}szz�ш��eh��؂��R ,�KQ�}K}����"~yf]�1��w[�+��*y����L�N�*�b�t>��2�tn��fV�R+�_l�-��,��	���x���=�9ˁc�u�8$�/�-��Z�`�(x䎄n��v�zymޭ����<4G�� .���.IJPFӮDT�a�F��A~���#� ��P��#v�>��ת�����G��Ώ�&�7�Cݏ��۫�R��7��^L�Fr=�'H�Oי�B����~!���ZZ���!'\��v������Ō+��B��ԉ�sg���S6���y�@�X7\Y�/f�&����	E�T��`�]�������*�����r��W6$��<��V�c�vmj�'��ʂ{����D�����Х���S�s�<���}�n��}�sa��Z��]Y���})��xΪN��fv��R�K�N[��aq哭ؚ'�C��n>�?�w��n�>��v��K����!qU�
_�k�"���C�4��K#��)U��C��Р3�o�p�w926i��%?�G�Ԏ?(�)��oL���������kHN��m-���zS��'�ms�C��p�)����E�uA��l:�ɋ��J�'a����CYY$8ŕ��� D:������!!�y��Hfxtϖ`� �D�Eou��G������{b�2R)�h�g.�I�Pζ0�r�6N���o�w4���k�J"H��yv*j�K�j�{�j�ş)�����ue�\�%:+ ��M����ʼ$�)Q;�Q��ۂ�>��-����Cd����=��/Z��˗���46.ϺjE}`o�ײ4��$K��3�K����b������L�l�Mr��;�Q0��g�Sc��Y���3���s&�:�Z�<|�<d1g�9� �b�� &��A�$�o���:Q,Ϭ\��r��˟���P����o��Cnr��k�̐�ZGmS�tXů���ë@7Ӿz�@Ϥ��
��D����)�@Ѵ�T�h2>ZHo�h��C�$y)�6����$������N�f�,���Wggy?���.��t���OU�iq[�����݉�M7�?�K�	�z�-�̈$&�k�j�^��]4�j��&��i�����U$Y����#Q-�R8�OXR�m��4/�7c�u��"�����E���������V�?�y
�P�*gy���(�	޹�g�ܤ���23��]D�B[�,�$�S~ߢG�I��1ꦫ�����B�ୋm�x@�!������,�u��ԉ��� i�Yf���t�}���vJZ��UأݵZ�n�!'�W%�"SпgCy���_/@�M��`���*o($H32�=���2�CEڙv��7�N�J����!9	�'��S��b*�N�_z�(	W �pw���{���+M�ҡ�t��-��n��$���_��ˋ���nA�`׼��nغ�9���q�z&/ׅo(R?=yט�dэ�낉��P3i�7��#|=�+-K�d������W��h�X�ء��#�q����� �0h�*�����u�$�b�������X\���l��E��ٙǋmV7�=�]#��������N	����]�)G��t�oY����Y��|��*xç�M�� �Qb��!eW��)���"Ƕ��`owX���Ow������8�غ��:��Ô�P��dҌ��(�X�%��|�C���:e�R�45a�A��; N����$�MF�4:��S����``�9�3ǻj����ٮ� /wb.WJ*�F�Z�N̘�<�@)�`�_R(R��5XQ&()�L$q07�'+FK\>1/�M�D:!V�������:�$��Ŗv���?�0���)���/����L�W�y�{���z��f��
"���5.���gj��8u�w�f�d��N�X�ݿ2l�q�t�Yz�cE� ��p���@f����@�c�K��is%
1�{���r��gk�J����&�ώ%tx��%X��-Kj�拻9�p��zO�ދOeZ"��(�5��(0j�*��CoO�����+���tg��X�+����r�(�[=�˖R{���fY��3n����Kh_)p��>G�����Z��|L�XX�H[̴���z�e�(�P��w��J
w�R�����|ou�����X�M/}�m{
����S����:ۆk�
.w����Gk��ً�m��?�u�Z�K4�y\�ߛ�������?S��:}�B1J�>��_
Q��ãP�G�|__'���!�ĳ����H�u׵c.sn�.zBss�	������s��*�B���j:����&���Y��צ�q���T�E�������5�@�_~���9&-�#XQ���S5���-��U�\h$�����n�#����^��]Ny�T\(*M�jm��v�C��Y�	��Ƒ�����_�Wpϗ�5j��C�gN-)�$F��hwP�//~�C����`%n%sL�u�V��~~.w��i��wRD��"(�����*O��}���[p_n1\[���c�J�jX����}s��=�����3�<��$��_SQ��D3�z�?N����EhE��ɳ�����ӷ+�GsE����ݍC��O�����֡1HJ[(���c��̈	�We��ϰm�A�yYO�aQ	4%#CW�bq�p�k�l
�>�q�s�V���YFR�C�V���y٧�n?I�=�'e�����BLN��@E�_ SG�fZ���]j1�3�q���&�z�A��O�s��l�oj�����A���T{å����'P�lX�c�N�/c8V��΀���'��B�5
T'R��y�<�h�o2Y����#�&?�L�)n"������:�3iB�������@Te���᳉%�Q��Y����D|�^�B���wW�.�U��gq�i%��N�AG�-$�̆�K:X�����1u0�>O�mf�胋;ssJ��f��7}�3G2ǹ7|'����e������t����$BF�� 5:��ËQ�Q';N�����a�L^��mrbP=V������'\�
J���$6���ЇƲ�.���拷��y��B�\4��w���R�@��:n��m�P��H˄f,(��n��WߡǛH`�����J@�ȍ��̂y��"�G�db���+ޅ덭+�x�<n�?@�^r�B?��6�t�E�_c��2�m��9�٥����5���|5�0�#8���u�?+�H<x��ӽe��ء#Oę�{�D�&v�m�����~��s^��}:Ě`�՘��1Go�N,�ڦ�Ο!�5"���/~ϭ��7��u��g~�g�^�m���:{�B��[O�OL^:6Od7PLū��`RbI:o�E�����������m*Q.�ˋLQ*]����d�a7]#����7Ϯ�����	�V��5�q́v�Z]������̻ϻT�k���2p'Do���/�Q��>{�Ey۲�O
��T�r�����{��h�Ne���3��<��L�ދ��	����O<���1����j����y���
�][�z]�6��ӣ�/�1S� �;ϛ�2�gh���ֲM��<8W��TI�Uu��_!K��͔�0���e�OmG�崠��~���N�s��@��o�	tP��P�!�ª�7���zEX���)H��F{z}4�0�ONP�vv���^�t��G�jb䝜7��!�T�h��gbRB�҇$�
w{0�h�����!�.-��"X�`�G]�{}e"�������X_�z����+y�Z5O� =�d'��Xsw�x�z�3�#0�e��P��N�"�-Xϰw��l=/��V��"*��y~8'��x�W������R{='
��p����:�j���spz�j[�T��~!�x�3�:����w���Ѹk�2���֕��Y������Fx��y�Ѩ�3�8��r� �@�����fd�v%NF"ml��ȟ�,�D���ËB�˱���t��Y�y�AS�)9˵�%���F`ȧiv���)U9�.�#�9�Ѣe�Q�Z\���	Nʜ�떿�w�� �x�P�����_8�<S��)
��w�$�#a
8����r� v��mi��4��3����S�Y<���p�,'�Ϸ�7
۶�#�h	��8譯���v�������������V:|ĝJ�>���6]e>5�:����kR;���sw�m����6��D��e�$B��������[�AIiH/����a��}:s~A�㝤$���<� G�}�JC�h��?~��Z�3y�r?����nY �X/�]��u��i�J�$7z����v� ����K��쬥,��g4)ι��W>�Bt�����J����vo<�]�ٝ"Q��0Q`���B��I)��7�ō�eܭ?�
���=]�}���i�w_� 5a���'!5Z���[�*���L�� "��F���h��-�d�P�BLVޏ��LC���8���AW�K����
_}>�
�03�>�u��r��wۖ�u g�nNU��XJ�������E���h�_N�S4�og݁]C�
�jE�H���&f]-�C�����6�M����I0�+����!r��fV�>�#�!Q���J��y��Z�v؝����hF�`�V��W��v��	����i����w�h��U�'	9�*�.:�sp�N}��܏��	�!��TS�;3�vq�􀎆W:�cw{=I�d9Da?ָj�.� O{K��Y<�4ܾG�=-����T�t4���HgU5}�nsp-�o�H���l�����k���,%SX�y�ǎ=T1�3;�^_�S)Q��$(�c��k}��5�H�]hѯ�1���<(5�������hr�4����'Z1��9��2j��}�p���T[����qa����p�+�v�C
!�H�}�1�B�GY@�����5�+�g�5�/���ˊ��.�<��>���.�/���ቈ��M����L������� #k'�����GϚ�q��ܘ�X'��≸����� ���_{�5�g�8���o��z2yKU�܈A���z�@+�y�N0�MpS��I����ēm!S���\���qqYUH y�|����ִ4dcas�U�I���k��?Jd���=�)�$g?=�l�{��A$r�䋭O�ߔƣ��R�^`�����"oG�/��3�W�,����T��c��\ƢV\	�֯j/w�c������٪ƣ�e�T��"����X��^�(}���T�i���m�=U���9��Z�%�:}5�J$���CG�j�TA�J����4�����1���h.�}]�?�2�n��2y[��a�9�R`
��* �0C�,�����|ę��D�)?�I�a9���\������Ԫ[2d��&�W�Q����UmC�G�^�`���W�l���.t�`��������u�Kk	
-��_^4��L�S��)�����.jS��nS��<�Ա�����b&|����{�6`Ou�hB����_������?2�L��#(8�{Փ3"�Y�ˈ�ط��k1���Y�OL�O�}ܳ��|}�2r1ф�)��^�/[͙�c�Y=�6s4 i�J��V�ow�䧚�rpR����<^�D����&���ff�D"�@�J~S�?��e)?]H�������ePf������vj�Doˏߤ(��-�Jm�������^m_J
(�NG�0��y�@{�L]�i簱=u��F�K�\���{mI���nNk�-3v��N���뵎�N/o�uv����+C�&đ�~��6��)G&u��3���G�s���(>h��M������3����{I-:I�hԔ�ȹ��sbM��L4!���_��;ݵo�E �6�5��y��L<I�E��U���m�)�rl���Z�&Ȳ�E��R�X@�|�ܮ�՜�	�����_'z�bB��zX����'�5� w+����T�H��h��G�����a�~x�Z2%��AX�FE��?4��c�m_��F�WG�Iߞ@��لqQN�TI�2=��-j�A#�t�z,���
]���\"�ܔ���X��k���-���(�5g������CUu�]��2�<�/$����I\�f^m��Ԃ��X�lb�a���+���ϵ"�H+����;Ur��u�\��SA���/�*��*?(�8��-vN�ڗZk��0��{7p"A�ɶ�sƑ�u�������\���Q�aB�\�6��G�'���V���k���AQ����W>Qv�+*I~R�96��6����eJ�FLh�(k�G������h���/���~2�?���A_���w�ϩ-��Ɉ������I�S_�2�Z��N��X��e��"�����(4�Q-��1���X���BFX������i��i#L2�cI
1���uS��Ӆ`�� B�B�`F��`���&A��{t���(�ZT��pg��u����q>��$���8-�!��Q�8��yT:�[�k������,U��Ěa<ej�#���c�rN�~������n�u�l���6�g��e[!1��{,hF�X�ܤY����xz�:?���{�&k�k�WSb�o���C�v�Q_$R�#��h/E��ؚ�Ě��|u~�M���2��hw�fg4�P1�R�Sx�/~��c��ئ6:h�]%��W���������bIqA�bH��������ũ� ����}L�}L2rh0�%xQ&|�|��_���9ê��Q�-�Mޠ\� sp�J]����)d�U2�Q�\Q���!��]I,y�ݘk�_���Ώ=�;�~ӻ�|^�@�A���=�Ew9���;[���mN�]�%s7�G���n�W�)�֕��CH{��\gZ�LY����~�.��~�M�=x)J�(�9q�¨��������9�ssfCE�̷����}���\陁-/bH�ۺi��U��!x��C���0Z�S6\@D�#����%���_��m��뇦�/��ʼn:��A�T�Wh5[�?�:��k[9�}n�]�H��F�rt�Ro	$���H���5^�3+U|E�^��8�ܜ&�������:��X��vl�\+��x�� ��8�۳#��l��ߞˀZА�����S��XE	m��g5�F����@)�JLx�E�Us�*���*��(M���7D�;��|b����&�_�tM������&���}Z1�OR�(�Ô�m�E�2o�_��A%V�����VW�\�Ey��1z�{Y�J>�sd�,%���"oX~�<�vtM�?��zU�Y���*S���do�� B��e�����^��LW+�<3U��m���lD��g��4�9���?N�'k�TX����K�O?�U~NX��¯�rv�����(��ڽ<Œ�;�tO���g�*ľZ1b�\��eu
����Zy(��E*�uM梐s�����WL��+�������K/�qD�΅>	�:��~d��CNL�Xe��Mf�<S�p���3���_� �yB�W��0(�m�P��_�>���g�C�66�@ȇ?%vb���xL��snOZ���{^�.H�6daޚ�t�f*@�l��Y��<^��]����mC�P�%��}`�z���}W�ͅ��l�y�
��N��l}}��M�Q� �L��b�
��Z�;����PD|rp~�c-/^Y��g3�T��08(/�5��мN��_�K��8�6��Z2���x<��oઇ:�Exk����Y����3_�Dq�d��vB}�_{�@�m >�m�h8�	�/���5"��n<!����󚏙�a��l���z	n����6Y)���C�+�kqѤؕ8��{�;�b;�|~l�1BK��@�3a~����AU*�(����-����Uw�n\�C_Ѭ��y�Ez	YM�MF���k/��!T��>�f�߱`�Ƿ$�O9I��G����a'-FZ��;��<�]�$��M���
����xU����$�p�1mk���W4��$��]��B1�?0���J8W�J�a(>˟�j{e_�n�� x����g��a�0y��4�����~�F�d��[�6�Vn���?�Uh��߮�I�e��1n+R��v"�����"}=1�f����B[�.?i`;��x�:Ē���~��oXd�Q���e��G���C/��� ��a�s"��|�wX:\�}�ϧw�%��������oY&[�<�h
�j��	@ZT��x�|iY���:�M�jn�[�)sF���	�]� �5����ׯ�Y��ź�%���O�4��\=g�h"�Z��6��__�:kΰ1V�������p�N�J�+��d�F+9�O>�yUq��(�ǃ�P��{��B�:[�0�Q����ʥ�A
Hߟe���iEY���pl��r�����3���[��9E?�$i�ZL��{��PN1�,b�8>��2���d��𑿿�&�/"'��D���_����$~�>�T��r��.w[��u �?L_ł�J&#�k��@(���*p��	�+鿔�,ko5��븮܆�)I3�U����e�U�}sNY��'D�W��2a��͜��|N�F��N�v�z-�e2?g8�3�$��f/ě�_�b��!B03�u8?_xM��S�����v߭Q(�������E���s��"5��e��%�0ba�3CfRѺ�U8�:*bP��׭��,���9.���q���zh��0:���(Wˡ�Ӽ�Z��/��ltL�<n���q��qp��H
���tY����N�ad`��;2����E���Y������o��,}R��x�����]�^�p�l1��� �*��J
�z�p1hC���Ig����i$���_�ʓ~�J��M��\�x�F(���s{�S��i�O��Zt����FQߋ��-N�� �QU+42`Rٶ]/�BU�j(l�[�)�i�4�ZHk96H�jz9:L���� آOf�F���[�󢴞��IƑ��97�6VY�.j��O~>�1�Y����+ k	�1�N7p|���dBψa���k�jQq�M�O�U�\�>�mSTb���b&�g`����B���6/!�Ni%�S3�8̹i�L�D��|ԅ�����e��)�o��;��f�Y���C�U�Ѐ��͠�7�J[�_�<�^�6k�����:u��P��3%�x�� a��k|A�b�$b�\�?kp	5��bO��Qk�}��M��a�U�k��}U�Yk����=�|;�E�nL����54��R#���ՙ��i�>X?�S۴{}R:Mm���P�ˣt��䘤(�[9_�?i�"��/B����4����T�7����2h1��Zở����aI|^�72u�ԥ6N6�+�=Sv�o{���N<ҝ/��=1}��Qۼ~`��-���=���9���ޓ=�1��3�J[�z:�*�O
"$��Bog�B��!D�����;]�7=.ߖ� �c��<���X�vyOx��d�*���U��	+/q
G=��w>�!c��Jr�R�����&�.�t�ٮ�7/��׽	V5���Bw�oW�H�P���1L���	�5K�5u1.O������@z�����M�м�?8�@�o��m�fg���s0"4x|����RǱ��E5������@�0L��/�/���-8m�(hњ�%s ��0=a�;I[��.M�SWF����V�L���楩���h	?[T���1��v�e�0�;m�8ryq��o��G����W�w��ێa�k�u�`��t�����?��D�矧I<\2�����{����T.��	]��7�>�=;{���YXW�sh@��-�g� ��g޽H�3ݭx)��[�����4L�:[|���t�.�N��գF$z4&*➣� ���F�
��]c��\G'Y�,����4�i�m)�t��o|.&�������	��x)ɳ�H�m���M$
6��#?�`~m ���#g��,�wK�ר�l��ct@j�P6�"��U%�w��*BC#"2�(��ͱ1�.��9���f�`���-���9���;!{B����t�ڑ�Ӯ6���hض	;�J��ۦ�n��u�7�	Goy�]y��uG`��k�i�̶#��Z���|z�8̝�b�rG��>��&VJ�>	�4����u�*! 8u�'����z"۶�V�&�X���Nz��yWӕVn��حH��v���+@75��)UKN�Q��S� �6[��u%�����rn:�+!:эS���_�;�-pWd5�=�.oM�`:��*b��;�ٲ��S��J���)l�w�&�>)�bT �E��v��s���A8o@�� �����ڶ�t����IId�+q�N�P��@o������i���$Q��avDZ5a&#��vz.0�I��ؙ/���Wӗ�M[�uJqm|]8�c��������]ϧGf�	��6S��	)��t�aN���)��P���k�����D�����4�䋘��l��Q���b`\����`g�11�6v�]�;�COoU[uIF2�W|�s��?�F���[WC�r�
�W^i����Y�,J������^i�	};�������E7�QL��}��y����w��lSא��v@&8�H�B3���-�HqC��۞P��&Q��G���Wa��&c��؈}��uRP�D���b+��}w��o���^�xW!G4o˫^�ׄ��_� �E�_&��{x�1y����-�-�Z`�LW�%��T�/�\�L�!n�4M�m9:_ı6Ø�c�/}$:�S����{pI�`!׉
��	���\�QH5�C�-��������a�x=`N6���:I{�P����W&�|"�_-���8W70V���Z�I ����g�!�~��9UX�:�+RV��ğ:f_�W,U�H�Иh�,��5�zչ��4�q����9�{�5���]0��|���Z/Zރ�!-��b���2T��~֌3���J�I)l�3e=�S��>m\�� ��Ư��ZS5S��� �7��4i�EG��	u��h�P\�2�����z���	�w�Y�{fZ���"-��Ü��5�^f�Z�
>1*�Hr�_�;�Y�/���#l��[s����0NU�]%y��q�u�~z�m���{)�%�B*���®��'�f���Q%�=����M�$�k.,���䁕���(���(��$�,��h�V�!|:�-\D���璟cb{ϥ�xK3�k��[E��b����<ǖ������v��V1j�z�h�Yl���`{c�}߀�B�O��̦ک>]?�F����f�M����&��ƀ�$8|����8�r&K��C��j����,J���btI�/lHp�<B��s �K���q�<wg��n���u�=j.!�r�MF�t�zĩ�[������՛��ӌ�򯆗���Η6켤��Z5�{�����8��[Fgk#���)L�����>�N��e`�k9���)�J�lX�����J=\�>+��2�-�8����F���>�E_Y��6A3�~��(����I��,�0������$���X��#��u�ˁL�'�9�\hW�)b���`�L�z!`�ϴ��j�ۥ�/�[R�$/1�a�;z��qR��b^�·�Wr��=2���w�w ��ZOV�V��,[���d�ɂ�y��J�7N0�7f��[.8�c�z�k��' ].�,��=�]�M+b�[�*�Rʅ�` ���a(u�Ge�*-D�mL7�]�������M+��H���|�����آ^�����s*})�K��[y��1#���U�ZMd꫶��2��(Nk��`�p�]O�%�� !����βR�%Y�kD���	�"DYǠ����+t�S��nͨ�8'��y�r���;����
4䴁4G���#�_�,�� ��,�Z���}V|�e��l��1�q���"��I8#���զ����~�ū\��2F�N1� 1�MN/mm!�;u���]Hu'��Dl��n���ƴ+A�kM����*_l��Լ��+�BM����M��K�T&䈘�B���u�ڍ���tK��|�MkSw�����5���!��TF轺��C���#[g[9�����ߪ�����/��3��0GoK���S@�����8�5E��nKH�jD�?�/B�S�Y~�N��}7$���qy��tI��50�X�Q�_��Ij��BN Dk�P��E!]ѧm9?�X���=R5�0\���~Ks<8��8�~�:���ٍ�w#~g���/7��1ݝS�����y����x;1�Z���b�,��Y��Ԥ�}����4kjk�u�^f�Dص_;�Y�����|�;�'�E82�u>�`A�>�PT��|�����i$[zr$Qj�M�ܾ������GiI����z�}�8ybx�Ǎ!���:�W���vS�D���qɥ0��2u*I=�}]��g�E�ab(V��㽍� ��e���C �񷊯;�0���u���߄��EU}<\���]wƪ�A�]F���}�i�|����4���o�jeq��ׯ�&I��bu��i������v��r��MG��V���7R=!�me��~%�/��m�P��g]���o�[۰�C��,�df�l���g���q��W�q3�h:b/6�/�f�~�K��n�0��N�$s__ U2ɣPS|>Gi��^�:�%;//Y�|�Bj����bJ�
�m�A�$@kE���}GB��>�dAqM�<�]�ְ��F^ 04�0؈�B��������Q�T����h��\�8�������v����ֿ����\ܺr,�S��ru��	9/U�m�ŭ� 8�a�'�jaNb����f`���f'�z4{G�y�c!f3R�~פ�/�W]~��\�Bb�
���$İ���|R���H�v��k}>/�Z�k�1�;�+m��x�/� �sekd��Ԏ7���z��EO�VD��f>p�gl��
R�G~��A���7��Z_�j�D/+n�ﴪa����m�(\(byJ�z��ڸ]&V�0��<�p�~YCB��:��S�8��T�������~�^���*ة��ԣ:K���_�#Fx����G�_�79~_���l_Y�L����u���:/��dwM�#���LJ�}$}�'%�~���%L�zK���g���E�=�'�v����)J��A_\7D�,��%΄F�r�޽�%TNq�!�4��@-Dr���2�����;��T����e;V�?=��v����Xn�'������7�M��oW'V!߽��LL��}���j�	��������墹٠"��;㽫���v��H2���Ǐ�6����yo߰kW:o����1�%F�	f#�8s���;x���;K����M�n�ۄ�8���S2�:�b\�:��d��TA5�OQ)���`�v��>����BT���t&:��F�O>�v.�H� 4Ԥ�4J�%kܿ곦�����o`Ax�5��l��H��������T�)���n��b���{/�i7�,.�?�;q :�b�LE�YMŶ�h:��)nR�TC�ٔG8יּ�6��5��f�o��&-?�lb<��'.?�^pe�wρ�`2ή"�I���k���~f� -�ǔ̻��*�Y��}j�_�=�1���O�Vjy�r�M�%��Y�]��B󹨾��Q�������M�a�R9���bS���¼՝2]�i��q�8���}��������\�|���M��<9H٪��#����Tq%$��W�qzH��}{ǈ����Hl{�������S�i���Ң�򥰵�
�#^��0�״�t��YH�Vh�Swgٯ�$�����{�lV�9� UA�h�t�/t���OF�e�Ѕ��
y�Qwޛ1�^��W>�h4�U��ʺ��8���y0t|vmO�G��R:��\#�"�t`־da��"�F'��|�J���_ki���S���e���r���c����:x��I@�3�����<R�Y_=��
��%�/�T����{�b��t5s�����k��Z�Ό���[f�~W3�����-rZ��F�S9Tc�~��Wʦ����uX߿	:��p�Җ�O�VuG��n�[�'��M�Մ�{T��* is��Cfs��T�Px�߮8����*���-�N�����܂Kp���wwIpwww����n��y����*���e�o��sz�e�����)PW�؂]f4H�\~�l� �_��ʅ=y�0MFܯS��׺^�8��8�NW�@�^�r��>�O���5���ɢA���� f���m3�w�E���t��َ;�2�����X4hƴo{��a��G�^N���*>.��UW�[}f��"��m�XoA���-��#R��qa�t&�i��d_7 ��g��Mp�g��S��+�@��4��(.�����9��}LaL;�s�+��	O+�dʯ]k����
��<��_U��e�ﾚ9�g,ԥl��t�����N����"G+��bS��q<Qn��l����"�_QZ�4�����aO�㧢t5����w��V�B�bī��z�0a�d b�{p��3b.����-��?�3oC�(��qThNa�/������u:�p�`A�A���*/�V���R�g�כ��v;�zSz���i�a��H��ˉ`Y5�&�q���N�+J2V�����4�e�X���n:PZU/3x�$�`�UV���L	�f��,����A�uZ��*+ $�^�j���M}Sp*��eA��48��N�r[�I�J�Baΰ/R�T"��_$�[�A|�}ŌB�l��%��~�u�KoǾfQ�����0{�ў4�\�K*1ڂsn�XT��hע=���+�&��,iM�Cn�����",�a
'�n=Ӿ��i3�%I̪S����R~A�P�$<�܋)0
d�O���"p,������$�#��r
�N�X=f��WA�f����5��<�I$Cx �%��ۉ��۲C?��'����`�f^^���^צ�����u^QF�7Bt�R7ƔޱE[�S>�SM�s�Hh���8
�n0{�z ����\m� �=�
6,O�S��ߞ�,2$&_״��nT�tFܓv��ʵ���	R��S�q����Oab��.D��K�s�u�T���W{�c�M�J����4�`W��z����P���+��!~h~X�͍˲���Nd���:��F,�ӑ�z�u}�+�[Uը˛?.1���,D�]��vB��\��mM/K����#�5�����V{��Ew�����݀���j��wȼx���M7�x8�u�5��c,MOku�^��-�g[#����NᏎդ���s�.�H&z���1A��ð�_����d�1R|�xٍ#�ʗ�s�e��5�U�J|��($<��_>���_*/�����s�F?�c �S]�C4��1��ݰ�m���T]��IK�����1���	u�c=5�I�t7]ؔ=Բ�$��0�o��DF�˶>�̘�X�16z���!S2'��.��ۑj�阷ؾ�s/���Ǧ��R��9��D?O�n��5�L�o�ٿq�7�u�qhH�,'m�u��e\P@L>!2�Z�n�!$s}��05	��|��}��)%;��>�C�Q�՞�콩6��t�{��m	_k+p��h�uIa9�J�ۙo���/�.�3o��E����v[JC��B���5hN�Y$�}��U�*=�.�����Z�h��ߎ,�X}!#�rAZG�����D��:����+,��k'��Շ�W(�J�{Kp���$>zW�ɰY��~���F1�d�Sbɲ�WZ�OW��74�Y$rnv�7�Sa hH����`��+��#���n_���i��+F�(4���)���Tvs�~ ��x<-�� �I�*��!�_�m,!KlGxG|җa���g$
���oc	~pW������/@�<��ag�5�W�I�����`W�vńx̝_6`��ZLk]��/(�r�?4YZ A��i��w�hT7=/�/��K���X��i8�� ��j,��xn6���P:
3�2\�����{�Hgp��������:���(��w��o����%���՟JY6_n��>N3�<����/{un��ҏ�H�k�h�7Q�3����+�cB�!�.U�vdmLy{>5��R�Syi4V��U$-��e��C�i�=�9��>��
,�'�&����,((�5|�)����G Q�pk�&����tu8O����ӏ��{�7t�po��`��#�+�����y?�K �#O��B^���(��k��D�
E�3{���������rxgu���(\x"4\C�G!U�����������服4Sp!�t"���-�_\���OKE�h����7U�'g�~
��Xp߼�Z�|����qS�O4 F�� _|�B�^~O��f����K,{�B{3��Vc]x��Vk��1F}ɮ��2t a�9j�P�>B�u�t|cK&�:d�P�Q ������Od���K1����6�o&K��4PGW-M8ve�S�Aڟ{����?|�3|c���{�y��8X��d,��V�k������y�P��]�@��f��*�NJ}G^��&�!��X�����3��������i�g[����|��J�7�}���j�ʪ����:�����ե��=A@��}��l���l�	P��0T�kZ��G/S-�	6o�A]L����R�O��M��ɣb����*Q�D�*b{⍖�3BȾ;��?�����(S�r�V
���G��:(aer	&l�1�=�2��}�m\ֹ7�Gn ���< �D{e���	�%knv"��{~@�-Z�h����f�1\������0�~���h�������u�f_��C��$)��r�K}��^d���")�4���b��vK�/��*<Ek;��B�v�K%�P�Y8�xx�6u����P�����(��w�LV�h��3�}5���j���>��vJ@�ʥc6ڥ��23�@�",�*�t��1"r-�A,����8,{��n�rY}z}�O
x<@�����$%h=�]�C .)z+������K(k��,C�J�����������x%<ow0�׸��p�yک�e���9یb�����(Xr�\��G�Э������}�16�;����w�!�Rz�Ej�& V�Ԙ[%T�M�i��L��Zp�\���cP��a-4��K�ct�,����С�����+X��9L��:���a��oO9�/:��:[����dNQ�6uWL��_����.���n�h̀�þ��뿲6�"�JFoHL��߽J�A�X>W��U��^ze�z����u\���(�	˰�����jAB�~�p��B	����M9�-�v6��8 >�������O�����:n�7��\���/O��/'{Od����$#��֋����ݧ]4Z�U��-��J˭�ޞ��5��>k9)׎�ۄ���w4�Ӷ'� �;�I�ڑmv�ġQ�u��A9���W{�i�����S~6�i8������>�[�U�~K�����.w/1�c^�(RS,�� � 8I�"�*m��K9�L͹�]o
Rvf��T�b\" ��Utܞ"����S��mƩK���K���2��lQr��o ���}Q��g�}��������iw�,I�8�on7��f��z�-s!��B�X���(�:r�U��Ĝ���|6o�N��W9�^�,�l;bp���o�7�RűHC��׿
<�>G6���YV�DXPO��u%�L���H��VԵ�n�� ��Uת�Y�0��˪v�ٙM�V�cZ��!Jr>7�kevБV�E��-iI�u��h���wfr�,w<8�ʆ�
B�S�n;�����ȧ�]��'�Y�V߅�g%1q����	ݍģ�S'���Q��z�L�H�}">��㛆]�.�Dv���� p����/��ĵk�^xG��bn�l��q4��0��n*� �̦���1�\~��ʧh�0�J�
f���:<EA\U�W�����XT����~�Ϊ8��Ȟ�@��8��1��m��6&"��ޭ���Y�V��;�i�ai�]tQ�T(���Y?���g�����PIU���y�?��n�d��W5��� �e+�,o+��a/�.��k��H��kS՞�A>:DR�YFm����SR����X@�C���!A0���VrD<�w6�mF%W�͢�a��ݵX4m������NM���&HƑ�j2�%�%�-�¼����0�V�ݔ�,�/J���;��M�'�D��?�r+�D@��X�OÄ$�|,ĝ#-oƥvz{yԴ��S�,k��ۮD�����M,�Vm����<�i�����l��b�=��Ԁ-<Ti�˄��aC]'}.�z%J��t,Z_]�����	=���5J\��Z�@i�by^���ۙ^H��1��  ֖�z��Q��9�ҵ���+b��r��ʍ����ȔQ �����b~�s0�jz7T3-� ���O���]�����{�o/U�������4�t�P�{�~�ܸb�Α��P;L��5й�}��,�Ȗ���X��q��s�=Z��e����M!8��3)���D ����/�쌞��_��%�L/5ߺ�)�,���?Z�^����-�2(q�y�2��
�~C�.4A�p�u8��S�`Z)caaI���.<%E���%��k2��k�PMz�G����r����
kY!��1�Ǻ[.'�b�y�e@�[W�7Y���?���W!7_P��^��_�?PJ�������y��ܑ��u�ծ���΄�DB���+�F�z����5����|L<���,:a���X�z���� !,�qI[ʒ%u���~}��X�,��p:�X[w�N	��4Jv��8Ek?c�R�x����*w��p���w�
ұ�rx�r�D���5�98�\�p�?���N��w����� �D�����!G��S}�5�1��w�-�H�J�!Qu1ǄY�W�2�)�C���w�n��y�4K�C���?�����غj�C}H�*����Ł�j��C��ތ��\�����A1�/l�%����K3�x�KǸ{|��v w�F�(�Х��r�s�A8����.���&��3���W�j@��od���Fk?X��NM��`3mN���Ui3�%f������o+Bd�4X�'�-Ւ�$���-���KV�F��4X$a�؉Q������O@��W��eelŵ	.��%��Sx:�ܥ��b��Ѫ��o�dG��M�]5�"u���-g}������Z��� ���n���}5R�������fW��<Z����9�{:ln�Ii��%�،ަ�E�[[�L�W��zj׬��6���zF����++B�$u�&�����o�=��W�k :<!�S�D3�O�����ῴ�.�Mk�n�?����+9��7C���,wl���uش����\��I�o��u
�����k���j���f��Dl483P�gs��t{����H��.����,�͗Z��� �A�~{T��'4YG;eա)~��{^@���c�:��  �%%*�"����ȗ3�!Շ&��x�w��S�ʭ�����c��5�v���^�}����7&�pofZ�ZչL64!Loh?�e��h����|�}���%
6�C�$��g�����W��^�c�J"���~�L_���2��G��#�f�tm*v������fA^:	������G��������렜�Ȼk�B =��P�g���6qo��SS��ݻ[���������B��e��۽~�?�5oQ�U�� "����?@3�Da��1Q�ׂ{�P��E����'�aGDP����E�]�꠆*�82l̓�7>1ɀ��7�o�	p �4��*�-�7��@�����p�_��(����E��Q:Y2�;����Rj� ��Р��)y�����������y����>k!*]p�ipS��f[	�7� �L����C�c_�m��!�y�!�Q�Ԋ���j��E�/P��´>��B7%4
WQ~�6rR�վW/��?Ŷ�Px(+;���z�����bO]�X��y���ܦ�Z��[�h��A��/c)��""߂�23�ld`��o��ǳ�Em)w�=q�ͻ��bQ�D٪���9*�P��v��U&`��D��������`��dE���TC���3jcn��'��<� �3
U!�G����9�
��w��ۤ��x7_���W�t�6�UH2�5o�O�$X��{K��S^��u� 0����v�h_?���s����N�}S"��^�Gh���V��͟�hqaS2����sA�����b+@��s��� �99��$�XI~��O��iQ���(�05}L]g5b(7=;�o�O���d�����+�@�q&�����T�w%J8	�/�(DW���Z��i�?�E�C*|߶����Ѫ�>�s�?�dԣ�}���<�E'w��lf�\�74��Tv��X #�����-
�FJ
t}IlTD(�,��(X��R	 �%�27J(Q��1�ÃE#G8��Z����ϋ��ae.x)<���]�T�Ct�6D�v�0.<yu0�h8�We������g�Nr��e���9ӆ�I8��M\�/O����L�I�~�E-�_˖���$]�g`�Gc]�=��ɥ�>�w�^@{�oP�é���)�����y}5�� ��PFR�ܦ�})�>'���@�C�$B��(P�I-fė
�O\�Y��Lq�3���L[k�r��.��*�T�-(H�q�<����9%�9kl�:��i����Sk�l��Q8�j�A���}�0A"��3�>�߼�ZRl�$sI��Nks�@)���� ?���a\��S �ԯ#��|�n�>��+u����㓠�4���(�y��������c��HC�gt'K���pS���3!�{�v�CY���ۆ�~z��լ�<I�x��"Yu%��Q����N�8�����Q�W�h�O09l�ٹ�OO�5�˄�%�y��ao_.4�6G�Oe���4��B 5�w��
��[�pl�p̙���1}P��r���	��%�!�~��pj��ϟ[��B}9�u���YW��a���@Ј��ý��ե�4(&Yôש�Ii1A�:�j}*ڳ�؄��а!�ȏ��B��c��ȥn��"�s�H-o��Z�!)���'��u�*a*�Z\lml�Ǽ��{��A��n����P]��/#�a���a��^�Lt �lmaDe��X|�(Q����k�����1?�"���
f�ڄw�6��ގ���y�p��n�M�6ʸ㉇���Z;DT�3���&������S���կ�t�K;���68�d�{���u��8�zWM�#��Es^k��?C8��zE/������~D�0��	�˫��[��oC�<c=�6Hv�3q�4x�� cM!��Ms���}��3z����m�ӄ�$9�U����[��Ԕ�8�6�|N�T��
�k8�u1��yI���fWԍ[L���>���L��������1�+�Ә��Ƌ@%t���fo��[�Y�8�!}F�پ����M})8�� �<�4������,(�{r)~�I�4��N4&�Bc����T��oc\9���%(���\�.ܤ�:BaG��qE�}H�K���p�-R��GZ �~@ Q��A�����t�BG��{Zc�>�@F'�3v�g�)��;AO<�:�2m�>�L�me�z�v.�*�sg ʠ�����Џ�/�������7W�f���ճ|��+]]��	�r��}�''���Ya��������2lfW����ۗ�`f�tPT��gI�ʅ;�*���ޏ���*Ƽao߰_��]�XD(t�f: �Ј�2wi
��z�n1j��6�%Ro��V�����{�4��:ݎ�>sy���F%�j����~ �x�\��$�܃⪙�������ݽ�r�&�C�W�(�ٙ�P��Z�t��k�ʢ�;�z�␵�j9�l��4�1�����*b*����8�$5��K���i�U*�����*:p��j��8
���X��ϙ(���E/R����K����_��V�Ϸ�N�!!W7��& ���kM�� ��@�×�4�8!�` ��A�\� ��UYV�o�Ց?��Pu�e"-:�����;}������������,)����0��@��I����߯w�E��>�M&Cx������˼�w�+��b�Q`@k�3�vs��9oME��U#,�V�[?��K�m����]�c}OK�'��&����o+SE����ngQ�S���W����l@5F�Q�}��|�7�03� � ��P��q�rYMM�S�}T���*�!�����^��p���s�g�n9fDʖ*���Y;������Uߙk����oh/f6����^~	(!������[�
���%�̜�����!��
��L�	'�C�@�����m�#:�:.)A���#e)^n+���ឈI�<9w߮�Pl�֛��%Ψ�j��5>|���ӈ��&�g� ���~�+�x�������:	7�s��:=^�wv��P8�b�9�" ��#^Gh-��p�T�O�m��=VI}7|y\�N�����T[�cƁC��g�AP1Tϸ7��q~�d�ҽ�<�~}kP.(a�[c�AY�����~ī���"�׭ٺ��L@���li�٧\���b�� �	�#rr���?K���U��iz��ռ�lr�M�u��ֺ���3I:�dBf���YW�߲�����G�H��*lfߦ��#���R�P}��Җɋ%5z��F��{��H�������Cy����ʓ�7"(�Yfg~#4��dg�wrs�+����(Yw~�Wwy�]^A��;*�>���L**��F���!]7gi_��b�۞��:�b.^u��'Do�m\8�l�5�5�g�$C�Vm/�n=����N�!�h���my�_+��O̹zx�smؔ��P� ��1,����_���2���cg������Ĝ0J�B<� %�k���WH�?� ��ic��]F&	�ѣx�3���;�������!���Y0 Ø��꼵w��Q��2!�ֳ�ͦ�DޠOuX�K�����1��fFo�dP@s�:����*�:<�ns� /9a�2{����;%�h����2_H����'^G�?��t<٭�=۪�W:�J�^I8�k6�������l�nԴB#���=�(��j�(�?�*���Z�\�ޥK�T���q��������֬�����~�}��Z,��ֵ� ��i��>�aUu��/��������ܪ�E���{�Ic4�rFag`�{�!>n�����F �K�a?R��X���+c�?�z�U�<)ь�X^��o��1�]D&���6���@2kpQ-�(�\H�x㚐�n�q����x[vI����EثO�G���k��a��x�?������Gk ��ߍ�Awg�3�;�����F�Nr�w_q�e���Ѥ��ҁX'%0�S����r8)��#[��`���OlD�I���r^5��;f�E4�N؎ؑ"����G$�#��䟭:Du�u#rNc�L�!��Ws��k8�V׃v4e�8�!)B���]q�����U�GA�k`����h���q�,�"�}G�7	b���yI����3(I��@��G&��{OW�?Sצ��ͺw�GUh��l�N���B�@A���� ��������ƚd'o%сO��.������͞�p�H��R���D���_~��wn��C᧢9�C�?��������,�=��\�9o dڣ4]p���/P��b(d���$���d<�K�̊{�8�͗	�ZJ���7�_g�\T؝*I�J����|C��=�h������,e':�v��+#�^��&��P	P�=Z���[������Jt����~-�	xyLl��k�\�M��@'o+�����!駼e������*xҖ>���t�����Bϯ��T�v2�������՟n�u�Y�� �wa��z�(,-�x�M�0�	��gϷ�R�_ ʕ�i5����;v�H*}��n�P�m�]����%t!A�o+��E�P7��	��20�1<��>j�A�Ф�5R�Sz�S�/֭RViu����')%��c�3Y��]^q��̖��y����vќ0�{��BDTT'�HT�K�\��'��"��6G��a�Gx��mW);����rJ�>�R[���J�5��[u_G[��
�4D}���E��C�I)n{�c�|��>�F�y������e�	�sČ4�3.ź�5]r��:W�������{��\����<OHoҩ�[2蘑��g��D׆��r&�󳑈ij�{r�]�T���𰰰��~�����
����զc��┖���pӊ����y�[H�L_ĘB�M%�s�d��*��˲���n�iK��x~J@ԸZ��W��Ld�p^�&��c"��'���4!�-��-�jn_���@2���N�q��	Y�M��W�<&Q��CV�jo/N�2�xG�g�֭�$Z�6��2��uȥi!���,jU �4O�����J�}��x�$�W��M4Vns�"��b&� ?���]�l� ba.����L)�%�x8�v�L#�J�*�t �ʗov�2�� ����7O%��s��-�~l�!tG�U.�s�l���.��:	���Rַ�;���͕��K�V�����El��Ɂ�#�Ja�9q�����>�bP��<Es�S��j�o��l��vk�K���.������7+*��e-�vW���:M�{��G ����̖S��XӨ#�A�"��Z�����f���S��v����a".���pnK	
r�"�j�K�\ַ�<��s�y�� r޻G�J����/o$D����0�T��5��aa<�/���c���Ф���aլxi���W���^Е�{OB{J�g��6���04�ik�v+U�N��Ḇ�p��W�&���j_I��uPm�é��[(��������)Y�8�'�zn��7��F�sf�Jc�=V����s��b׻�G�V��:�(���%�>b#2�����	��_����	��P|j��ӏW��Gh�+�M#��;1ߚ��t�Li6�?8u���Z����8�?]�T�&���[��T������ݛ�j!����:vD���R�G�%��A�3�c�U��4<3�w�a���U]ξā�P+�f����N.��WaaD҅�!b�n�Mt#��}�zf�U=?tO�2+z3ꤵyJT������y{�瞢5����|a�ڇ�_�"Gm4����Ҽfg�}x�����P��uY���(p��C�ӧ���\�{.�O���ĚuR��{�#�[�ߊ�+�����X\�N��z�̰�y�<?���8<x&�F]r�F�c�n�8��-��FeB��l�e�[�6m�p�-�d@93�;/	f|�,!	��њl�p��+���������N#^�!��c��+��Y/���y}����p�a-I18�	UuS���搪�r��y��8Qlo�����XעS�N.�7�8���x���W�������J�z�!Ή�!���Ls��Z�mM�ܽ��S�|;M:�m��vՋg��˕�8ShDϣ��U5k/,BV�E��(ߤ��"�����Ǥ��u�(9��%�!�ے�Z�,VӴC�y'Ċ���Տ���	��'ڑ"z��l��y�Bxܢ����;ÐK��ں��`��V��`K`�[]-ЉK*P+��
��6 �؊
�z]w��	֓r<]��ڌ��+���/��\��p��3uC0�>t�X�x$�)X(���M��v�� 1x|Rm�o��#xf%��md5�?Ѓ�2L�+f��nU)te	s�6L/Hq���c�!r%V��/t#��o-%(��C�(��}-��|�#DŅ�ח2b�r�B��F�;Gzs�_�\P&R X�I>t��	C0��[^;R7.$�[£kO���<I�U"����BR�M���*?�����zY���N������Q�"v����mD]fw	�M�I�	��{R���	#�U��v�$N�̤ ��_؍���	5^r�xemVrq��������.��@�TM�Zi��6<��*����k�;��}^xg#\���H�RjT���s(�-�AV���.��Z?�˚mD#��#9ccB�!�w��P;�^7�p#϶�Žnv��!��:�Sp�ߟJ��H��~�ȅ&�ll��Ź�Ь�����dU1q�%>w"��{���}7E'��	�2h��=B[��^ ��n�ݿԹ��uܿ��.1�g*MC[��
%�+��'�XA]�v�}�d��ͪ��R���x��P�0랛 RhWcƌg�>�C�l:E��R����o2:3X��Ƚ���076��.Ug�hB>�f>�a������;Y�����ƌ/=�b�Uh�>�*A^�D�W��G��u������2���uZ�(X�� �J��z���抍%�Fe~��<3��l�!��+��6Z�k�=T�Fگ:��7���+:��@Xsū*&�`���ͪ�!���oYM��蟖l�3C�Q\�3���x�� �hG�MeK��dK#�J��ĩKZ��=�@D��Y�fG�p[�&����m�w�ZJ4�g���ZnV^���H*V���FfÝ\
V�*I�*1��9���+[����݊�ӯ��!�f(鉒#7-��+?)����Ii@k���a����u&�q,$`��<�Ҭ�U �a%	1ɩ�����j�'� m��*ɪ�:F�+*Ħ���3��Q*�kI�KY�E�
Κ�;�ٔ��~��Vݎ��l�w>,oB��N��2Q]>��]��غʮ�~zӄ/;�ȋ�����u �αb �[A��6H�eAk:Qg��5�&��,&�WS��4m�z����[}9*N3Ϯ{��I�$Ьp �h����G�e���,��G��o�\ �FH�~FD�'��SK�*��|:{+5f�`��ie�<M�+��9S�;���hMҒs�:�1 �Z~����N���A�q�]�ޞ��Q�Q�����:�������z���ޑ��*�F�s��<�gƩ-w�����������;�x�p�K�k�ٔ��V�o��lO4��֤3�����O-6�nǵؖb���߫:��^zq�pfw�l���?�=�5X,&�x�%_=1p?��ݽ,�L�e¾?k]e�k���p�M��Ւ{`�5�߅&A������5{\t*�>�~oI��b71�yg��|9I�� J�t9�[��zV~RT�񚸋�����eK��ݭb9p�q�UP��QI�g�\�l$�5/�R����|�b��òV�Hm*Ģ���(.�R?�b�b��I�r����������x+8�U���?*t���ʋ��CӔb�zF������,X?aJ
���k��;�X�h�Ӽ�8Ϛ}\�j�m*ЀΫ�T����$GB�?!��V����{c�7g*ߖ�G����s,DíP-��5�-����s����C��FD�x�#�qN�S��6��(:��Ƨ���\R2\FV��9]ZEӎ�n��N���LY���O�x�Ĵ@,�ו�sr9�]��%qnk�������X��F�R��[m������ɕ�J{��)/+�Հ�M�]}�`��2�{o�fP����H�4"��t���Tt��^i��b������Tp�@��G��Y�����ObV��0�o���;��"��X�f/w��Ny�"N����e�.�k��_sH=`W5(��oPJ�>�[�s��o��V��R�;n��ٝݞ6�\��<�[wv�ڡ��NdH���/
��m^�=J1I�P�g�^&QD�g���ʥ �"=^��g��:{���|�:��B$����b]��}nȋ�,%HD;�O�����j�j������CPi}�I����tX��|�6]�zA���{�^�_��P���Wt$�W� �1����M4����ϵ�&�3d[��7_A]��2p�!��B��ف��)p�1����0�������پ7����`�55.W�Q�hK�NC�f�F8y��;1�Ԉڨ�q~��̎��M���`�?��kY �M1�2J�]8l)!�@��v�/V�uy�OJ��}DD���KS���oO��R��B,����aC�RCT�Y�'D������#����.�(d�g{N���g��Y8�t&������zk�ӗ������bH�q��:��,�f,��	q�Lq�������NS\��C���$v��c���Io�ǲU]�$`'�1 xv5�t��jG&.^���c����6HWř��y�f�3D_28�^vtT�LA߄����F����<O���GXW��/�_l:T% �� �r�YswT7�Z>y{޺�OIj��s�{�X�2\�4�Lo��HFE~Z��}�(�٠��(�ے=�؏q�<��#,�t�x�uD��Y�;
�&��:�o�-�4�~ew7���	|��|v�e��V�1�,�B���� �;)Ī���h�ZhD&ɵ�k��2*u�7�8IB+~�T������:��X�d�M`��#$�9F�c8g3�@ɾ��[�����/0�Lz*'�[ͨ����P���_��`�~mn�ci#���-��vu��<����ӹ㭫����H0U-�g;������3f��r^��N� /�8k�x�~�E4R
��dEa���͏��^�I����k1�����[�!�������|E����G/;��s�+��jZ��S��w�����>�h}j���C��E��Y��34��'�[���OG)� �1|Rŀ��q���{:��԰ӟ{┈�E�0�>�� ⟚u�n_8=�.v��j��߰��k-�h�����!�Q���#�}QC?�İc��mÖcP��@*g=f����H�d���k*��,��  ����9��^<���P�[ěO_�ȕ�������\�US���}>tL�
��%��5�0L$��i���U��hN��k��HQ/q��Δ�s��(��#5:��[���l_ !��PU��xL�úo���L[6��XHy�>�� ������]������P����B�}7��]cz�
�G�N�h����Q���n۹(D�ln�O���b���sb��CBU��չ�g{��U�k���;����īb�|��G'�M���ˑW������ &,�7�y��|k��= �3|.cdA�/0�%mϩ�])�c W9�xvaa���B�xp���g���	�����r��0�J_>��b�ZNޘE_���v��b�U� 1�-��}�Tt#!�.ذ'�+")
;��U5�jj�S ��Ŷ�#�����%^��o�X�W*�.%<� :}Ap���?O��y��ju0�qX��r3U������Y>L:Gf��,'`}��dXh<��{�r��m��ڿ���%^7��× 9��	~'��F=���A~K��̞�0J5����^�()�gv��	PK�BC��o�� �!]	b��n�E�c�]�����'�3�{��ӶT�3�-5��m�5}.����z�{n�0a>�@����$x)���n�����x���p�S
=���ԄO2��+�G	QQF!i�~3'mtmW)R�G��ҎLL�x�x�8f��w$mA:��s2W�W��ۈ��I��s�lPr�Y�s��V}.������v�q��9~8�_���X��i��^5m����?�����Q�&KiJ������X�e����D�� 9��I���\ �C��M�Bԍ{��оew"�oR= ��|Qu[BO�v�b�'f�ok�B 0�G�֞��3O�P ��c�ᵏ: f���_΅��vv5��~h�������\Ϲ���T��٩�h��{Q�Snw�Ï��\w���O��yS�i�٢��Y~զ`�y�(���jm �s�����d�fvO+�}x�:b�-�	8+��	����(�AEg4�� �"�S�D��V�[t,�Y�����{��F�k����$���4|���R�zZ7#+FU/G(�[U%,LL}C�����A���5�� ���wM��ݘ��oϊ8(��t�`Bk?��"r�5<�I�ȹle�.��v���N���qT~3Ck�����ܜ� Ҙ_FvTwy*��r��.gH��Wqm.J|<4��٭�/��ۖ�����.׾4Ă���)���T޿��!1Ӳ\�RÇOǲħ0���U,:�ɫrw��P���b�	��y:��X��{�y�vO�X��b�m`oH�5�0�Dpo�� 9��3|L�#!�۶n�����?TY�����Տy���n>Ĭ��j���tŉɽX������E;!�b��/�V���9S��K�!*˹O�r�P�����N��D�~�4F|-�����V��3�f'k�(���x�(�m�Y�`�:�䜋K�^|5|V-�@e�������R
��q����͹ ��[Y��4��Ή�X��杗��I����!��f���lD���g7�>���h&d���
U*��11���u��)>3^�9�9}WX�|��}�cM�vH��`����4G�ca/����O��1�;��&��ņD������<�>c�:!!�s���^)�#"�~G�3yN��S /�u��"���^߄WGER�]ښh���]��-!�w���3���n�z��}�xC4�8`�޾Gt���[sH
�"@Y9�\r�N�t�v}���@W��Z<���l���F�_�Q\��Ώ-䜘�6��/i�
k+���2?wYV(���8�Qn��ZǵGc��<�ݿ����x?^?�����z�ޟ��u��@�� �4hJ�FH��ρ�п8.������f(�Ҩ���`��^�&J�-+�i,׻=l��
�}����mҲ�h-� �n"?�7)��wob��αe�L�	-Z~�T��.�D���itL�"u��F
:#��ÃU�=Z������St�El(����ш�oi{���r���6�_�~�o����g�]:����3�B���ĸ��� �"�9��2\�r�� gԴ��o��?�����L{oF;򨱱e���Y����RO��M"�அ��@�@`��/h�o��,_Ӯ�~�A"%���|�ʪ.��̅grU�WKr��$���K2jp|yO�_�o��EU����(�N��;$mS�#�<U�^�f�2g��̫ٜ�e��V�ĲΓL�/K��>��L��%�nʒu�z�E7H|Ts��7�'	Dd�#�󹆜P|���e��=lg����.?��x�) �t�a����=Q/�xQ�*�Z�~k�^騠D;��Ƕ~��c�5/
��b����=��"��e����0A�!�����<q��A�����+�蘞��>�l��x�aK0[E���5����9Q�{����R�	l�����P��x���N������t�DGJ?5�w�X!�,�T��F�qG`��#�����Nwmo��8w�Δ�V!��0��ܺboMȑ�mx@4G���ٴ��3Mt둋�k~%�+���#���N���28̊�T��U���J!��V�>��q�B�rBN�Y,M�r�ڶ��n_�V��t����'C�h���N����ɉV��#�vis��f������a�A:X>���؅U�,�8��鴺��~*�|��ټz����kM�d`Ԇ�������ǕLZm{Hc�xo�s+���w�;���g)�KȺ�+t�&�2\��*�j���m�!'��'�R���l+��� @S����i��m���Y��Y�nٯ�&��d��I5����������4���{V������2��5b�.���@�.���|��y��3P��Z�?��v%�0�Z��~6暈�d��o�*'�l�9��L��#B������G�	^ό�n<��o�v2�Ձ:[Y�
����T����T�q�����j���>�<��I���E�-F��j��1�#�>��p��G�^�����ަ|�y·���S��O���b��6^���p���=P�l�i٩�ؖ�Av�w�9U(E7d/����ZJlb��X]��a����+���H����}�f���Eך�-U�-��Ʌ�F�S6�!w[��Bd-�#R�V�{������cLܟ�XgF� ��]�Ԧ�?�$еƕ����ܧ�f��޸<xB>��C�����`����H¦nw*�W�x���۫)��Gu���9�+��ۡ���,����R��X,�����hz�v������)���3"|
��UxN��	���x�RL�0Ej�=�z��� ?^��"��l��5\2R�u�&J6H^B��	%J�Kf�_W�)��fp7���|sF��r��ӃFv�+G�9E�QG��P�T�:T�F/�9D�]2��	���O�lw�j���v�`W�,`����ұ0��Wj�q`P�/T��Pؗa�kQW���բw���LQ�EN�l)�̏;#�:��������7PK   ���XvnG> �? /   images/61f4766b-b131-4d1d-b591-12c82c44e54c.png�Z�S��Fw�8���k�p�����z<www$@��ww>��#��ں�������m���:):�"HN~���I���4W�88�7��K�5�뫢���o�Q7�7����Ъ����ݹ�֛���Zʨ�tM� RZk�	�u ���<
b	E���X��g�ab��<x��~T[v���g����U���ϟO�BcGF��M?ͽf��ISHCKC{ҽ�|ۆ�
@�"5	�}��� ̸o��QÀHo@�/�E� Ը�w��2	�päP���qQ���	�E������a ��I-)�bZ�ÏYK�>�j�࿯Y�X��kԿ{�T2^H;daxS�<wRy\�˄���ەּ���m��J��������2M�L[ ��],z�ҥ��%}�Ȟ�����^u���޾�+�$*��<���U�:�.�
���f=�X��������4`3U+��¹�)�5򴲲{/�K�]^K����j�{� ��u[�Z��E�����ά����͆�)Ѷ2� ��}]N̈́t�쯦6��91[[69��6���Ƞ��_�n�	����=���jS�J���-��̘�SzP���<*����:?�z�/rz#��Kx��ǥ��^�%ZFFd�ں��Q�M|,��)�b�է�bB��ʒ�]/�/�Ռ�X��>������3o=��A�:L�S���q=�o���KLL����0�]�E�y��R�
�����|v5���_
����d|��"���ev� i���i��.�H@@�!>�o}«���`Z�m��E��H�����n{/#��L��e�� q��ß��v����|��<���b�6Cs7�?C��K���c���Kfff��M�� �������M;U��V�u�KB�z
n�L8�=<<^0 
pԠ�.!�����:����X����z�2�d���:|��A'�����2�i�?e������+\M�%oonZ���떚\-z�M/<� Ԙ@1�±F�cy]�{�>e���)�LŘěZ�vZk��ɢL�Q:�u�����[w���AAAcL���,�Nl��b5�TI�z��lllQ��u�oP¼��W�,��N��ŚJ��cn�+O ������ ���:�������V�]Lf�v�DX��a���\�9�����E��VF!��\S�H3���7����<�}Mz��X��6�M{Δ�/ܧ�Mv]�N��	nRU"�zk�@��FF+�E���`�Z���-uN�h�I|��R ---������@R-Қ��E������2�g��/����qf�T��G#/���d��_�q����"#��Wm>t�*p��]�a��{�|f����KT��<��M5���O��2��ҷ�߳�I4���fg�+��F���؈���q�t>F ���U.��x��E�F��/�oL555F}�T��)sYD�R��"nذ�W�u��M�Y�v Q��.��C��!����4C22Cv���	[�����n�j�
�KmC�����ݟD�`j��ǽ��P����0>�ב�������L?\꒩gYYY{__���_��ӓ!��v~ޥ��H��jp9{V��qؕ��rO�н5q�|�t��}���A� )j=����m�#D6w���"P.y�������$� �� �-"BZ��rk�ؓC�^����-K�Uٹ<�=:�^_����GP*(;d�'�^v��#U�;	.���U��잲T����?��]끊a0%�V$q���cYc�C�篒D1M]]���_ �`\ksWWWe7�R�4t�HH�v�㿘���m�����!~^���>)�KQ#ˌN|c�x::@�H���%�|fƍ��A��O���hZop_�ޞi��90t�oTcZ+Q�����634��*� �zA��SH^"�
7=�LK�2"X�i7&W,����ep�G��&�_��g���|ٸ�k�dN�l|�WE��������X�ߊ���R,c���rG����Đl6]�^h��IP@U�J��~O�
1-=i������,Hn&�����%G�����G�p�4��Q�|�ɍF<��/�c�,_c|�Y4�0zuv&�W����I9v�`J9?�C���q��Z�����������q��\\[�!!&&�"%U�K�b��x[��<F+E-�ec���"<�7��'}-1�ow�*�P!������ݍȣ�˒!�RMH�%��/c-0m8���`�Y�a�ͯ���� �|f:�*�k̒��B
<u�&0��,�K);N�S_o�/!~�oa������N..'���O~e�-�ES�Lސ�ˆ�nspss'2�(�����3hCE�,�5F��Jg�X ce���ޣ��98�WH�U:f��k7���1F�M͌��f�&[�/̒G�s�b�X> �zd�XXٕd�s��������Љ�q!]\��lZ2y�+�6.*6���� Ɉ���X��7O.����n��7�p*>�YN����JV"p��T�Ε�/�V��2F�{��������_ Twk�7J�fb���W?�n�M�a���r>��~{s9�����K�2�G3=�ɟY���E��]{��g��5Nm�8*���7��<Y�������mb�f����^�N�:?�Z�ܧ��U|��:�J���O��q�ڑ|S.�P�͑_u��☧���7*��l���������r�;}���p퀈��;���`Y�X���G���-���:������R�#�-��fFIA��%��;��iSC8����߅�J����tt<���:Y[o��<�mmi��'�'<����@Hf���hG�,�e�Tx#��$b����E~jx����5��Z�/���Q�YԝX�2�����)�)$�O+�tԖ��1���(��O����_�6�����OO_iŃ_P�?+g�d1����D[�����ޢ�va}S�?k��o	KHH�ʯ777_{�{>����]������Ξ2��=㟎�^�jT뭋����7�N�����"�j��u��:�-�s�Z�}���iy��ո:2�
��y��Ŗ�w;���/�<��2�o,���ϊ���{�|x�������=>䖓�s]��D9a�񆑟�����LH����K�3{p���)BJ*�@ >v��܃s⊅ucCCMB��8���c.E��`]�y��N9��`��� �nf�"�c	��xǿ:|P#N��@^1�q��H�e�y���8�MW)�+)�d����Rxb�s�r�~�D�zu Q��?9����#��7��)�;t*=F����v�ah��e��8=c�N��\\�]~�m���=���!ǒn%c��=��M�Z.l�V�B��"�s7瑿����~��χʉ ߤ����-�*vQ[0FuR�Kno�4?K��%1�S�,��jU�	�4��Џ�ab����D�/w;�����^^^�^�`���B�[.>�_5�2��te���BJm#�-.�5 j�71|�<T�b�'O�d��F�u5�<םe���|ڵ�KxT�^x9�7���J_��29(�}����"�4t��ͱ�3�_��|a�G�B�I�����'~G����Fs�C����-ɵC�8�	��cݟx��%���h-	�H�g�+29T�����%�$�jd��ldo�0��+r0]�Y2%A��g�$���MѮ��fYE0�b�0h�!�Z5��%S����#ޛ�\�R�7g�3E���[uls�Ax�Y��L��
TZ����k���7��#&�Ч�陸�?�k�D�1�T�@u��o�����B���I&߼E:�Xk	sc�v$���G��{���O�����������L�q��::�E_�U��R ����'�� uv���g�aBc�Ck���ॡֺ{-<��x���PE��n�9l~�ٹ�M<�#Xo������Cn�(�n&�\���'�Yz��<e�K=}�؃x��t��Ļ��&R���ϔI���P�W�@Lү�5�>�Y������*����M�h��y�E�I�)I,D1�4�\�3���|� -B-n��g0�>2R����3��|Z4�d+��\��slj�����Kz#99��q,x##��nȘ�����>���a����y�	<E()D-��Ȋ�#F/#����U�A�	ON�|6�� ��-<<d��1oN%����n���
�f�*��<<tP�'���� ,.�D'�f��ۂ��tx�]�� ځQ�դ˶�W\��g�[1��f��~O�5!ݭ�i�$Y�cHPMm"�W&V��B���;~�Z�8�2����߿����a��a�x�`?O�$� k�H[�;�W� �.����wF���W�Qi,p��֟�4���+^�uHvi���f�т��|k�u�ߪSb_8�9C��*b;7GGco���3��z�f�p�,d_n���*��cM22��l����o�F���"�d���7����Դ��CJ�ș.��B�dsZ IMu5	Twmr2!g2���% 9�C���jQ���}R(Qs���jsGGM���@���(#�at�V��Z�ુ�H4����?�\P(Y9�sz:���|�F65�7�<Ӡ%ZcU�cZB��Z%J$!���ݏms_�;��K?�nKs������{�y�2�Ʀ���Y����F5���s1B�w��'��&�>g�w�_3҈y��*�a�\	��2����S�V�h�Q�c��{p��-��V6���4��98H݋�<���,������٫ӻ鮅BLk��M��D"���_0Y�l "F�98(������,�NDl�Ai~����DP�)Wķ���vƋg�t^�2�b�)ڸ[�R�|O�#�I [!$oon�Wҫ�=�~@� ~~Ԫ����k��(�	�h�UK�>I�D\�ҵy
�W�����3�U�[��2��,!E��sS����������qW��Cxs����{Ū�q82*�L�.��F�FRq��^�J�7[���I���9� B8��,3�a��|�+V� *rr�p���l��4�=b݅�u�Z�oz3F�HX(�9��n�ce�	���K����r���bN���V��S� �jNA�q$.dk��c��e��3	��N5P��:�6�W�,��m_���M�m����Ee	.%e B�-�X%8�3J}>#kĆ���5�]q����Ro��Hj�wt1ʠ_3��!�5�@��n�ti��F�|���HAl�#t � G�c�L���%9����$�[�D�F���� Í��;��nOO˰'�LA��7���^F�mn����t�B\�Y�]�~7���H
�Q��ɣmo�?E�o�*ML��1��<��Hn5��5�7{�b[�;	CkL�c����R15�T��deeL�#7����^L�~�C�G����Q�:���Y���
�� zτ2[�f&P!x���C�c���~Z&�ڴ��XzW�Qd�� ��,m��Q6#���*"����0:���x9!��B���ڶ���X���^��[@־J����}����堢���5
(���������2��k0�\;�#>j~�a�UR�n�$����	Uvl�thL�7�	��#��>6*Z��1^�=���ۅe�޽ծ3��PP��N�J�!߸-w/�0.�4��ة��#etB2��`~"�D!�|W��eD"��#J����&7�V��b�t�(=Ӿܜ�@j�����x��,]B]d��-&�����H�z8�vYv�� $�d� �%l��J&+�t(��m܄��X����|8
�045�J�5���4�8��
��hM�~���G0�G���\��]�[͵�]_�f:1�9_E�e9�z�5�{A���߭��<@���n��^:� �e������+�V,4���i#W{��Y+�GLe�2�/竑VM��?aY�\_��#Y�3۪�,w7�h.�Q��+�/�:��覿1�����P8�����m�S�\���F]���Z���lQ��C�G{�X?�l�����>����?�;����n�Zu�Z��N�}���L�(J����4�H
j� ���@�0���e�	����"Ke3�^PIկJ����vH�j;,�e.�U#�D%$J~��V�FC�Cs�qn|���8�l��O<"�{�)��m���x�W�BDj��D6a�ل�A�D�A�D�S<�ꞻD��%t��F@0桸&��8$$�\�H�[��5\VmQ��R�U^~o4Ԃ-S5G�pː%��T�~tx
%A���6 ����f�K��t"������vi8�l�?�r���̢���T��fGuc݅���I�����K�;{:f�j��Ήt�Yd&B�1�<����q)d����)��@r�n�Ȓ@��ӓ�)$�L�U�!4E����Q�c�챻
����Qz��刺�Aࢭ��M�K?�'.bd�]����pJ�ӔhyTtp�7t�)�W�Ү�OV}2ũ�P��n�
J(�[���Mא1w�����
��m�9����#)M*����:1볣͍���'�~�ed$�>�4���/���{b�3w��
S=�>���� �ٖ&�p�߭ /"���q�����P-s%��"н�"��ʒk���m�s'X��[���Z�o9���h��Y/�� [��Ą�(mMݱ�O���1:�䒲?���Ndd�Db(U�z���5��^���{����;�z,�#�h� v���7r}��Q+ԗa�j**i�p�aW_&,}��D��c� �|��Y�#a2���Ƥ�y%)����� q� ��7���4i�3��c�Ps���?���O����(�È�m�д�[��H��N=9T�&	|#Ӝ�~q���ܐe�j�*Û.�ʁ����?�,�%�o�W�p$9t �D����?/þa>Ҡ&�H��:P�?��	��ʃz�m��w��=ؙ�㪆^,:F�8��^&us[�93���uQC��G�4��%���� MY|j�z�"	�z6N臅�Uő��WvrS[Q�0O!X��$��^�Q7ѫG�v)S�R��=nF�>7o�*X1:�c��jI�&8'���>�S����\n�r(�,��$0��/�j~uB��=�O1q�E�"�ߏ�vL�ڑ���'A��@��2��!�=z6��(eW�93^?g#��B�����Z~R�GO����8X�<�ޤ�k߉&8cF�)ю�k�C�(~iȋ��
��U�l�ݛ�mx�ɼxb�8�>۔a޵�^-PLG����gF�Mc���}��2�ŏ��ؽh���D��n?t�{�I#Kvs3{s3R�8��9�zxQ̱.���e�W磌�1�%��/���4�/r�!i��V6>���\+��h,P�8�M�ڕ,��]��l��Ƃ��C�^�[��|�>�4٢��~��wa�(dO����ND?�KLR����"3����Saj�Ej��p�j\�<ΓG��BB%ru���j�ins��<�H�`<Ka\H`m�L�|ҏ�ڜ_�>aѡ�fx�r�A�����+UE����+( ���S���(|����,���ڼd3�oG�>L|�	��̇-�V���ZT��
Qy��7;д��#��+,$���*b\�g>[����g����b�����y��٨j��ک?���;$j��`��H��\�/=�w�4B���*e��7��ڭ��K�1uŒ���E��3��4s6��E��JS����1��[X�}zq���C-Er���,����+&�>|[�epi� v�P��|��~!KU����{��*�/9%%�n�y�$�߬#ؒ���m\^��yo�P�6�N�X�`��}=�*Z�ێ	[%��pG�Ǩ����Z؎[&Up����9��a��#^��]�;��ALn���Ul��]�"�{�f�oق��jM@��
_�W	�Ҷ�Ҋ/����ʜ���SlZ���'b�R2��ɼx��������Q\���u� �[�}��@G���[��-��fTm�eꕝ"��/Dբ-`�5�g��d�?�<ۢǿ�a�z89��G��%~�Ux�)����1����A"�HPS�Qj�E��HܻN�$�N?}��@cZB/��e�zsze�ck|�(�۴xp[e��n
�
�����W:hv�*
��Y�"���;X�2��)J�.�D�t��A� ��Ζ'�N����r�[�t����&h��;{�L�
h])�&�"�
v�����}�#񶙕s|gt#��x�xK�r��+19����0tW����CjP�~�}%�o��9n����g�Z�>^80������	]*���c�	�Љ�ag[������R9�$y��&�LT�/�?j�^{ѿ�� �B����K�,�~�,�l^|�f����,[qq�P"q���{�̠0�%��U�7+��O�P�����燞�M���7�ry��.;�j�q����mϽ0���Ͽ��MIۡ��V�@��qҩM/����	,G�OrGk��F����JϙQq�8ѻ���H1Y����uW��/��hG�&�����|2)���'��5$ͼ�4�LH�C��_U�sTW��'V��q%�>Z����m�sk�ܾ@48���������nx�6�s�s9���oJ�_�Ů���7�9O5.�J�:�e��Қ�4�d��i+W����m4'Z������Dh2�����qY�fk�����yԒ����P�C��/L������:D�<
J�ܜ�`x���~vb3��O��T�1�=W�
{��ۅ��˦<%��Bw���>�Ne|3��b�K�-E=�����a�d��|{�Lw��wY&���t�z��~&���Ag�v@�_|���$���-#���`�/G����2���ZK7��G�V�3�.�H��A� ;������>xE3sxu�Ђ?t��w�Y>:V�;��E����ʂ{�-��xv�B,�n�\��Y]����k�U�ȋ�������?=��&��9����d�$��l��֨Ӷ�)E+�K�YM}v;��ӾpV�Tu`��'c,B����FRQ�1i`�%�I��,�K��F���������;�@�'��f��1jpL�q�D�tP��a�b;Z��6D�DB	]|#�e��"ȱ��/��+@;,��ܢW ���p��I*=��_׌��`�����l�F�{��|v��7���jy��NZ��b�hC*��m�5>$�CS.~~�Fc>����a:��w0W�E�q��7���
���J"|�rş"DtƵ.��*��k�ՋB����\�����ҧ����a�w�t�v��0�ݿ~ 06��Rڰ�F��̵����}����ppm(����a)0V2�
�m��W����8
��L��զ=L}�HI�m���P�?~����Cf�ҿ~!F�Dж��:���R���
�Lo������;�EYb�+g�ѹ����3� ���/٦��B5�tlo�1��v�~�	̖������ ��D�_c�7����}i��^�nj^!*>�4م�h��<G^�ϿY�(	Vo%���Xok{�a���8ڑ��k��[�'�9�c跃�4���J�����ٯO���hZ^"q�/��͒t����aJ�x	�j_��>�7o���غ��Wn��&�U�z�ǰ0]_��)GZ��T����-�|�F��Ê��z �[��̮�ɡyS���,���@�822�:Q�����TZ&Qq )�޷ �ɞ�ԛ�R�"t�O�ΰ������������(��|� ��s��_-�G(m�9_tǯ�o�z͘�~Zi7���FS����Es��$|�Su�����H��D�d�^%'�␥ ��_W؊�9�������r�!�������gl������z�ϟ?T+�,/���<�O���#o��j.�m�`z�:-'��]\\(022rV׺<Ik{�$Ns���wq%2!�q�28r��b-�C(�[���*�A���K��txat�	x{x\�T�-�I'@䦅7�Y�}�u�㞷�_���?��a���8炋�4߁$ū�_��5��n��%2�lR��8z�`�f������ה��fc��&���y�K��wu���ȸ^m�Av�DXly+WxE�3_����(�4|��	����|�a����r,�#�M�+?�˵ ���	n�����6U�D������Q���҆�99�ك̽��׷B�Df� � �����9�fa-�wk��:�eU�o���^��K�A��J���Ju���sugg�O�!r��Y�`k�r�?Ԓ��N�ʯp�Ɔ��SU:q!�D�+�:�?����*��p/�G;:::*��,|3}�ZO1 �t�BC�k랖�Z���7/�}��Dƒr��I�����*ć��������)�a�L�t�Xc1���7�gm��7����<����ǌ�)�gO�[���%�Lܐew����q�y�'�����N.���4_33�����V}=��:��"~i^<yymy������ڠZOuU�zotwAQ����R=}k����V�PV��𴨇86nnZHz���N{��0Lĥgf���<z�Qp��K,���ExA�߷�?!���s����Y���Je&�9�1`�'�k�hq���mg�ut*+�e���&1�� 1���sc��v�zϪ4IT�dM��sus����-�>�\v���v��ƺtVؘ�2��F�G����,ٿ�$�z�-�)��L��Ȭ��-��P�NV<<g�vo~�\��.����������mc�U����U��'ƶ���Q��`��ن)Y��-�Β�:�w�BMx��锋�di�їQ U�ݫ��w��r������y=>n��`ܢ����};�8Z��"⫑�Q�ݴ��v��7��׀��/}��W�J"�*�\r��@JA�_��XU|LP<�a��K��1�s:r�6@H�R=�tG�K���U��)���(¯�Ὂe����.����۷o<��5&xT6����&]�VS$��4�Ѥ[~�3�V��;ꯒ1���dğ>���ۺN��`c�uCxj_�{�6%pU�%�O�L5�:��%��Uҡ�1E̸��`:�O~�����f]Yg�(t���w1�dE8eB��w��p��{ǘo�%S��.�����Zf�� v�
4-��.�_���,:��ܭ7��_[SYY�����b���O����.���x���>�+�֔qy��yq�7ׂr�r���9}1%Vy��O7�5�Ăӂ�t�f��R<]�k������Z��ğ:�O�_/y��t��s%�W��p@�(^��
�ӫQ�8�wX.�'�Du��D-3��kXS/n;�I������Ȗ+��Td?�D�G��֩��j�J�6��^��������%i���tX{{Q��,��v�8a8�e	\���X��ʩ_��D׎����!����7�b``4'&NA�Z�m��z������N���oF�g���=aa�������:�u�?4����)J�*��a��5�( 3'�����&�<pwii�҈���5k?����L�B0�9(HI���j�+�����c�q6 f�q��T<�@a"��4��θsu�듍ͫ��]]��}�3��L�EI�z�,�7�n~�!�u���}Ā��eA:�ފ&Ű�g��F���|+wD���C�����%pDl2�ڌOU@�q�ߴZe��'}gh4�����U�����.zf���t�bw��t�7>M�g$����g,��k��ӡ�݀O�$��#��-��w�6^�6uY/
˾�c��(�<HO��T����3�?���b�A��'�/`B.����S ,<���2H�){wſW��OlS�R��۩�d�
��@o��~1Qb��N것��:��mS�����N�������tr��*z�mR"��������M\t��1�UU���@k��p�~E(.:��&�4Ch�TCHƗq�'���;Ġ��^2Agb��ݝ�2fp�c�3��Ay�Zk[[[��� _����碌a�g��6{��nt�mtCbm�{�9���_ed��1@��G	u�5������ WU�60v��=\ ��;���� LB��̻�;,����̵�9yG"� j��f�O��(lUmȑ�@ +�?l;��ω���y7�W�����T8�.�5;�!��:�sQ��I|ϧ�y��F�P�0���R �U�nŽ����a�4�;��ѫ�m9hȥ��� ���p�����d�㯿�j>q���ūJ���w�k>"C	9�;��� ��|���׫k�l*�$�fS��pB(����#U����<#ga ��d�C��4��ȸʼ.���Z���P��Du�''!˥%�:���ɺ����dPrgC=b�C3'�̎�:m����՝��4�^�8u6]%��q�
b����#-�@�Ƣ,__6<�XC�R��mvX��^Z��UL�vp8�V��,t�q�B��ۣ�=]x;�U.�_�`�[M4ꏏ/�N[H�E3n�<<<���#m�$s��e̧2�GHn����R���\�_M��-�@nnj�n�A��/�xpp��2����9�n3Kv?�Er�6�}x����m�t�!���A���쮙,\E�q�����DTǋ~�G<Od����9�%��kX8�%�V�X�reO�HKL�Wx ���^��v�R	�gF�/���Xc�>��I`<�2rK���d�}���[Ѝ�^�2�n=<<ĳ��P줓���ym�5��/>֑,���ӵg:M�.���X��U�!hC���B�q�G4��k:�U�����4_n��>���W�}/���Zl).裚��U����U'���A<�}!ax3b揹���k�u+v����d�Vľ�y��F���b	ԋq�bNA���� C�cP&�Y�0>%SD��f=;+^�0NJ�]ҩ��ڪ'D�s��Z�1�zD�������<����v`�_�����pF� @��5���˿�(���9Eozv���7su\0��`���������C�{R�kR**?.��rϡ�"8��==������2J���X�5_<��-?�g9�&���`&Y�p�P�< �E��<G�\�Q���軱���8ö���wxn&{N��[q�BK��G��hŢ������
;��e� ��J���)P����*~����u�8�(�W�X����N�O�N��	�ڽ�GZ{�h[�=%Yx�n�ʿJ���)	�������NU:�9�u+���U��a?N�6s1c��Y��gst�s�]��6���Zh�Q�W;�5o�;�a����R��	Z�3(�ω�C�i�uX�d9��g�󣦾��������W��l1��3��O.��[��٬�'~�����,ʍ^������/%P��c8�ύKY~���m
�U�Nz��m[�/<���6b�^6w��	w�_T��B�?���9{c�c�
^9;�rP��ZÜ�K��_`�r��3�V�5����a'��wۗ+T̣$�Ryy���2��������_Y��7s3\�#��`wK�M�ښ�����wX	N����!a$'�iBtF�x�,x�H���v���N{Ų�܋�����i��?gZ(6[�ਸ{��Z��x���Q�V���C's�#"�ĝ����4J����`������� � �

�8��]��)�'�����������~c�g�8�Yes�\�s7�Wr��z�J{k#�źQ����I�-��\�~><����t�������2�����m��x�ͧ׽�	2�B�!�L:��2�������6�U�ӳ`��*�a�Q�3w{�~����x���챒�b�p)���~UֲW��i��ƻ���w��u�K�=+�����q�O��o��M�z
�&|��O�!EI-�%�RJaXx��M �Dط�[W��c����V#��6@�������?��/$?��l����{<�-5ڼ�k��^^z�,4��	&��U�ʼwip�_��/DV��(�,>6�] �w�:E�Zo�w��<��h�MA�o�e��Q���|��*��iQ	Z�$-A�m���C�+�x����^G�\,�ξ��!�J�#�1iP��kp�}Wh�;�/�d�L,�w�2�l'�t�_�c_-�̒^�v"hZ�o�xe�Hd�o\��!.���϶pvEv^P���a?�������dɱW�ȼ�DA��폺'pO.&�gw\(Q��V��1�i$�pÑ=<>~�dIp�m�h�Z�	�N�ȴ��Ҭ���&�q)*T�TOl����t�ޡJ������I��J�k͜���!Ͳ�>�k��m'�!Z��:��&[i�;p�"+�Ƌ�!;F��s�f~Z��`�&��f��Ll�!X�F���4�s�ҷ�B.�6ߕq��La���|'�pY��#‶UC6��.WDd��`l<=�ɾ%#�ǧ�*��d!i�s�Z�9Ņ��5����q�O�i��������g��)-F�5r��2V�zW�Ln94�*Zl[ƴ#����!������y�5A���d�R�"�n/�q�zEZM�7��*�~.:������P~�K�P�>9���k�S���Ҧ�2�T�w+"$T�aڵ��6�s���m��hn?M����F�,�ҽ�E�9b�_�ޚL=7IxtX��YKH�=~�;�o���;껕����d���l�|���&��&i��*J�&����6�^7 �уzqq����/�/SMD���:���?}d�ѳ}e�Ⱥ�M�=���bЈ���( ��ħ��2w��7�/Іǎ��X�E[RfM�Խ�g�X��j�
�Z�]�}�;=���#�Ŗ�S�IP\��J=���E�5v]�J�*�s�k0��/���u?�ʾ���?Y�SX����:*�M�ycO��ؘ��t����Zj5���I�O�^��zd��@�*���)'�%VK�GDd���k�Y��%6o��b4E!I�|�Y�Z��"�W�ZL�j#2�rF��&�~ �Ҭ,��>�J�ʻ��m3 �t�ޟZ�}}x@��6�sC���!�$���n_������P�ƽ�ƊhW��] ��<Ɓ��,O"��-/�rjK�w,�U+����D��k���Q��1>0G�њ��D5�V��A���I~�ғ:�(���u��1�e��IX	�����ڋ���dq�F����Z}@��XH��;�:WIs�$F�.���Ꭶ�-E�co�yg㉘5Ux�b
��SH����b���$�I��ToOz%��5��m�!�����c;K=��T��;���-pn>��Z�����v�sn.�ai��5��-)!Q,:mM��cS̷���b�v�y����xW���٥���@v��y���W_��s��FK��hA?�����݇4�_ ��07�7Ŧ��p�w��^t$y�{VP/�G�h��!k�PD��o�����(�Z�4��a�9��/���h�d���q5� j^����0-��8��P��q���U���o��ӕ����^Y�C�������DEh�%�Y�d������]�|&lˢil�����D���i��K�O�S䡻�<E�)-�	mO9V��}�u%(����a9�\�yDFF����y��]'���p!Wl"�:f^�O_�r?�����C��-,"�M��ӲKaM�����<b�����U$�'����5�C��W�".�ؙ�/�>}�;�.6P^�����D9�}<o~&�}e� �H��ktD;(9I���a��'N3�^8�I����q���5N�������A�;�h�~Eι���/*�ķ&z��Ԡ���8����u���R2a�x���ܩ	���X����%�ׄ�E�Jt��3o��uFJ���U���k��F���[����h�H� ��d�b���}��q��p[,�N�h����I��ⵡ�W�D�'�ّG�ևFy�r��W�9 D����~��R6-CB�b�V��c.K	�՟�� �h�f��߼[��VJҞ	������C�h���"��I6�y�m7;�\��f�5Y*��W����d��dDeFV��W���
�f���:M���c�<3�-~A�L!�8��|���w��獊��3���uP�З��E���dt
z��0�Osu�5�NL�g�d_��������4��kF,rA�-Qn[v�;����*�sϾ�hވ�(�\��!�?a�$�e�ׄ�$9�	�⢅0����3��:{��1@�ot�����p� �$j�(.ňg� X�O��I�yR.!D��%TƯND�7�oL(#ahm˔�L(�> Y�+��'��W?�$6&i�,�,o-��Z1ٳp/���+� 
"M���l��
���i恠��������LaM�
c=�֯�0
�IIy�B��������^���~�	��ԡ�\� ^@�������Bpc������`��Ƞ
��ö����ͼ^���t����8D~䔄w��#�=�����I�o�u�vRB�}8L5�J��p���?������hK���9�z��e��.%h�SO���-�N��b��h�X	~�Ơ&I�ӽ��.%����aV�s�6\���]����џn�|ʤ���M�~��!_!ʣ�z�n���SΙ33F��n��A�==I��z���+��ao��02Ļ��eW	�R6jR%%� l�(��k���탥;�p"�vk�1BZx�Ğ�a���`��>1�v�����%�GFF~lmm�=KKK�J��� ����S!�V�5T�b��B�ȃ0�x�)#��,Z��s�=Mv)���saaVw�%�E����!K۶)�y4>WH�����ؘ��]6�n�x�I���NO�M��?��T����*����Ԭ�`h�"&3� ��@,�j�<���iȹ)�&5gw�������� ���Q�)�]ʹ7���Y�~WPŊ���ya���={�W��i��&�?S��8���D���=�(cǸ��WmR�����꾱�i���9�7v8�؎<X67�"���,:+'Wf,::��WV�q ��A/I��a��71����N6L����y��#��������3`H��=@oZy�R<`Í���t)�Y0D��������',�U�A�������CP���/�N�̑n�I�I<R�[���)�*U�6H� �`Ld�_��Z�����oћB�mp�	R7�����R�i�H���t��@h�����ku��^�@�����J�tx�G%����6l#@4�1������#�B�1�b"6��������B����u��3�֭Y=���w422j&=������%BL�m��'�JG�I�]q$Ē��R�Em[4�T$�5Bk5�Ǟ�6���c��\�8d�ARA��CbL��llrC���u�V���^mE��J��� u#�ք�� �~������'G#����ظɧ�(
ߝ�n B��� 5n�P�r�S���x� U�0� \jؕ�%3��#��S���s
F�cF����+WL��B!��rV]����i�;wΨ�8�|�e:�o��v�v@�����J}WX5��?�tNGR�b�1�V���.���s $�Ãdș���J�^����c�%������)e�i�T�ȱ��3J��� 57��%o&��k�v��5ς���89��*�,�r�y�Sԍ�H�"�Z��MI�m>�:��L$2nV�(@��A��Ĵq>[��$��X�6�HKe= ����8¸�C��u�i=P�\�����?e]�U;�U�v�$?�
G�#�o���p'6p�%�K4�p�V�8�}�����#����AR�F��dJ&�1�t]�:��f����&F FL���.g�i�V�f;�R��%h�SM��#��,�jM6=B;RluL�@C�0Һ�qs��i���A<�9�J!�Mg2D��^q�E"ԩ#��Ƞ�[]]0�.��iB��:)� ��,<�Q٦�y���SF07w]-.��\�##Ȧ4h����=Bc����~�v�UʵZs���%���G�)YEԴ)Z�c���J�o�e�}�b
޻T�Ts�w�	y
ʎCd���'�HFZGL.1����eI�;�mć=qD���*}�(�OX���H���j�v�8�O<�9%h�SM���<��n�h0��K�ABz����a3dTAcGL� -Px���yv�ױ��١��@1�Q�YV[��D��nii�y>)��{4��P̬�b�����-J�����{�{Bb���u���O����g����ܓ�<I/����M��sl2���@�A�@��F�^;ًj�u�j�E�}�;6C�1�K���y�h۰%r�,�<�N5G���T;��Ҳ)s�IH����O?��z�)u���b7(=�oh�f�gL�5	�NOO�߸qcC	Bq�	�X,^�3�
fl��c�����$���}����,��U�y��k�R1�/}�#��H�g�r��Z�l��*��XQ7n���G�|������+��R�?$�|~���nެ���O�g;��V���f�mg��^w�%���o��a�$��rJFX�Z�A�	; e�!"L�JH�8���|��vmT��-��
�+a F��w�i읞�V9���D	$~�]�~F����u�4}hh�MZ0xzff���<�̜4�����"g5Y�����g�x��}h@U���dw�Azh�,9���f̚�I�����V1�4�,w��� �jc�l1�]+��v0��HQ4% L�w��<	M�lB$)�b�)���'�����񬩺K2�\�Ӟ�co����v�f'
��H��T�T��?SIH���(e�o�l�ңT����CRHp�˹f4LW�\1�N&E�֌�bDQiMdF�����D���^Usss� �Nib�����?�����߯���ՓO>9��� 5Ŵ������O��'�|b`uu������޸��-�G}Ԕ��*:5����0�c��5��3o�$T*��E��Bl�(��<��ѢY �X��&1���� �h�fH�`
���q�<k�o�b�$���+r��u���D�ȇC�(\�'hTjR<��nsI�$��,�Vi7�X=��p�<Nb��¼�c?ԧ9S���~�{�*����y���������&1��w����y"^�ҥK�Z�և�].�R�k���I�CZ�����[ׯ_/�S�M���q�~�?�]��]߷��6g��&��>�N�CV���/W�~���C=d:�����;K��z�D�ˠ���'�')�`a��,l;���:�Kw��}����Ai�4���(�Y�����I\6�t@�؆
�Rk*+P�S���D��Z�����IauW<�^��ɶb�1��[ܨ�ya�j(\�+���X�{i8�V�1`-�)Mx)�&�WԥT,=������+��c2}��EC�����3ƃv�$�^[S�n�R����V1�|�+_Q�a���z��e������+w�uׯ�J�_��׾�����?_^^����?~����=�8qy��w�פ��R��'G�^733s?f]�Pu�ᇿ`b����7UH�gh��=����ƍ��&@�q�v�8��ݑ��m7hV!��a�T	[��6:�z����C�|đ�8`���C����D�nR�!w.��W׏�RW�����-���&�#uf�֠a�"�:���CN@h�����s��7Ix	W� �~
��n:?��"��2�D�"�������n~W+I�q�P�B"��8�m���ýi!A�w�}f�!^�W������|�h�Ц���Y�z�_�ީ����ٹw/..=z���?�v���\�~�:8�g��ox�mv��]###�ֳ�,������88��cu��Y�a)�T�m�h` ̗��e�[�����W��Y�)Fqm��d���mV���q���s 5*���+��8c�Vx9ZﻓI�x拋�L�(@�̶�0|\P�RLj�Q�FD�.���* ��I�g��z��܂K��Y��KvX����N1�{>|&��9�gb���aa놛�)�N�k''�G�+�fh�T7E�*��UǮ�G�s�����w�� br�ܬ��{{�'L:�׼�5f6��6I d��<����-@��r�̄���z�&��={Ƌ>��/>���x������O�l�����8w�&�w���[s�ccæ�.//��W�5�7�}�sMcE��K�na@�y�Ha��g>�Z��>����M��*���;����A	=��bϸX+9wl;��g��[1]�/��P�jb�	mQNi$��!91I�$O���V�֜p�,�xC�T�*1�#o�������τ�Df˿ů�K��s�W'�V�z��tz'�3�J`A��w���ʲ9��@27���w�>=��g�5a�tA�
B���6�W,��׿��f�8`�c�<�7,A"��׾�5-(|����k�����>�գ����߽�%�Gfgg�ӟ��Q']E��5��/�-.\�'SSSY���c�=f��x�?��?lH�6އ���`���ozӛ�B��yAPȿH���������ҢwL���cl/<ة����7� �Y��$>���& �Y��!L�RN*�\0A�����a��%� y YC�{��Qm��|���VS��	�7Q M44��'1���A�o��n#��̓^�������[+I�qOP����i�	�~��^�z��VU�jZ���8�1���W_�җ�8[%�>�c'Ϟ=�M����;���T']A�zt��+W~I7����&G�Yk��\������_�B#-�mh�@�B��{L��O>i
T*��CN�"���@�s�ٝ��ٮ��7; �⼒&�5l����m�g77W5��]I�r8��-MxRq�ۺ�k�#b&��[�3#ۉ �lG�#�����	v��qn��y2���Ғ�\�D�# 	R��^�,��L�FJ܉$���}�>�$��^�3����ِ���w,�@8�@ �$h|^��5/g :w�ܛ/]��"=^����Cuб�	iR��wh��z�r	3HJ<���we֍7�J�(��*�@1Ic�F#A���g?g���蕑��~�1���1�35l�J-��yZ�n�0̊��gX(�	���,��Y�$�7�ނ��N��MXp`x�b2 �{.���BD<"�r�6�̜5f��j�{����}�$���{���^�F�i�-oy�јq2��WQb��������qjf<+=�N=������]�O~����rtA�?�I��l�D��\RD�eU*\��@���w�B��8ض	�<H�:�ʤ e�_���}���;O�v���g;��V�Ta�?�`@��4A�P�}!0���������2���y����$�+A"h?e�$�X]]v%(
���Pl���Ϟ;7��]6��ݨKw��Ò$�w�~��kaa�,���$8k���,�:
���1�?X0�_t�CӦǑ�w�w�_?��'>��U]��!H�`/jb|������L�	e��r����ڐT��¬��$���g�Pa�ڰK�~�΄�"�p>�⬰Y���<���X�,{U��^r;�����}Ҏ�Tx�mT|�lf��ˋ�G'��)�dr����W	�
AG";�4  �R=HH�Ђ�J�r��L�q�!H3�͒T���Ȑ�4G�ݗ�ګԷ[����h��@?��B�A�}�0y��:b�Y�)���ׁ=D��o|�L�!e�:�%��ևT4I�;ե���R�722�64`��J*�d�O�N��/�H�p;fUj+Ϭ�!�'g�`�*�=R�7�`WW׍��U��C�B�ӹ�O;J����K�P�fؼ���P�hss�Wg��䍇�w�ʳ�RX)缴��d�ynJp�۲��${ Ś�����%����{e�	��`��Ǳ��>#��7eoR?�T�ı��{$�����Az��&i
��Bcc  �c&�8A�Y���/6�ЃJ����Wx����o��\��Z��-�j����@u!nA�wF⻆��~F���F�Ⲉ1+�a��Fj�}��:|��>@c�'`�uD�d@���n�}�sN�Ȅ�-$ef��	���G���G��.-���Pwb������H!1�1s������7�Owc_l�x�8�����f�N�ڼ1�$,�_3�7�A)l�P݂}Ip�L&�Ξ��퇜f�<�u|jM�U�&Iz�jF\__3ml��
5��M��̀M�<&�<�;��_0{�g��� ���a"x7�}�kA��0���/�%��^�z�A-ev�w���e��ο�/�'z{{#DI�:���!��%c6��Q#�Fi����ɞ�)�l�?}n�th(���RR9+er�BK�}ѐ%~ p �}�Vj���4
�F�W\���K�L���>3��d��Zq#"t��=�:W���8բS�Ma�21Re�������|�����>�ظ\׃\[[1m���՞�KgA�	�g�A�W�M��$杫�n۪�]<�n���'��k��y6N����	�9�!A�PJROyZ�M(�F��u��th���AV8���#�Q�m��g+T������~ޮZ���&�T]�c#�s������\�zI�e���g�`�zw�HE�8r��4^*�M�A;!��zնDM:14�ry�Hd�y�3��J�U�����`�ۛuԗ	�}Ķa�|����S�!��1��>�̰c�s��㩳<���5�� �-ϋg�}}9'M������>�0�����n�����'BԦ��d�mc��M����r{2G�\��dt!���۟=����<�o�xx��qL�����H����oя��6�D|�8�Q~ޘKl�� ԩ33�݂�^��6�%�	��Ȓ"�3�
Cf�$T���� �>~"�����?���{����w|����U�X�ҥK����~i```z� 1��іA��V����t&��}�s�m���;q�z5�\�{�@Tr��G�%�}��dJmn�:��*�S=;,���+���$�|`.7��+��;A�`��%�jn�z�/���F�v�I��B©A�&����漧 �NZ5�vN]�ߡ⊗vΎs�Zj�`�����.^���S�Ԟ���{O�m�^E�3��W��|o�`�)�"l�l���c�oK��϶��Ǆa��󬶊��ܯe���}6!.1����O����'?�I��W��m�y�k���O}��U��H	R��w��~ ��vF�/
�����VqT�X6�ao�ĊF����K�h$�8��#q"��2�;�Y��G�M�a�ż�WP�`��3g��ң;̀#z?v�x�� �mhhL8CzPC(O^@�n�[ʠ��q%��d 6l�����v#�?X�;��qF�S��3Q�$��֕a؆�Z�u�`/$��Z���X�-4;��`��6�Ahz�� G�$O�2RǍ��6Bۍ���q�5��|ĕ2qNČ[�z���?�9�1��51�&��.\����z�+��Aj��MKK+Գ�~�t�5%�0r�/�z\��*$V��w�P~�s�����=l9��1�BeU*m���Gh�Q�(�����L��]X�ib,�2�z�'�'�xt@�C���L"x�#&9(Y���h�����r``�H�"�5�v�"{9��=Zæ.���μ��8"4��$�����*e"D߇fag C$�:�Ƅ��^';6�+|�t�s�BRD[��4��y��X�Sj��D��/�4q��P����L ��׾��A��;� ߤ� GB�##�o�D2�����'M�A`){O�j��e�Uy6t��uA����̊ݦ~)�����F��eln(���3���AC�D��S��zd�H.O?��S��%$��ޜ����&L���f�2<<n��h���z���nK��!=�܀Y�����'ȝ�d��$���-U3��)�v�ԍ %8ߡ��-�إ#�F�s�Kߘh����\�OO�r��bK�����;$U��7��}� I��ׄ rTޭ�} ס�{��G��{��>}����	rttdB������DPH��z�[���$��a|ի^�T �(���Y �	��2� T=5K�l���t>���s��r%o@� ��g�������S!���f�}���!MJ�9��ϓ����W�;�C��WV�VPKB#����0ZvTi%�u*�N�"�������:��m'�ۦ	|Gh�����L�IU�ڜf�E�]5��Р"��ZH��U��w�^� G�;�&I��q�$R�A�w��?�$��W������y�y��8t���,�'W���^�Q�=v��ZΟ?��zu D8��Buy�;�����f��_�ZՓ"��@���ol��%?)5Z��LM>�-�6�$�Z��֍�.t�7��!2ݠ�����A�ԅ,�<@P��f���u#Q	byyNݸ1k$�C����Tp�#y7�Ihǋ0��(}b͉���I$BH�X�vC�r?U�B*O��=�i?J���YD��S� U��֦�Yh��1Fq�u�qh�Vy�S��"I|&�k׮���#�B~��O?=s����	�GU�P	Rϊ���捇]�jC}�[OB���O�H:���?߭�x��@��V�߱�O��QD�튓( �z/γU��l�'�`)*\���ݎK�y��yn�Y MB��
/Dy��5��6abN1a���7���y��,�8c��k�;��w}��$ݰT�Wb�$�B�0Opx>c?�f�I�3���&��H�x��9î�BVN�ur��d��`�&U;;��ީ��z�Y��UH����ݱI"q�w�y�:.�9���/W���ԏ�ȏ�]K����?�ա8T��?��X,;�J�A.�u���}A�|0������|�I	�+����_}v�v�kt
����oT����@�=�S b�H"	ϗ��Rn�'�Xe:></�?3V�)a75�q!8�F���0�����#�!8T��~�wr�CI�h�*l��-T��	2q@"������W���MǍ��9+_�ŝ�����Y3}xx��4��4tL�!E�;�I�+;� �~#��9��	>���5<���}Oд������dOO����)p�=�y����
Ө�` �Q�m��"�j�pRl��&TR}&M�'�;�(YE�_��Y'ΑN'��t��u%L�[F�j��9��d8��@��F���԰��D�/y����|llұu��z䑯�����c�B�%�6���0�KС�����
�N���
�H~XC$�`�;�߁��x��S��%ܫ���ݱ"ui���C}�T�p�bg,���{:(l'F���>'��$b7R$����� 9'�{���x��}���)Ձ8dd��n܆1x���4I~N����츁{�TWaj�0$��$I6Ex�a	Gx�E�)���_������}f		�L�N <c�p�����j������L����K�t��ʝ"=pS�����`���=���n�Z��5f<�����	���G��={���(�j՘48D��\���&�]�$��N�M� $�P�V<q>�p��^�$;e����X��X �a��R���Aag��*�����n��z�&Ŷ]X�O��կ~�_��_}[u� �Þ��F��v�	�E �N.͇&H�Xl�j��9����ձ�����X�Ԙ�����af��FK�ڌ8&Pɲc�.���U�� ��T*k:�a)�]̨bA�p6A�HվO�.�3����kmm���>�ē��'�p԰3��Ux�~3Y�[�U�k�n��M:�_��Z���-x��`Ւ�N���H��G�8W0ԣ�yzz}�?�G���m��l�G�ńHH�P�b"��.n���?�ဟ�k��"H���bA��N�� pndCe��&J����z"��{ޫ	�U�᰽X�v{ ���A��/=����Q�����9�43�0� Z�i��R��a:f�0H���S�H&Y2��y�v\����޷�옎��6�Z-��òZ^�7�=b�t�����a
�����1����*jii��'�uὒ����7-�)k>n{��=�!�a��7��J0h;L�Lj��	[ҵ�����T�E^�1�ߝ��n��Z��|���<<U$/.����D�6W0!z����=O�a_�8��p��	�����9�ժ������c��8�����Em]�-�ސX�8������ ��U{ ��v\�����z�k_�>򑏘��!����._��~�������[r��,M�yh����s J��`K(���%?����΂�Yz(��*��{ �U#]�>���DbH�p��f��M�m3���A�!���>�^����Q�=�m��nj���$7��u4\A�n���̯J��{$=��z�A	�f
z�G����s���ݎrɪQ DH���)��:)38C������$u�A֜�ƈ��	��Uý",	T�i��`�j��������=�� ��7�7�/}�o|Y���h�|�� ��gfCC^XX3}HG���p>�B�n,�&&�5z$׬>mE�Ab�*Y=���)�g�t�`AE
��U�v �3թ��פ���t�����g��f���{��]1���~Ь�d�^��B�I<Pt����AZ[[x()��tŚ������Z�}�ZyG�RG��ً;�8��#qG�$�J����֍D�Ar<1�ӓ���Z�-5��VV�M6/�@Rqh��J&��4��߷+v��$��ߐ�Bx�q�]�S�� ��R��,敯��_��O|�!�!8l	r��F�J���R\�&Ȫ�L�@v��z��^f�x��1w�V�S�!����U�Z��x��$ft J��s(��^QY�����?{j:eLX87���n�(Q���_q��sL���bqӨ�H=�w7Uq	k��ʴ������o���yj�~��'ٓ����fb	������Ï�M�	��%��щI ��#E%�&��˗MML6���{ �>H�k�Y��5äI�#��RTǑΓ��OM����<�h<�$�����%����K~�ᣕ�v�C#���h��H�G�!ﴌ�)M���)�8�� i5I�����/0i�fg�|�B�q��e�v��D	��B��J%q6�䆀f ��u�� ��N�5�Y`���X�쭧��	��Q
�a�\0v�qL�E�jK��"�k���<�=���������6�c��9�7�jK��*�I��0I�=� ���6�a�5���̻^\\r�� A�+�V�'��0)8��q܁�6�`�G���9"��s���*d��cO\��߫�=/���~Z�ſ�: �F���Ϩ} /
v�7)B���C��iH�A�h0 e��իWM� �����Ը��;s��[)�
�L�#Ui���8��$b}�8��ɶAz�F�'$� +��'�A!|Fx���ss�����I����A�m��bd����گIc��6�>��e��+�T<0����O�c&g<����4)Bf-H���6dԚ�����N���� ���DoO�y3���  ��$J$E*�
���,[�Z�kk�����A��'����d�\���O(*��"E�������s�w�s�ԽU]��3�=�P���tuuOuuս�?��/�>�� ��.�B����XN$��Y4��@�ښ�S��w���7�zZ�a��۷������N�81�.3Ribű��2��~�:z�eu��99r��R���J�$�<ƀ;u�4}�9����Dfbm2�W 	�sqq�[?�(�'C���/U�ƚGF��H7.��j5���܉k����A�\�;��s�[��� �'Y��{��AD��?�Ke%�����N�~�h9�	6�"R�6'0F��q�O|~�#����ͬ��瞭Z��M� E47�"45�vDƲ���`��B���T�Ȅ
E�J�\���_�B
L���	A9��|^����rDv�q��ҹ�[���7��&�O�ˌd4K���+u e��z�u睷��o���Q�E
:S�F���E5a!m!`����"�ɧ�Ѭ^��U��N�6�����F�8��u&�4}Nj�"�_:��3�I���n�E�5e�d��юl	B�P��#���T�D�Bp~��X��-e���3�;h�.FN!��Ȍ�ix���jz���*�1��ߏw�k�]�SN���KĘ�0	c�ؾ��%DAp@�A"�����V�B�s�N"���ϻ�	@�nmm��|��^GDm��2�N�<I�.�9Q';XG�CSS���6AB�_)Ab"��r�b�:w�V��Y����Ao��rl(��>L��P��#M廃���7	�*�^|�>7 �:�Ҋ��[q�+W�PfͤJ;ŗ���r}��Ct],j����`�^|��|�&�7�P)�*���ƨK^_��&g�����o;36Dۓ���~�<����s�X��D����K��[0Z!^�\J�q�G�@@ ���R��Ƀ#l����0��;�{A$	��q0��(�Q�	y���!��@X@V���mӪW�����[�����?�.#R�AJ�E/0���^"m	6vh������ַ�E����tA����IJ{饗��=G��;v&1��<?$��O��׼��F+R>����'�da��F��:~�LG[�qR��mFU
n�����@j(��%6�EH�o�k�7e��s��{$�'����"���7�qoil3�D��j �|ǰ��2�5�/J�R��;�2w�UnVr^K1�JG|?�"a݂2�f�B������B�Qk�s��b	�G��m\�o��4Aަ.#R�LY�8�fg3)��mo{]����Qaߣ�>J7j{:�r\���w�M���M����MG0�����Q�gb~�������i$0� �	�� K	���sZ}e:��d���1)boRn`%B	��o4�^0Y��%�XM2�v�}!���oh�I�ݢ��p'�VTRR���b�k2��B<�i2��b�I��
B� m�;)hJbZb2�w�v�fc�1�I��j��m�����7��-o���㏟T�	�$Ȕʞ����#Z"iQ���i0C2���[)\�.�/�v0�0���&W8�����9��PkH���5>��Ѯk��ߋ�l|����80�Td��A�]$eL��p��d��v�u<ha�E���Ԣ����f��Ն�JC���c�6����B�q�J�L
�	L�H#)v"�K�*;t$+�4��%����>+ rǹ��Pe�
b��s����\h�H�I�-�UzT��:��N��ccM����Gon����vzz����~+���0��f��Up��Q���9�t@Z�l��H9���}zp!��̉�ei�Ń;5����*�g#���>�4�yH}���ټ$�-&\�`��^��)!�,�;�b���s_���H}X|\;v�rMa1AoH	��� !۶ҰL�	>��p5K�Ń��BI@T(�� v��PGL��Z�Bv�/"&]h�PT�/���������k���>��_�˄Tj�шq���`�bQ�I�Kuuu��[h�Hs�j 1m߾����?�<��(��˩_�e����lQ�x��)qQd����`�e
�,��������eq�w v>�H�#&��ɒk�j��F�&�9`#��Î�����!���2���H�{BJ�e��<̡�i�e�Y.B.�_/��_��U����b�3H�p����)�S*�I#����s#g�C��Y�&G�&[�l�~��W�;v�ث�2 e��*�����̣Nؑ��B8��HQ�O�V/��"�^���q-��� K9&��H��Ԩ7҄d���,97,6W1yrLdV5��A&�#�&� ������L�<C��T�aӪе�۝�]�µ1!ZJ���&9��&�O޶[��r֩8�fҽn��xFc�yy�n�
ȃM���i��/�n������!I���`W�9K9:<����7��B�6��(
�FvZZ��k"H{�JD�r=n��Əh����H��!)E�"F����/<OE�aB�8L*������~�3��0��Bځ��M��#������ҥKZ� l��xU�GeX~�X��C����	<�N�,q#�]�y r�YY��di[�r����w��xm��҉D�fA��B|�^D]���m,�ׂ[a����[��cΌk��Q���3y<JڒR�Bj��Iu)�SH2(�%��IE�������@3C�+\7�V�t��n͗�
�(8��H��[H�����"���_������������Hz��A�"��ZP)'H���R��ݪ��ǕZ {��BD#P�$�C��O�M�F�hX6�ז:�yq�[	����
%�z0��`��v�]����Im�%������-8��"�6E����-�QNZ_&�(�����6��4�,�jC�^�b��g1���<�f����F�noI�O�#��,L�,xe��]]]EA%R�N3A����h�D�8�-�$�
�8�|���`���wd�E&T�!�O4��E����, H��w�q�w�}[�)�����Z�hЊ��_|�e��H��u>��7>>Ii��I�?��H/�$o��6r(��	��7��M�*�t���̸!�ˁ}~ &?�/8�1p>�U�4;:��3ң��%�U��I�e�e�=,F���ԯZ)�xd;��\3�H�ޔ�� >W֔M���W�\��Y�S���G|��f9��C
��)n�}O�WQQ��(�GƬmy����@����j�&'�����严_r�Md:�kA"Ђ�Ǔ��"f݋ ��[��J#�ʶ:aM:v�	�8'�WH���-9&K����V�} Ə֤e]�Ƽ�QiT�����$�V�/O&���T&=� A���~@�C#YB�� M�֖� �a��� &&T�YBjC� "bq�C@�z��Z��E&R^��%��`Mp��뷫�_�T\x��B����������Ik;h���t8��h���~�KEE�[N�G 2ciP��WLpA�1ϙZ���im����#��L<�ha܍g��D�9x`�@`��D�b26))�1�ʽp> j��s�螋B�F7�l2�+��b���C�qϭ������2 �9�<R�$hE]]}df�M�o�M)j��v��&�)�m1�Bۃ�d�J��%�����[J$��	�.��>::NZ"4���z���>C#}�Hp�w��GuUQ�fũ)��PS^�5���{��_k�mc�L̤~){)"E?�d���oܥ��j�#�i�!�A;�)H�9�,,`��a���;�s�p�'bmAb�����=�u�-��TM��?�{�o�i��~�>�=Z��kii�R��T�X���Qi�RVV�t /���=�3{�� %:t��a~��
-�G��ɭĶ	P�c��7yM� *4Y@��x���˒x�|� ̼�W��^�hH�+7�E�j�������M��U���Q@�)�ł8��&�/|�$�7��%B2�~K\K���F�|̚b�K��)qxk�/�C<�2���a�,;6A�&
RD�L� m�Oss3�bH����-ǧ���h�����y'�����B��.=ߎ�UD�R�K���6��%�b[[$�7�0m~	>�k�30����I��5#m��I �?DĂ\��S*�?[��ƪuuu2������=}���h���ĉ<Lȶ/2��`�_W��-�58�M�d����"3���������]^��$��[�%�Hr/A� B�
��.���޾};i�n�1�o���e6�'���)�t*���	b�x�ͧxƘ�s�ͨAڡ�S�	��D���{1���q��\�	LOONBˋ킞��啪S�^����!�F|9��_����@��"|( �Dh�H� 9ap@�M�i���j��ߏȹ_ytn N�"a�A`@���:��qDk�m��3�ڪ KhBB�r|o�H��`��E��7���f����jvv@_�9�`��B3RR�哤I+�׶�D�9�gXp��&���V0�!$C3�k���t؈����v��~A�G�)����7 ��x�9s�Zw����*�gb�5�".x�$kR�e�rm��r�~��ZE�� �E�Z�Y(Y`�����ېҽ9�~i���?�1E�~����͇d�L��@����)�'?�	}D��/�d�rG�G�J��� Dh� s@&:��_$������D{��q"K�+j���VP�e>��W�>|��E=�u��Eu��*.��������s��� �]^�t��ҡ�=-2Aډ�_
���o�4-lc��(p?D �y}�z����-��!率�Lq�x�D��C�����a��Z%8�\̥��5��McӮ=kr���E��a�y�o���B��)��� �#�B�h�r�]C; �{��v�ܙ�êE{�� gf&�egТ��&���
dٵk��9��4��56�ϞL�ф~��M$ ?h� n�H��4E4�dq�1(`���,�[M׭���.wdpww�	����	Np���4�����=���V�������;$�c,O!�b��<�u�A��i��?B2�fYj�o���M?C�k#}��L��Bc:�t@P�%-�2�O�N[���垐��(XK����W�Ɨ��eڬ�E�Z��	�S1ߪ�0)E_s�M���&��	�9�����6���v��I��J��Rm�Xg����p��BlC�������6Q�甘���![��bwZM������;�d��|�F��QK*7N���|�E�z,v��>�K\�U��j�]��1^��+���Cm��4�O����t9�{+[\��﬐��V���ˑ{0��
�G�Y�X�.�,�'�G>���>}r�}�Ǭ�(Z$���N����/)�W��p���Q���3����T�6��PD�K�!��S���Q<	wu�$��_/Y�l��:�<J��	b\ʆ���/<�Eg��?ɶ77��8ɕ��X�t��tw���RI �T���!�I���E�q؍Ġ� �v��+��8or��<���f�s��5[�PT��XУ&�"
&�>�^���!����Ў�%��	s��z�א��ٿ�,�x��t#7�$+�u@0�Y���<���s�/�#����p\ė������n���r��I>�u��������ca��f�-�w@p2���"[h�����#"i~�g��!����$(��8>��-Kq1��ccY���MMr'��̓�5\�+�1�q��qc3�9�(#�:b6gf]&'`wo���$~�!��!S���0~z��n%����P��I	i)x���W�˂�Z�O��>#����O���%<չ6,H�D	�}(��akl�k2����0�l�S�6a]��0L?Rj���b*C�(<5�ٶ��g���H�
��o>MzO]�����j�.b��ʢ�;-�s�6f���N�r��L	�=�L-ޅ�C{����x��\�0�����V_�r�����U:fn�dk���H��T�|�y0�;5�İ���*h�"�D����P��YTׁ ��$q�t��Kl<�n��G��Wm�9�Wl�I�MV2�����qu��G�KP�g�%�,EIIACz�@��Q�Я	�&�1U�<]%j��V [+[寀�X47�*��*(��q���͕�q`K+�����b���Ka"���?�������c����_���~�#G�4(�Px}�A\��ߴ�!T���J��&��+����y7�1��d ╨��8J<1@Ȝ�o���9�8��qo�@�]���)9���p٢@���9E�5���O`ż"�\NP,�`����n��U���MZ�5�eݹZo=%x��o�8�_W�|�Ĭ?Z���d��+Z Ԏ��\�9�m������ag�N�;~�\u�'$\z��>J5}"���,є�SZ���x>qpƔ*�B&��觟����m�<W$�qZ�u�$��m���<Y�� 7�xI�(:^nn�Z�؊v�1�k&F������<{���@�j�u��0�0�c�g/6�Ә�f�G�se^���P�^��ݵC�RH��/��D�\���H7�
��Z��6s1s�'��_��xٴ��83�Է'�#�%�
�6(V9�����ƚ�ڠ��{���~>�O��ۡ����h�mvU����S.֔��e
b������0+~�ފ;�s��vߜ({_;�_I�}��-�U�~ޖ�(��_e�[��_��/�sʹ��+M�93�
�������R��S�,�����>8"t�/��P��e�Q��6��89��ṖW�H���p�#��2��nw��.�`�d?���dt/�f�ɽ��A|+�'���0���!��"r8S��| o�lN�' ������ؼ03�)X���e�Z���Lg�>����
u5:�63� %��6ط���ga�C
��Ckb$��E�n�p},2y�(����\�x���'���S,H�o�pL�8&�c�@�Y�.���]�-F4 ��q���L\��C[��Z����5�R�&�������cTCe�����V��!)�J�t)��t��lʂ�A������9)�X���<����F�[�w{� �u��F��hv��̃� 8WןӼ�\��|�H�::�:�����!�i˯��V|]����/��p�#��
���_���[�%Z��3�Bͦ�h7s�5b��/>[q�kc�Q\�-��"Iz ��X���=nݴ���F��3�Y7g�Te'K�����R#�1�^?8g�X��NA�8�L��M���ZS����ⴑǝ��?s������P���^D�¿�Z_�:l?Ԇ��}˞���3��*���\}_�e¢�ǵKijj�\
o4�V�4R�CG�\m���L��R�	Tj��^sM9�S8�چ]B|��!/����Lk�ާ�҅}D��N6
p�._NVW��v��sq9�ŒIrR��b�!Q��I(|�k�ց�(l*���=Nc�K��̜vرKxs��x���39M�+�7�2Ȝ�qt!�cC6�q_O��ߤ.��f�(��+_`[���@��O5�9�\F���e�~W�{m8F������^}dO_"��)��o� ���h�w��&Y��g��]�9t9��J�L?�����|�R���m�!�����ng�'��[�ۊ�K���D�}Z�Es��߽�Rn��ƣ 2�Dߏt�������+�PJ��%;�Lbg��Ƭ/WK�g����}���}��I1���h�2�R�>l'���q�U�Z�w�vQbj\�J���}-W�K��)�fOk�N���n���R�z{�&+�=ކhR�?J���0��釾�8>b:_I��[FE{� (x���a�T{��H3�Y�(̱����!9|�(����	ް���q@�]`�Z��ڿ`G�mZ�a&�W/8!��f�~?��ƍ'o�i`J�ԿyE��8����?%���w�E�v�5���0�ָ�y���s	17�s����M
��o1|�-�_V�㣥�w�?J��p�o��V��.��:!+�\��m��)��D������fycC�+��
��l>0eQT����ܾ�K��xD���a�l�>�t�κG�W�N���(}�Kq�"p�./t��.}�>>����B2��`w�O��}ϝ�_u����h#v� �#o'��6�'w���ػ��lJpt/Ӊ<��_����
�o�Q%OD��k���+
C��^���`�m�u>/�oi$��mSJ_𸯻/%�!���s��/��;�F�	G_�K	8�� ;sw���!ih$id{ &���b�l̃��w�G)�"[�1:;��"EXK�u�$������sN	���T��y�Q��\�e(uI&���S�&Ч�f]ۖ&"� �+��x����1d/���o!��L��"H{a�Y�[Vu�C,��E]�z�ޅF)��	.���2�i� $���
�f!br5��s�-)s(�;e��*(�cKߩ5�If'�kI����K�ڠ)�x����)=S���g�Õ�����m�F9�c�����@ȯ�ƪXO�t���k�P�fR��O7�љwj�.l�׃I�4�t���V-�^X=dǂI4�0���V-ůQI�߰�������F��8�����Z���J?��pH��wY�	���K�ć�*'�(5�f�r�Qҗ�?�"Y���顚��b��_d</q�+ Dq��Z��m �1�SZ�o43�p�W(SJ�.~�0�ȸ�rAb�)4��9�+����,�&sv�E��3�2�t@�;y����!,��Զ�fȣ��(~��2(��_4�4KJ�2��c-Ѓ��7vDG�:up�{�˯����1��̞76��E
ē���b×�$�ݫ��!�,�)�)3TE���8Sd�^�L��C���j�9E��M�K?�2��?�L��e4?i<G`K�K׽x4.��X7��N�U�!(U|zd�g��^}ʎ��'�yؙ��x�:3+k�:��q���Fh�A��3��ʒ�+�$I�[U�@�����a�����T�Λ�����d�����Pȴ�ق����G�詽6ѥn���03�\�*(D��Ü�Njh�0o��G��������	��%�+��N(i��D�4�������,���z�:H��N&5�?��hnoŗc
�6t��Dpt��R���U>#3�Ô���q������}�z�4��(I��4BC"��k���S4�&���pF���ȱ-�o��Dx��M~��K�	�R)���|�*�y4�=	cC�{}���]�?�k��˩q�U�X�W���p0�C���E�&m��c����x��M�Mg|���0L�W�8u�,�ݤ�O�6��D��<�o�����V�[�v��u��7�hl&�l%��(��Y<Wl�J����t?_o�k:�<Ln��EŬ�d:ae�N�L7N�G��0bm$�J���C�H_gG��n4��R��"=�dx��*M�eP���m��
�� 1a�p@79��>���n�*J�U>�U�YYZ�����>��V�} �}�b�wqs���HH��}(lۉ5.Y���Y�����J�������u)[���M)��,@b���)�Y "<�b�tG�þa����ά��J�"�X,� Ϯ�	�
w��|c3c�ݳF����Y ��dX(����	*���������<S����1����~�\�r���L~	�J8l�c�x�}�;�ϔ'Ka�w�����P�f�g`215~O��w����"O��a������X�2 65DƢ��Dp�܄)&��ڪ[��^��S����jVA���_U��b�'!\})�\�K<�hޝ�8�������<F�3}���n���J�C�n�iv|*�����"�KYa��GZ(�Z�&bc���f*��}bws�43�����"�������^�����nt7���̰�Z���@��f�[b(�{k�-��"xi�>��`CA�y�;S]��A�U�FN	�Ґͬo7�/No��/�����{���}�u�?�!Ĝ[P��e��xH�~\5��#>�'�\������A�!v��C'��N7�Ճ��BHlal|abjz�{p`p��Uǈ�L�0S�)-���r�PA&x��T�Q,��ݚ�XSm�/s{�_�z��E�z��ZS��w�D��79V�4;���Gj��!��/�?��)�C��3�~�Z�z�ɡ`9#�����u�i�s�Ӆ����=�Tz�:Ie`v�8����K�>�h���x�L���=��@��w)���� ���6SWշf�(���_lfp-Ԛ����o~��D|$�	�o�z?��څ5�ƁǗ��E~�7��-G�D0u@�IC��$��j�'��<�L�S��T�L�$���r�]y� �ᇋ��i8u=)5��1+������1$��!����X+��QĄ��n�8��|^���hH��~0%%:WTңh������H�Ơ�=x��'��n�3FE[�'fDRg���X�"G�jdu*dj�(�@�s��R�/���ڐ?!%e�6�ˌ�m����q�G��`.� ��Ե99�?]��s�� I��~��&r�俇��O�4�\���T *	AEƌ��	4�\�s�*n9�R��K��ݝ>�7$b��c�d>�i��;�
�x		�`//�ܱ����G�����v	���
����ׯ<�6J(��sr��g�*j�T��
�^��:�ߜer�d_+����U`�"=�k���H9���Xp�	��З�YFn�����㹢��3�1ѷ)[ۻE���o�$%`%Btp~��ú�����¼�7�u��h�<@��rw���I�~*0K]�N!�O��.
rў�O�~&�v�j�m�@*����׷58��PxLV,,�Z1�ZgQ���t�(�"� �K�������;t]f����3�NZ�yx[�<n���wpP�~�5����d�aZ�y7��ܾȎ�Or�Cg��+�b�&4�յ�iugި�|ĥ�"���D���#2�1S�JR�s�jQ��8��}��ò0�]V��j~NP����2-��x���A��ys�/`����O�K9���oN?������p�%L��A'���0}�=���Ww��Ƨ�e�M��e��E%����?
�4�͚�~�I�*�w<w��kb@��e�j���y����Az�pv�����)�<~�P>[�,
#6/H}"������"ax=;=][*�(����pp����;��"��ť�P�+�_C��0n�}��#��#��	�B*:ofn�����>��;#��	g��fS;�X(Z�2>>��KXME%1������C7 M����Ƌ�^��z��}���T��GB׸�x�]��&�̇��^�x�����e ݚ����:�G�Ih����%��е�XO���M���%Wmز�?;.�����*�䖎#W��{���ր"E��R��û!_�c�ũV8���8ɶ`R�|�S�,h�`ܪ��SU��5𶖔\'o��ˠ#r��C��K��[QQp��q��r���}��P�6�����얨��O."���k~q��{��B����λ$�{��j%����Q˳�DkѶg�Fb-�o��٪G��Fw��������t̓mbv���Av6iU`W��si0��F���+�D%��V�
����ta���h�kJ
�fl�0&"⾘�ms����r-�������ۢs�R�;]��6t+u����oSB7�m�w����!06_��_/x��΢��N����Ǧ� &%�ML�)i@�����J��-��Τ�l�UsR�ї�a=�֊1���=�N�u��_hOL�J�����)F;@��������j�Ѕ����E��3i�0��#��e���+#����ł�p�� ��}W�]GSK�meG��Y��r�=������ႊ�A��ddg֠����C�å|��zZe��V������oc_)1����1�C9b�g�8��{_�P�Ł^w��sߌ��o ���Qmr��!�Cw�/�z0`�̝�_F�+K]��d�F�8pH���NN�<U�Z��D�j%B��@q}�A|��.��W
�[hͥi�"��i~~~|��^1,��r��a1|�6������oo���Ŵ$Ə?LMGe�G��C���W7�zn#S@�@�~Ǭ`R	p#W!	�:�u�tbo��uɫ�(.,\����\���t�C"��߆�-8�[*���c`N㏥ZD5��_^X�ږ7~�������d0y�������g���/��7��8]O��ƌ���¤eb�����!%?��)�>�&8�5��2�ot���q��[���{Uan�����O�b�CĢ���p����I>N��}�x���4��(�{����QRL���]�W[�R��g}���G�f{�6�KJ����ȃ���Io���V�+��E�E1���b�ǬG�"���Y7��.l�UL	V	F��0WR�>>>�s?]��~=C����~����������m&-&v�%ۦ&����3s����Si!$��	�<o�w?��v\�>(��;�U�V��}L�����G��gd�j�������~YP�)��栖�v`R����G���Gp���
��N��C�|������,���Ί84ӫ�~m��υ	2[���ᕝ4O���Xa~�r�C����͂�,����W�����[�<
u��)���2����Z������V���U���QR7���������ό���x���[[��d��1<?h�������q$,�(4l�_R�y*q�$B��׾8���a��VT����]��!�/~c��>Q35U�,I��aia�;9�0���"'7Z������z���o�|1_���߭���]�b�s�=������C�OG��ַ�9����_����7��]D�\+I��d����É�:�ML����[~ee��b��_�:C�G��PZ}J"�U�qD�qu�F!1Ie��L2���j�1��@�'"3�x��چTς������:@o�So�L^w7H����l�����Y�U/�l�c⎈(!�z�عU�.���^���;t55�U$�N��q¢������-(��X�ӊ�����E��_|���!#��I�4�t�B��-;sQ� {h��i]��{���������߿���lOUC���'-Z�=ܵ`�1S�Q�,4�,���Bı�y��?9�^�����sC�C_k:��x�yPŞg6��d o�qU�5�c��vW�}��B޷�%5"n��7����b�rsT<�yh`B=5q�m����E��bRRGG檝skc���{ǫ���X���l҇]s��}7Gp9m�[���O+����:��RW0N?U��1���`�1ۤX�Φ/�+ÒhhIz~�/���(�8R�-�*��ʑ�鸮��׈��J�L&��9���oۻ��1��1��ws���~R�>gvܪ���@q �S�o�سT8[a�h�/_F�xxx
�rE���or�����G��sHs[H�p��}���z���OH�-}}�޶	 *��#��X2������g)MMMyI��� �Zv�Z�x*1'� �- P��&\����4��$��zb6�ʀ�"b��9 ?��Ikk�1	!��\(���VF���ΐ�����m��e��]9��P�ʊ�:<|Jy]��E��A��1�򈚇N e�3�x�{��&ёn��6qy�[��6_d���Ɔ��������6
����~�h|� �Nt�E�2�~3u���S��E�k�iQ"���Դ4��Ჲ���n�vNNqB._5?RyU��fad��Ə���*��T�a:�~��h.�^���}��[��!�p��7S ňgR O��K�lT򋾱���VG�WcQQ�\�����G�X��*��m:E;xo(��XŻDt���lRSR*ff��sr����|0nGyy�b�S{��=+<<���Q�	mSpc8e{W/��x�S3��Ц����M��νbq��S��ӧ��GB,cW�$���#U��8�7!$�~���2� ��72A�Oʻ������E6]`�5���kK&��oOeH�"K\�������e���
�����ZZ^a�)&� (�xƑ�"a��{@�K�,s���]�P�xw����&���hasS^��|ix�ttbB�T��xi�)�ͩ��Ǻ�W��:�"�C-���OYc���%�E޺�"�-����[������i�q�ZMq'���9(�Tq1�&0	��q������AKp=D�"=
���\7���(i�����/V�d�6%�lOLFF6���L���Xn��������b*�V���Cr�pǞ-��I��C�.��N�h�)��uI������:Ϛ<Xy}�, VBB��7T����42R��f��5T�no�!U2�	�V�����4�'�n�D��JŠ��%�;��>ኤ���p�Eoo�ű����q��DqE	C�KĐG00�T:�bc��W���0��cf!� -��W�ð:=;�)��~�֩��R�+f~����&���+L5\P����,�F�Ʒ��,m?R߶)%v��  �2�t���j�2W��z�������_Nř>�?OG9U�#�V��$�.~C�ںȰ=�[)�Y2��4��!�C*6aC-�I�O�u��I�h���h�Ħ��J�`1�(����=���R/�۶��S�@���&8dyIAA�W����r�C�7.ڤ�L3!�YǊ3k��K�[6����XBO�wI���J���c�o+vT����6PWz�>��>A[CCa(���gժ'c�v>��lG\������A�#	:�#`t��� nX����[j_�;H���X�m��������{��f��|�z��BI=������o ���y���8o��@�1��k)9�\�Ia 7;xX�a�u��K���x����b_�X��T{��f��/�����k�0� .���u�ܘ\��{��N��B���Cy�S�pH Z�y�H�I#s�
�./U���K4���d�'���~蠞��8�M�'��~fv����=��	u�cٺ��>��$O۞_�����:�fӿA�~%9��y��~�Z �|�r��Fh����H1ٰ�q����� ����
�"|z��9h���=N���?�%�#�c���!������)Vo/_�R��@�`�h�KJix�Rk�/,V�k���$6pKA�7}��X����o���VVڔ?�~��I��6���O���`N�%�,,,p-��e���4`��#*��9���ut�r������D&�5'㑨�W�"z�cC�gfz���I�HO�^���y�Zy�
N�8{�$�V�^T;pQ��\9���x�(���ߙ��+��� (�]����8���]e?���;�(%q��!/��9Iq"f��������'���!�7�1�4[ʶ0b�>3��C����B!
����~�����nV��Me]���ߺ����A�~� �|���k��ƒdh�~"���!�3��F�c�����=(yy/҂�E1��͛;�"�
�����1ix�e\]�m�""��Z�t<e�0��F[�B�؄�e���Iވ���W~���\����'pb_���)^�ҹT}��]�c��jK>�BU"l�q�WX�XJ:|�sJ(v{�ư�;Qϛ�ߝ�W���B�����D�U��M�L��p��!�݊z�qv���r��f��wێC]i�B����e��+k��~���~�e�b�v��\U�)g�	���f��v9��نPul�,-)�轢?Ң����������򝅭�7M�Td�-��{�e�B��]���#*uk��0����� %v�FF�b�@©5�v�"IoZ}�O
��X��en�Q�ǳ"z��DN���P��	�R�A����7��P�9g_�qED !�񯇶v�@���쬜 �n���gV�Y���;�	BD�L�ɾ��f��es�9^����_M0��e���6��Y��ݏ�ԅ��uH��@� ���`��|�b���v��~�J�2����
��^i�,��<��O,�W�U&E�/�����
����`�i���P��)>��-�� 7w�E��]���#R�[��Wj`W��H�監�]�������#��=�~��~��8^����e,�a�A�l|Y��yu
M�D)�x��?$+u�c~��O�����Q�����ٽ�P�#���?�/%֊_����e�5���Oɛ(�*����!&^�;2���L�:J���΁�U=�߇�T�O����%�@9� �+rg���d��s��W!#�s��C�9��E��tO��ܭ-h��]��SOO{���m^��ʆ)�z��ͱ�^��(�;�vo��u�-������_��Vͅ�P�4����?�Q�pE=S���C�	;z���b�	.u����>^���˻��&������!�V���,�(}��z0G�1/y�����:7wR�)�@�P]UԸ2�,���L���u�<\?.� �ص��x�c*G��	�����hko��_\|w��X�h1<L^�J�/�6n߽�����*���뛎`�^�$w�ݢa�?C���'J������5���&�r��u����U��H8}U�@ʓ�������GT��ٞ�t��ғ��X�rY3�HؕT�]��Uo����~�Q��p*y������.y��)Gl������1l`�&ai�ν�((XL��-��A�.O#�����V檒7���n�J�u;NH����I?�m�4Lm�d�y�Nn(�@�*������\�
X���т��Ș�yܽXR�����;�5��I�s���M>߯�L��q;��R1��Et81v����l&.�Zh��Y.1533/������P�rL��b�><>����:?����x�������n'���?vt3)�]�."��@<�Ԫ���1���215��dafk�87H
a}S�;7�Yk<a��?�>���I��Z7���r��S�4��Y��0[ćT#~���˞�T�����������P�T�t'2p	K��i���X�"@︺�� ~ ;�b���~��LW�uƷs/�`�S�L�ga��%���Q��^Q�hx���E�^t6�3��j���#[�?����	���o^���2���-�-�-ڞ�����O�t�
�j(�"��d���<Ѡ͇bɀ���r
Oao�&Nn�ۣX��Z�RC�)w�
oZ���x���}��m�xcM�
��+3'��t��r�%�Kꅏ|J��g*����8URV��5�'���8�`վQ�p,�����8��� ���]��]z�G#R�Q;����i�AR�$�FR~Aʭ'�Y��Pg��=���q=�e��.��)mu�F�O��Ղ�$Yl���D���f���3+�����!�U"|��\G��n�|\��շ�1]�����4L��i_�p�����f��}���9�ՉL?�\�����dff�+]�oW�d��\^^�1�Gbb[�4��]T��t���fgf~`�2��]��*��E�f��j/"�Be�\�.p��e��7�%������}�x:Z+��z��ݧ��;|e��D�V���8Bw�����1�P61�zp�Dl��7����i=��8'لȒ����]]�d,s����V@�J������{�D�(#�a��_�#<plGf��ǔ�h�=5_��x��0�5Fģ���f撲	�T/R��3I���*<c~��6ُ���fn��r���$($���~陘.�'oճ:��υ\*�ۅd��W�35�΁+GŊ�.�Ls=��PC.�Wt�}5(���ѡ�.�?QK�r�f+F�.pH�u�
�oJ�n��2	�z����@�Q�˩���/2E�U��sO���L��6 �1�� ��B�܃���XfZ�"I�/����QS�N�����}IUu��N�A���g����UA;d�Ș�����胉<�VW2�4������V*)1{�#��c�h�-i�s�t��@�]�iՂ֒���&�VRU�b�YxZ�Ya]DH#B5���z�vT�'"r��C�OQUH���
�M��W����ڰ��q�"y��_�|��3�i[T��g���I����'�p�u@��%����ǏJ|G���I�������dy�x�zLG����^��<uRP���MM7r�8��Yy]�kk��`@��UQy�~����KU��7Q�������R�9̴ڬ���V;�Io~2j��p���+���\_妩�dP��K��3!UUU�z�:�<��i��i��G1����
Zv.��,�h+oCq`j�����R<D�ZvvCI!V�GPl����(ZS�݈w��:U�$��*����Q�op�v��9p@������+���4�C����Ix��oA���v�.�T�����.�ǵ���Ȏ���yh�#����jh��[��^ebN#�~~��u����㒰왍�e�㏁S�<���j;�6�q~����w��l� �����>�E�f����Cn�o��>��:8$����`�)��W����]��ٙ�BIm��7�;��j�a�vg��)�3�ү���R�g9�D��U[���5�m�����k�%**`%������)�b8�tP�ǗƓ�:�z쩪�z^tb�{D��L���T
��s�ヷwExbB�"��Zv���F�Q���${�v�yIQ��ϛK��Y�!ʝ)�	���HŚ�mlsoC����-T�0Zà�\F�G>������*��\��fS4�I.HF��3^iWp�I����m�� 4��=�X�8?O8)R�tNd�R�e�� ]�{�����#�Å�S7�c�.\�tW��:#��5SP�d-�1�
�,�w�|dQ�u^[��X��gSRd��q��k��FKTY��<1G ��C���qM���Ąr[���%|/S���E�z7;;k�m�x�jjj���̃U14|�R�}8�գl�|���	4��a�iIVr	�|�,q{R]�>�m��[�&;w(��'z��Q8�W�F�%�t�4k/3�Ύ�l;���R���)�>u�sØ��ҧ?Bܰ]g�}s��d�H��<(q����q�~���!��xn"B$<9��@�eQzD;���&�w��1s�FxU���BJX7i�Ay�¤�>T�,Gu8�8�Z�o#p�n�G�B���5��^�;��R����o\��=��!)-=d\�,%r�(+�	@�(@�r��_�tp���^m{��𙨨�t�`�s��p�ά�kE��/l�T{lcYmm�*
�@�
ћ���"#Y�2mF��ALJsw��J��\�W��ϙ�-(������������Z�_$)eB��l�7R0Vל�Uel�I�M������Qw�z�t-���yц�k�~¯�f�[��_�xX�|�he)U]�+�0m�����0�=�Ӆ	]�x��>�E����${��%'ԏf!m���i}����m����Y%�R�Ƞ蹾~V��f&��t��������d����Ie
Z��1u�ڟ������RS�#�d�kEa��@Acla��W�w��vXa����b�3Q����M�ww��(~�܆��C�!P��͆v�=��`@(��g{>�{��U���C �pwia"��k6>�,<3_�O����C����� ��{m�����B�?5�1M����g ��U������nR�p����_MNU�kRѼTC���1U5%=�3���Y��oԳi�����pŃ��6g�OY_�z�V=Gֻjy�C��h�cYicR�q�� r���9� |��

&&��2�s��mmt���/Py}|V�
��
�554J���C�օ9����z7�X8�,[Pݩ#�3�_����R\%9�i���s�t9�ׅ�)�%����jf��C������4=1��7�2+&�h�H�o��i�/�b!������^��Sm*��A9|�������V0ˆ
!���2��IЌ���Lb��T~���7x#���긭���t�FE��D112�p�wM��m��������ۇ�|BB�"�C6�X���S��A�bt���he��=�Ǌa u�결�@���/h%Z�i��B�0D�m��dannE[U�W3'WU/~cW6R�!�X!̏([�����Qk���z&O��e{,+���7����U���My�'���r�߫����L�	�d�#������� �g����5jb�s��(�w�g��[������6�?#8ĉ��V愰L��p��ּ��G�rT>�C�$�#����`}x���io�x�ciճ����D]��g�b_f?�[B'V�1G���֜�F�PF�EHd�|P��",��wEs�ҭh����ݰr��փ3y����9�Ӥ��dM �1�!�[\�"~¡�O��<���|V7�ɾ갨;�"�e��-�ï��X��1"�7������;$*rԦ�C����S��GsŒ��"
yA��'T�wJ��06
d��R�t-:�*�����B�,و��ĸ�Co�
c}��Ċ�~�~�~����GF�$A������eC
�?�Ĝ���,r�^^U�����U�`�Q��p��e��ў�~�A��Ng�U��'r��r2oQf�25�Û�Ĩ}��	�;�&��
1̻��ؐ�0k���(/�UCV�����Aǒ��;��XM�.:�]Y`�*���J� �.��k���0��q���k�Re3v%3�=5\�c�_��5H/��i�?���'�h�S�g�Ág�&�Z�q?ݾz�e�����~�˚o�b̛�?q�/� ъaW�h��7�xgu�m3u�"r�;=oA�����a��.���K�D���m��@򿼼��P��&�Vh���+F:���No�G |��p1uu.Q��0��
�@����l�	H��ű(!!!ђ��:M��P�}�	*���P�b�d������������,�%o]��}
��n�6���Տ��t#b���+����)���&?�ukK
{�
5���p� �iO�>�C�F_5[�
��I��1q��S~��;A'1�aHX�Z���� ���t{����-�C��z��薌m��h?���fU p���n�?�t�,�����j�/=׹(��p��ͭ,�!�YZ�l�����|��`.�����Z�y*���<Ξ�S�������I����W$.N�N�n��u�o�l�l�}�!6Y&ŠC5�_E�#^A�Q������ڥ���� z'�c�K�2��&$�Mt�)_�ۼ���N�������Y 6�.˾]��u"q�&!jo����{P�ey ��ek`�+\��m۶�۶��fO��ĶӤ���n�ƶ^�}w���k֚���O9��֦-�εB�I�s2)6I�z�6.,��O����?q7Ϣ"�W,/+3x%��׷��ͬ\���6���r��a�\I��(�S�g��4�(�F%�c��! ��zۭ�ͳ��@��q���i�e�ců-
�c�"������~�������nK+A��[����t�V,��:���m��m5�ҭ�@M�[P) �1[H�X�.�X��F�&3x����x,�=,��-~	J�S%5$���+���+����h����g89>��y{@涗$�o�]�B�r�5ܓP{d.j�ok��M=)'_ja�/�$�Ʃq	p���ګ�ȗ-b�����Q:��g-���WHM!+�o����9#���=>L���9/��[f���n!tWe�sq��L�`�h���T&�z�Rxo��`�ۭ�A�!� Y�TXH~+���B�D���v�N
�B�s"���bG[Fpe����o;�6(H���d>1֣.2��Dk�O��G(�n��G߀���x���'�&+�hq9I�ҒVI�Xx����jO�Ą�ul�Q �i�*��̃�1]�0��_���[��+d,�Hp�5�+W1�,5�M(�0�˃1ہ?3�ɐ���Q]��=>���`%6p:��C�7�
V�f �rBG� ��	"��%��z�qb�����s\BBT %�����ͱ�����=�g�_�i�ϑ�#�[�:td|b||�	6$1z��jXp�$(�2e�2Z��p��pkei�m�)��,&r*fxٶ�ܬ�L���Euz�����:� _���hAr^����[9Ҳ�q�O���M�orh�TM���s�q�"9�-~|�DY,�t��_����P[��*����d�>��B�~�屏һɵ:b���y�Z潲�f1B�����&�A�Gl��K�C���E>��5�}�PRR"�Ǣv0��+1Wכ�{S_w+��tb@L��S������x�xdzR�)�敌?��������I)Gٞyq�I�b�)An����1c��xy4,D�jؗs��d��V�ܹnH�Gq��~5�1�E��U
�F�B)�7"����:&��U1e��?�!=��9�C1��&���7q�%3Z�P<N�DOvƕ��Y�^mE��MѬ�y87  /PQ��b��l�Bθ�'8O#�yѸ^��L�]�{G
;S�_��T]]]����E ��������mL�{���;��nf�In憄��秭-�P��Q��jWB'���y��ڗ��[�)�̣�>���4����.<�f[ǄM �B�dpGS܉4s�re��';['���:0?�ݿ�b"nsӂҷ�����v�k�hDY��j�%�R�� up6v�@8�I&2:����!"�D̋8P#
�6~���RZca�&7��y_(X�: Y�A�B&��O�x��
��\\���[�?>�hjh|�'���j�׆R�s��t���$$�'\��f���m�����M9:�*����U����͛5�<<yk�Y�&��QСH\//.�e�'��i����h4����p{;w$�:qd��f0}���v0uh��'�=��K�[^��9g\<��� ��q9M�Ge�
4��>�w��K�t���H����#d/���k�0�9>��_�T�_���!!!s777�ϸY�iB�Ȉ���E��h����Φ��E�y��e[gڠ|%�L@Zů�����1�����6͉K�%F����M v��LH�$���!܀��SZϙSi�=��g,}����8O�����ѕ��x����P	�TJe)Ѩ�ʣ���=~U�|�þs�ȍoD��L���-��C��o��V�b ��Z�! �i�rrr�v�J�Ǌ����@����m��A�"!�����T�c�aR]Q��/A�2�t���q�!..����z0n�D)������l�k�ne�OP�I!�����-��Ǧ���6�2�_t�+�jE��ӄi��ßj��~zh0:�0����y�ܫ��(*�{q�S���䏮0�S��tn��܁�,�-��5���O�&"�m1k75���.Ѕ{���)��
���g��t�'�V� ���QIA����|S^I����,��Ʀ���:	'�YZ^ު*��~?�R(տ74�!�V?�a*'���1�ɢ)��e�	&�-����� v�>��Q78��m^�F9}�#:9uɗ���0�q��Q�3��n����}��o.�#��L��Fk�+4ӌ��<�=v�\��1Ʉ�s�L)�xl�e��k�T�/X���w��T߬z2)�����_�`(�8�>oW���<��}������V� HR||5��9�%3���ȷ���rp�`~�-N���o2���R���%�T4���^h�D:���cv[s�mC81�!|k�z4\��I�>�IDS�L,�ZV��Ԙ�@�1����@ى�%<̂�!�n	T ~��B@l?*9��[f����
OV�������U�W�l��+��oHH'7W���R.MjCi���p�;��������3�X��$I�lJ}������(�YZ������y"�ۗ��]L���#���C�d�域�?S*� ����Ϣ�&rW���8ߝ���7��������ȷ�����Zuf!+�u�!��� R�^32���J�ʑ�A�,����%�ju,8fn�7���ʠ���+�M�)ă������ "��ي���c�G���T�Z��I����}�Q�d���A�z	#����eFJJJ����Lmmm*�P��ߓ����_Nۋ��\'�sss�i9\����:!���7��c�$P\�J�:u48
N��lC���r�Ry�eO5�7$<�:�M?�6B�Et����\|Ud|�_VD�;��PC���y�0���Q�r�a�m���L��Ҙ�qT���\�8��9�,,�~��&-��DZ��Id�!}~��Ae��3����d0��좋sǭ�J�AtZ;�H��ط��f�@~��9���z�p}\�&�ɝ�t�������~���<����L�`�L'\l����5,���U��c���!������)2R�Иq��kq��~��?8��ǉl_wx�pc������Z�t�vЀ�Q\���:�iP �n�w��-c�W/-?#WQ��-�%��W��L�'�2-Վ�����	҉��NЖ�ղ��%��$�#N{i�𶘘�#�CC �4�J��xd.^G���ڵ�6,	�H�����ʢI���Ð��������� y4˔YH�ތ E�ALM=��l�uf���d�D�d�)I@X��kv0U�%��x��ߣ
����an�@]`
N�d�DOqw��8����![x�F>�3�;�_BY���/��"��<����^]ЋK�T��qa���E6-/��,Յ�i��S�c	;��j([ȧ6���������R���ZSZj���.f�/{�n:�;_�����3u�#�C�m|�yxJ�)���ZH����e\���G-x�����a���p�(�.��ă��|�ܗsR��0C�/��&�p�ԅp4i���xW�p��/Jd��~ޡ<�|���K":"`P';�+����=&ܘ�����(O+��^�&a�vrr��0�7��J��݋ۋ��Jt�l��Oy�}���n�B������l
��l|Aˈ����:j�0^\�#K�=_N�8&�O{ۊ%��-ζ@�oq��d��DNNj@Ձ���!��2�"�y��d�wņ�u��.�����4C��C�U���h���$J���!L�����x��X�� �҆_N� j�)�G�#��.��v��hf�2��L��.~P�C�(�YZ�O¹3Y�x��U-�<e��,]����++�`��H����%���f�6��6f<�)�$�����4&���o�����Tt����������lo�'zL��Y�@��p�=+�a>Rn2c�t�!9C�r��*h�
"ȸ�=�b�Q�\�Z��Y�4��Y~�@չ���)@��ފR'�
��dv:X��w����m5s����t�O�?���14'r���3H(���z�r�߂�� ���e���T>���pP,�1̇x>u��-HR^E��LL��^_��[[���R�1JPZ�9�b�������+���PdZPVƒ��gQ�*�!�������$w���~#��;։2��P��w��V��Z���Agz�t��2�T��CC�I,�m��6���2tsM���d9��0ܒ�d�d;��K���Qh���|�Ί��¯�=�i���x ڎ��nk��M����D�z�������,��@
B��Lb�`�wwh�:a�k�Y��-l��Z#[U��3�l3��z�g S��Qx+a-AU����X�5>>~u�p���LT �#�͋-��G�����o�{!N	\?'HcՍ`бZ�Y%���_�@��r
{SS�;�z�����$c����0G�>6�@4�[�+�Bn��g� ����6�,2�Gh(�(m�NVq�o�ܼM���Gb��o�aΏ�;��e��`��j;�Dgm^l�gn.Lx��[��0D�oh)졯A��"r4W�a��	5��)�l��0$3�0�x~za-~S��_�6�O������UO���&R�겲���_��PQQ��������*�hꩂ�N.�;���|4KSE,W��͉�V&R7%�!Jy�=����L�h\�O����%#�5"��+n��?���:x�����8�]���bq��bk˫��!5)|d��,���k��%Sjhu�?�1�d>�p�|���?��|��>������ع/
ۋϙ�-H�ʛ����G(���7l6���C6XY�_�E��l����]�h�-���ʊ_/}��#lS�� ��uA&f���v�;����E3ѫ�_�rO��΢�C�"�6n�p�p�8د1�|P/VQ9U"b�CȤ2��s�=�CῬӚǫ������~[��Fɒ�r�+��g�$$���x�GTwr��h���4�幠��Y��^S��l�\����3�Y�a�0�ۉ����e!�O3Nv�X�
�=**my����	K�i�$<ʕ�|�Y[��W�9�C�*V�`wV��!���'"��_����{����O����������f��O2Nt�I�`R�k?7W\h�	 ��Hnf�ۣ�@�b�����n��p���'�~����x��y���z�:,e�� ?L����V��U`�f�������Űw��\�7r2�R�0ي#u��{��N��#�׃�!�,�붞n�����*����q�G<�qSv���"��{dA��ĭ�#?̵o�b��u�]�T4ԧ������9������k4�P����l�
�~�uJNAsB��w�d��;��3���ň����$�2�wϲ����/7�X��4�pP���D�9���ά?[/
*�jkbf&I7]S䶚������A��Ԩl֍�{�8DQ(?1�IB�
����^��}8��¢�£����+���?~���ġ�i��޴4-@�G�7�w��y��1�f�a���,���������=}n�������9m�� ���T�Ng�]��c}m
�LP&q�5�����G�5e+�bь�0���N�b��J�B!�)�
��Q}u�W�ŏɣ�{a��J,��\Hjmup"�<8�u����▜Nu��������7�_���Bf鄲?�m[�-��|�����̤���b�1��نD�
>$�H΂E�LWs_�������CR�I��W������x���ϔ��T�\.����ɼ1F�MQ�MO��j3���>(G��#q�vx�?�7��k���cp��f��b���o,(*�_���iL�Y���`pC�d�'9��0Q��Gn��ei�"�k�h�ى%��b�Y`\�1r�s���Q�;�����j��L)�TW>�?�.�}X��b/�k_�.r ��Wg&���o���������C�q��2���F�Ԡ\��c �#�|SBگ�Xd�x���)�»��ڽ�t�5��b&��6؀�X8W��,�=��f�A�5?��U���֖�Ʊ{f~{�n�^S��!���z�֥�a@'֢R�Q���܂���r�'&��}K!�%q����;5��.��Yu�@@���^�(�P�K�חcO`7�`���:����bD秉|�}}iC@�g��fu&�`�iJ�eME#C�t�&�hH{  �u���Q��7=��~k�994t'�Ttŏ���Gz�E���~��r5+<�R�Kd�ە��'�gIbvG��PJJں���f�s�D����w��6����8'�	��x$�PG1�)�Ruwm8�1]���k�'0r<5]I�
ʝ(�oS�~��v;�DY�l�Ty�e0�<\Z��7G�O�:4������׶-�$���RN����R���R�XNMq�2������j
��کh]B�{���N��Lӂ�d����i�`o���q��<�w$)��_Cg��78G-`��"����i���*�Konc���ڗό�+����*��@ui�=7w�oB% ��
!׷��Gv.�Q��<'l�n���
θc0�$�M���@��W�J�:�$L�h��{\�Z0R�ѯ�s;0�Z���q8UB�����{nbb���V�@\�}���� �ލB�De��k�I���z�I$'�TX�0�'� �
��ʣ�<N��.�����"��A�P�M�3C\���;�%���Y����\� ������d�OY�)(�}�:L�������*�����n�$���geP��?�^��}hQ&�(�q�Y���>Џ�%-}H���<�����(E�z�F��T�y!)�B6�)5�qΡT}���9}����1������ܙ��=�ZMzR�"��hY�5}lq����&I�V���ij�hq���ҬQR/�g`�On#R[O]]�F����S�����_�����\���� 7�8��L"I�jQ�6���6zz�ٍ�3#Kf��~�~���c����2���Q\�:RR�������D�'mpnt�#���Z�]�kCl�DƘ� 9�!ӓ�^4*`;C7EiB�xx\����0V0C�}4����%�ɵ������(XXRR�Su�M�$��$z.�#|G��"޾��	O.U�$����V���Uhs�bΜ�'�mT\��%ta��������Y���;���+�Y�F��o[� ���-��f�8���?&�54��t�/-+�I'�G<'�}�b�Z�x�ֶO��s�ޫ,��-
��Hb�������4yOu"��Ba\����q�x bяI�Ɏ坬�L�K���E�`�q1+T��=8&DtKѮM���4��������E7l������l�%u
�ԅ��A5��m��e4��\�Q�O���ƽSj�V�]��Բ�9��Z�w&�������-L2\����Ύq<�x���8��+���c�ߜm��w�V�_��ٳ������I�uD�lq���[Vi�SN���k�*��amx
J&�f���p�t��8��~���X"���RӘ�@����K/[g磯p�h\q+�CD&�}��X�`ָ6@k���1�G6��#Y
&�6ܸ���Ý�����3�;b���%ۏ��VFBF��0s &��ɾ��I�X�;��u@�|;�	#wV���os��t��:c���Xz�q�v<�����ݟ�ߋ ዻ�������]����o��%۱&�e7
O��;�|����zU�?;]�й:����GG���U�q�3�.B�"=�0a��� �*Vh�?Oį^�-,��YX�A�u仝e�LXv�ȷ�����c��n���E�V��/��H}.9�����&����1P�b��� B��¿���U�p�<�`B�6�-�ń2��b�Vv�kR̼jMu��g���R-y��.���)�6
��:k���]\\�M;[$%}e]�.S�m����\���acȢ���nOLO+Xp��j���7W})>_�d�z�bG/�I�i�C)нÃ�2d������>�=�l�kɃӿ���f�����hr�kF�C~�;��=�[���
��c�p`T�O\?= ������@v6Y'�k�p���?��p�a�4�
�°D��L�,7�v���e�Ev�s-;�@>ζ��"����z�6������?%'������WV�p�}��m�9�%�U�:9��E���y��H��t��p�"��).��@~���k �����"�?��I=���������9���C����j�E�p�ȴ��b�6��_��`$;g�{��D"E�T�^�`R��s�z�ޘat,~*�A����>d*�׉�R�`��x�	�,�C�1p�����J�2�,���9��MLͿ��<?N����T�B�`�TIAl���^h���*J4�O��FlK=W)�J\����S��E#M��8������E��9��`d����o���PCd4EB�*�:�A����o�Z��\Zs�XT���C��@��#������V�������W塧�T~��F7��瓮~�=����M��W-׳NS��,���7b��k����DЍm>Q��9BS���c�h]]O̖k��>읥�Dr��4��8;9]ls��C�Y�Aq�iW?OY�}?ŧI�6�7��č#Q���د��ѣz���NNM9�
���}�1F9D�С�M�H�2	Z��xK<��\Y��t1O��t��PR9���B�K����\!�ڻ��׿�U�|�ٵk�@4S7<j�N�bÿ��uEd_�5�6ה��1���F{���.wE�j��?%~D�t��L3�a������\\��<�z����@Ѣ:��[�qE�U��7�+	��56���`uT���YU���#�eʨ����^{��<|l��׫l�[ԕ��A$�z���"y��[K��dV0�AKnP����=���K�I�����x%����SbJl���G����-!#8M��
�wR҉�0����2�.#:,F�~A�I"����e��c/�.�s�~�7�D��aQ}��|_��LZG@�_М���WR4ꩫ����R�b�>�w��X�FF�/݆�H�53m��-V�������C�BPr.E�x���z�<hE.7��>��~��9���A�E���C��7�e��=����d��*�v�Q7{ ,g�X⏪&���&���M�yf�6y�4sR��k�I��"Y�~��OπSS䇞瞭�����⛚tyF�6QvV��f$A�u�~�Ds L[�*������Kq��>�xr�` =3���y�F�r��G�f
��<	����Tǻq2����ˉ��~ (`H��{��}b�����t�#<*�b�j�P��51��.�'��ƍ�4	�X�N�ͪ���KV����|_f_I2�׀I�w�k�-܁lb��=f�]r)�L�-�IU�"{;��A��S��RC�g�C��I&V��NTC�
�GuŒ`������]����k"U�E��WC5qx8� �d��hNjj�kѪ����{��6ĢO-�P(�,l�"����}��n(t����7jp�K7���胒^$ 4�6.VTc]��N�C������M}W�d�8��8VT�Z���O��|�d���hV"w$+A��J���`T�Hdr���3�����s��:+��`c��ޔ$�>�����b�ƄAHހ�x?�该۞��"��UU$Ks������C#�����u!b���~X�_t�QR䈆�}��� gYA�$RW��8�nO5�kvv|�"Q��̱���	D�N����յ��Q
�$���%{~P��K����KY��׬�g�⢥��O۰3�5��+md��@�9�>����"�YjJ�L"��}͕�������c��r"N?ͱF��[��ޒ4��ƒB[��U�E�H�ƻ1�����rXf�:\�KU)��{��*>K��&<�Q˫!������5:�`������g���;&�Z��Ԕў_��my�7M��8��{�a����Z�����1����HW-�YJM�ѮFB�>(�7�Db�3U~g�i��lU~���v��.�ȴ�թ`�	q�C��K5zo�nZ����VJJN���K^.��t]���j���E;���ǽ��9�)�J�>�{��p�E�a28
�+�O�:����I]Uj*�L[_*AQ�4�Ų#�)�Ze����V��&\!��S�mR�NV]�AR�F�V��A�%�+��0��lRJ4���*�Fl;��/��������ܑ�������ۖ�>�R�����,�5��?�v[���a)_c�Ӹ�t�B���0�/�+�{#�g(�Hogo_m��tAQ�$&�tW"F/A�"�A�M&( �ϊ�1�
f����a�e������hR.�|� |f����;��O�-Kg��R�/8E��,hpi��������w��d�p� m_!��4mu��6���B����	��3P������m�OWP5mm@V�1���S��7*aҩ#�R��ӿ:�1m[�8��FF��B^��J�&ӛÕ��D�/>����Nb b�1��d�ÞV�R���{����s�h-޾�:���j>YYq-�q��PAϻ̲uꬴ�	h\֓��)sn���-��Gȱ�k��X�~m{DyŰwZ�F.����8q��ζ�����E���y`��߶��+��QM���<�Ki�Iܣ����zr��/œ��o�($ӏ��d�������5��M�L���ֿ$R�Cn���oTE��H򊋍W����I���hjߡ8ܞ��S��-�=�t�QHV�'.��ex��[Z�V,*��Ac��3$sKaE�\Y�p?R�HyV��	��9��|n�P$��i{bxp.�ɳ�4����M䍔K��1�(ji����-o�8T�QJ��<��rA��;譴��+��H_��I2`]����U���u.M4 &3�5�CN����
���Uo��"�l7F�.s��Z{Dttp����":��	1~Wŝ�KRe�k���,ۧF�aCy�C;	cl,���pRᦆ��o���SqhS�i�[Zq�m��-�����u;<r[��15�5��) v,�#�ptt�GcBuNN�?;w�`�L�k�1�������Q�Q�y9�X88�zkLW!����8F��$�%"J��ǯ���$�����s+��86����r�RT��ѡ�ع�D�捺/��C�z�n?��iKm����@��*�Idی�`���a�t��y���x�sՃ�W� ��~���S[����%G�:3�_��D*β��J?AH;;?��o��T�[/g�Fm��Ze
��@��A��CO�7���}))��[�Dz8�v�"�P*lO�3��G[9������ 7'mr ]�&囐9�A��ܥ�bԃş;���l�Ӿ`=3���@�X$�#���7�����	2�;��A��#�3����с5�w���)�r�0O�j��j��ưX��'f*��y�y�S��:��� �>���J �U�k�}��,k3�J��6���¬U��jv�K�E�A��2��_���x���O�-t(2�׋3��_�5ӵ�SGV��c��m~	8ߴ�sP�B�mƹ�+պ��/9�b���`�_���%��'&,��z%-���[*�;Z��X�*��^�\�ܾ�LFI���vj���y��M���?f��|��J��E[!ؑ����QhE�g%�ޞ	���ؕ�K��^�~\��~��R������8�r9o>%����p�ԭhz�?�gU�����v"�7��Ҡ������bJ�O9��>�{����[�"��_�kF/��)��^o��[�ޞ��Z��˻bsAOЫ�����@�����Cz�?�֍&�z��2���G	?���(�)0�ˣGe�9�EG�!	\�~���3�F ^����cn;rx�T�#t3D�k���EK�FA���u it6ǐ�@���`H�����I��@y�r
���k˕q���&}���h��ih3 _O�l������U��y�j=���ūg�P����;3�f���6�f���j�[��&�;p�3!�iV�g���%'�a�c3z�-�7��,e����>��f���||�}�`ŷx��Rb�1p�=}��n[�
�Tx��.U�2�
�&��X}&�QlV>��ж�b�:�ʽ^I��N��?���'�9'�I���i���}X������Iס����JQ´����,C�:�֡�-��4����ot�����f��Į���_����cF���~����w���������y���x��X�K1<�Ę�+�h�@s�+�`��RB���J�����ރ�VV~oy:*	l���k�?�R�#���i꤈��mN��c\[�epq�	KU(Lq���
ECT�A4��+&��j�0��ލ�ca9`���� ���#������-���of[jO�e�ӿ�!��r\�Y��b*c+�/6K!@� ���]��̇[MH���#�� 㫢��Zk���zK����?��A�{�9��Z($�
 jr��c�!m��/O�	H6�
�q�r}�M�B��N�F�>�=��sR<��vd٩�d
	�Z����/�r�����T�Xɴٲ�8��yq�fp�����X���X��y1�k�,� ��K�x����,�=��ZEc��8{^��^�����Qn�?V6���|�¹���b8���f���V'��OF�io�$g�IW�md(�PjB4����=��9�c�r~����-ɼ|FS��$A�N"Š�P8�2K2�Ei�����M��pd7�H!�������@(��|�3"II������ծ��,�g>'��-+
��x��)�<4�~���òԙ�����q�_d��"����Q����/���(�b���F�Z8�޾��
�P�pf��% d}�������=�_�ET�M�y}�2!�`�"��6��AŽ�0�.�6�Ѵ1fnnY6{�;�Bj��	�$j�"q�19Ys:�m��W�HQ{P���S��`j�^�����o�''�y��0r4���`�SEf��E�b��,+�1�[�c��SI�]�J������o�T����wI��FǾ��v-�1��8?���mEՔ�F0�}�G��Xc,V�ʵ��}�'����5@*�O�]\$���紖�a̕,�8�>�J��j͊F�W�Ih����T��_�TV���ƿ��Brk<�v������ ��^�]�88C=����7+���v	�ZY ��ڐʲI�G/bi��Ǜ�%�زa`Rr6ڣ�1 j�@�hm;7\�m�L<	���5��	�0$��Ľ䮛�1��5x��Է�����%�[�O1u{�sR�r��Ԓ���i��Pdʒ��\��M�����w��[B����,k���$5!{��v;vxϔ�D�#t]Bw�s���1�s��Q�f(�:Vy\��W��:�[�DN9�&���g���&x�����c��s?��h#%�R�.vR������=�	�SW��Vo<�
��=dgh�����ğ�Y���Ӡ0>P���n��>������ϵ��TuҐL�LQ�ݶxũ�������0�+�LcsK����e������F��(rqv�����C�B�䴕yt�_y_`K�!{peH�_Ç���W�J��q=�Ls۸��U� �1���9���4��2U�9�GE���|�hi��9� V������(�����Y�]#��+����H�r[=�R�䋾�/3���t⸅�,��B��D�_�Y��c�T�O�~�1-&�1��X?y|�]R�(�^������^��)ns�BG[�n�x������"�Oҩ��	QSg�L~��?��q�4��I4��p��(p��CG�#����-��Z�zz���1��ҧ�]C��QJ�>|D���/�zIĵ�sT�p�[8R�����ےk�R�H]3/&�2it�mS,�a�s�,�0,�w$	�HF���!���i�2���,��Q���A� $(A�!��cl�8��+IY��^���@��"�"�P�w�s�#zIϕ O�ܒ�@1!���i�_���O6n�Z�8�S*5���	q�3��X�z�<V�<���2�7Y��0w�y��l�uޅ��-��N�gw��g�wE��zY�[鸪mDZD���<M����Vlf����7�D�����	��_����3\��-ʐ�-�CX�K��Q� �[�-�g�3�ܩ���9��2i��ʑ֋ǭx<t�I���p��^����\y���i�s�E��Ϳxn��9mX�i;X�&b���*��څ.��r��4�Ֆ���Ӹ)jo.��[I���<W�=�Kg�*�y�D6�/�k��~�ߑ�ǻ�:t�p��nf�RL!�)C�����R�����lkR��u�aׁ��777iٹ匶�����3N�}qP�.{`q�+ؼ�DCA��Iӌ���s-�Ճ�f�g�&e=P�y*f��`�Z4��;Ε�����Ⱦ�j���յ<���i�RU0�辪Q�Rzso��jD�Ir��>Qk�L1S�ɊP�-#d���=y��#� D'˒iܒA��,�Zu2E՘�g��ԁFu{��E;o�9��9�Mî�MY1�?ȗ,n�	z�Ne��	���K�L�l5)�:?c�A:��.�.՜�ܦ�&�Ok���L8Y��`TI�E���+���;g+��h�6��xX��@��O�"�z�/[-����]��ӳ]��P��ٕ0m�Y[q�B�Mն�2�4�L��Sj_��>��$>T�μu#�x�60��I ?1�I�g����U�#��u���Q6]#���Xa�Q@Y�uh�'���|E{��p�m�x�V�I4(v�k���c���ηc1E��(����JOo�,/?���V�����%�j��JDWF�BG?m����fd<j��`a����ͅ>,�"���>t�K�M�^�3wlh��������ť
R�%+n~{��ɞ���eq͋k�I��M/�(�87J����`5��u&�zދ���`oL�ά�����F�������Vj5H�]�S�E� 0t�܇jnm���ï1���5*Y�3 ����REN����D��n|�x��Y?�$C��	�t_\z��Җ��w��p�l�H��U�>�h=�"KF����A��p���~�q������[�B;�S�Ԝ'�F�'���#=�nYt������~���;���Ϙqz�է�+�%��o�6:�}
�)A��ԟ..����K'�ØU�
C�M���ְ���:tSSJ�<��/w�v�s�}o�M�0�����>����ǹ�����vp��~ww`"-M�T�)I���DY?��I�����lw �O|�t���i6/���@\3�&IL���C`u	�f�fⰻ����C�Ց=<M[O�]/yx_�mƙ�k�.�����a����@Ii��z$�R24>�?w�OU	��]*((,=>>��,]խR����z�+��(A�&0�|'^����is�����v /j�8n�k%�M�s$�}r~>ı +�˖=-Ţ�5�cpU�*���e���%�1��q��m�/�����=&�]淋��8xZF���=��Z�GN��O��:Nli��i���5A���K��W1�:��<��*�C_����-�xD���&R�B�r����/����j�!���D���f��(]ܳ(zXY�?��l�\�ktqgH��O��-)y�R^Rbt��nm�?~��
޹+��� DPk���ln�dq�9X�vY�	�7h��3l;)�nC��t��kÿ�Dk�r������u[C
������00��k�����5�}�le�ee/���ک��CJ�� ��~�����Y�����*H�b��*n��;P$h������pK޻�w���3�9Ŀ�)b�*���2��FFy�>;u�bckȀ?R��_��>���z
�X"h�@�9���)����� N���w{� �Y��ιs�-
�������PYim-~*D�a�'��傜���/�J��W}�����
W'��f�o��O1��S����ÖlT�s �=6��}.2`E�c��K�����O77>�n6�ssۑ��)��X��!���O!������:�h�{	Q�i$(������l#���0C#�Ɩ��z\������(}��D�k-h
B&��26�CJߖ������lh�i����]K��.E
E��[q�B�+�^�kpw�����M���	o�g�cwg���M��v����}n�cb}ۘAs	�1q�~���q/ҧD�z&Y��8q��h �7�7���r�+:�ß��+�A!ӁCt��*Z��mM`�'�9SP�i�2�I�-B���ʲ?�#�I�>��u����q�V˔o`*�1��0q����U�	>��w9r�aN��zDw7�G'�SE{��^̓����O�hS����O h:s����b%VC�,�	��B�d��qIHmO/��?mI�0��O�f@���x��,@+ME�""~��ӆk��n	F�� 蛋�P�z����Q��z�
��ǜoطrI�ⷎ��� @���t`d�2� ��ڃsPʯ_x������4}f_���Yg�7��
S� 7���%\H���/&I�/>�#��;�����&���$F���JׇM�]���:�$�O5�H^(��ZӠH���D��b��}q��;�����ʻ\�t�G��8(s"�&���KE�s�LN������1:@�3��rS�Pi��_Ґ���3䚡��sB�Hb��%�0娐��y*h_*M([�9h8DDV�{vIv�#�ד����يy3�u�H�*�ҭ��A�.��ZD�l��0!!E�*�yQ�1��ny8������@-i���s�I�k%��E0�^c�0�s��a�Y/�΁A0Z�1�!艇��]<⊹��������،5�>����O5/���4�sD�O�-`MJk����[�?
���ƨ9��U�=~C����d���Z��)�F.90Z����Y�����{�������K��A�BI�(�Ac#�e�nڮ�fL59Q�h
{��6�Pk�?z��]Δ��P��M������� �3�ׯ��͟�mk��]�^�� ��Ob�UvR�gw�9��7�N�S�$���9�׀ߞ�E�$���t���;��*��`�w�(�Fj:K4C�M����9���&o������R�u��6�����(����\�.�&B2��a�����0_�fk|�2tW�ꈸ���qh�.�!T0f7���ܞ�(z���P�aF�a®�s�(1.1Q,J� MQNm)���:g��Lj�}���]}2�J��?�%哬��|1p�>�����"[L��3
�=���(��Yu_X[?;^L{--�~*	�C�A|�>����&k�ћ��0��1���c���нHl����%���L�~9d��>�s��J����秇�ė��\\��@ӏ���<��aq܂��Z��2hRR�@`���S����ᡸ�OC�S��%�jlj�e�e#:�.��'E���� �@�ǝ�
�Ϫ	o��3�t������w6���Ǚ�[y��f�4�}��	�V�Z��tǱt���ps����h��`�ey�ck)3�6a�q�ȁL[L� ?x��}��h>b����n�3�+t��U����l��{�~���!tGr=��`W���	s���o�Ed�>(�0Ag�r�����_	���m����o
���.��被�)�}N`њ K�]���;�]���<GKΛ�����w"�I�t��'M�&�X��t����"ONgfq$,�7=mݙ"3�����+qJ��d�cw��I�����
���?t��l�?#�,����	Ý?�68(���!�HO�PtZr�=����P���֢��٬r�؄r�U�����Y�on��"�dP�xrI<r%��G"� �\btOxɵj�zɏ�[�u�z�p������$I����tq�͡�H;���}���Tt/��r��1?��DӢ�+��i�x�#(�_.
�%��>!B�c@�A��:��ꦭ�������4�ݍ,���.�i����o��FV~T��#�%�l�-�h��?�NMa���w�~'�	�̙�|�T���>�;-��ّ�o��������竚n?$�$C,[��K����}����>r�̨�����gWKC�����/�"U�I��g���W� �8�y4d�[Ea�۪5T�X|�^�KП�<��' ��"&eh������")W�1�ld_5F&#3��Y0;ͻ�$�]�q�f�M��q�
fK�;���9M$L��Q$:20cY�/���mm��N�e'�L���<�n}ؤ���F��h��㵠�
�Y�zM�ؘ��ծ-0�XS�7
���+�~���l�L�i��%�����]��!�D��6	b��|�"V:��]gŮMʾńE@�ǚ�n$�,\o9��v	3�g��������!3s!�#����3C\>rp� �Lk,��a��[�lֻ�ÈFN>�v����(���m;:225.���z0QY��	���,�t��EF�+B&��:(f{����������t�ͨc/Ǡҫ���}��e�ܳ���"83��;�����C�� f�R����HF��n�v��6��C�p4ʽ��_���~�ǂ|�c�vQN&��\�J�fd����<#xKז{�C
����r��+\F%7�� �W���h��+���I=���e">�s�����J�/�cL�Hj�= �'4
���Ö��u�K�fnn���rU�H��������b S���y���壜���ݢ��dm��<:���h>��q�� X�ǣ7�s �Aǩ�[��SS�N1�q�Ź�ƻ�������"���M5��^��ɬzu����F.�[���~~cA��O���wK�R&`��+�Ό��g�V��'o!|,�p(�.�)�5�SF
Hw�ml�O֘�������FD�s|�Lb������h���M^�M��\]]=l3% A�$�m|���'$(X<F!��$�1��[D�������_����U�[��μ���%��M�#��j���YX�^lEC�����Ҷ.�#Iz�}��]0��+Z����7���q%�%JfmR���?WB��G��k[��/q�h���3�X��Mf6
� ���6屮�;2A7,�
��
��s��l1�r���H��B��2W)9#�ON�J)����E?�/��h�F�ώ�Z��^��2_�Z'�m0V}7�kg*YA��������5�G��g���ֱkek�V���33۸��rGq����3�˺Z:,��a���r��>�**q�����Cֹ�7V">�0ѿ-v����9���R3P߄%�TG<̝�	�􏀉��������w�� &�=���L79!{�˗��ZG�e�!�">�1,�K.�ccc��l��o<Yl�b�4Y�~pq�Od]t#�n �����u!��'%%���r��Z};_U����t�����|$���;���|��Ż���9��*l�1P�s}Λ�]K�C�<57����[`�0�����Ky�~�x���	����)����\�Mi�A��b�+����=�q��4����{�-.W������Mq��KK�����bE���/t�Q5�+K��5�[�e
.� ����+�+h�W�Lɬ��ܯfҝ�V���r�����ߕ2���(�_��ߌFF ���rh[�i�[�>�AI,Z5��[݂>ܶ?��w&�E�H��u�"�$ B�Sk~�!5A�rB[5IbB��b�������l�ۧzHK�z�����!��ƦaEJ �Ƀ�Be�N�#��J���;�	Aw��3O��u��ȏ��c�7ݲ�C�������c�F޻;��{�U��Ʊ�@�(thap	��9f�[��ٟNgT���6�pr��9�Uo������Χ�Χ�Ye�W�V��wK��4˱�Q�y�HE�9~?_ʱl�P�����.�͆�l��L�l+�`mdiy��Dkp�N�Q�����ӳ�ZV�-@�J�rz��d��>9TuDG��!�j@#A������/w*��%��� tg[�pi}��]Kzee�	3���RY�8A�mR����D� _</�"C+��2���$E��H�e��co�qJ�O����'?Y������H��OH�0��XC���p[%ٯz=+�ˇ�{�QXOT��1'E�q�뭱��|�;������c���s���!��0��%-�L��V�zƼ�R�t�+w���=�ZFg"��L�j_;�������:F����|���[��������	�-3(}���q%�޽��.k�pe#�C5+W�V�1b�����`[XXt�W轟��~���ؘ�����?�w%�D�ݢ��h�;�#�r��U��Z0/s�|���O�LJ��cO|���8��XN�gA�����3��	����Y&U�1�DT�!�1)L��y���igu��\�5w���V����AQ�> tp������l!r���6@�tztԑWn�j�ߞ4�R�-h�?a_����!�P{����t|"#�_Q��]����*��@���[�L��$w	0�������˨�\ �v�f�h.c�bi���&����-}��>5Ω������Ə$�r�˗)�~�d�N>{����E�M͙��m��iqɧ���=��t�����\O��z�R���|r�}�ïv�ԹT�����>hE���v����/b�!�bEZ�k�������r{�!����з�^�[lT���CcU05���'�����T`p��c�$x�0��׽�8d���(���i7��h}A�֖D#CF.�� E�������-��K_��h`2��1l��:$!!m���%��0�g���Gh7O=�����	�K�jm̌�l�xX�
P�]������0k�B�������@��0�1���auo<#����2����J�ZC< �꾀��@����K:$�H��ty|8���w��R�$Y>����N{[�2`S]Y�C~���t�#���ճ<�g|�Рuxȼ�'2P�*�{�h����,.u3�>"��Z.��9���ώ�h�n���$��1z��L��;�x���,6ؒ�H�'s��q�SbH�z`�	�b���r���+O)|��[9b�P��d'��u)������,|�Z��QQQA��|�����������*�`�J��o��v�y%�j��$V�)�h���kf���������w"!�����r�m�斓�������e��O�m.F
hq3C��7�٫�c
"�k~X/�=9��n��劋���͚�*v�Lq�۴��(x�� Lng&���������\���tA) оl1Z9���͚M��l�K�]�DdkQ��3�`��U���-iu����w��Q�¼�=��N�q�[o��÷v�	�߿���V��PX�������v|h���Q�夲�<�\]벀kg�(���p�D�~9p-��E/UO�y�=%-�wt�D�pGP���;11��ŦDĀ>n�?�Uj�b������A����t�R�_�tz���2���f��Z[˅zw��j�:fjx���&���'f��캼�B�͝$�o"�*>;�(�[7qd�#���,uFh�}Q������*�4��;E��0�Do?����τظ�q�� G�Ch��lGB��5RǶ�m����Df3��>Rļ�s�uo��DR^�^d�+��^ �IR��S|PZ��-曬nz)(�8ݮVe(�Auo�?����YE��ϥWYy]m5�*�߿�י�6����7:�Th���uVbn��Q�7��(����j*���ii���-��>���O�y��-LA����q��ˌ��[�W#��fT}�[�X���e�F��	jm�3�@p��y
�	�����uߚk��l��y��Ѡ%H��㤕��<��I�`�Ko�A���D73=����|b뒨�&�ylO��4�A��&KɊ�Yq9�����mT�&v	O���vZ*�s
���;�u2hX�gK�z��L��ڈyJ��I�[V ����������|��u�C��c.-=*��wMd	�+[����T��B�R�@p��$&K���"vBڍ�!���͵['���������}��n�m^��@0q�&���⡘�ɍ�;ϯԄ�a$H������4��������v��>�r�JM+���b�'�+m�����k/b���7N�Dxͮ)=5f��<�m�HP�1�(<���=������?�:�.��*T�EЖ<�B����O0QQ���6�/1)��	k��!I7����D��CB�-]���X0�A>�F���\���������ʊ���j��-���We"{����ݝ��0/,q����wt���{m���C���c��]?S�)9���Ö�c��m8���#K���s���xE�[*$�BQ�-i���lí=�Q��>�z�c����U�R130gR����y�� ?��eb��_K�иAr��iUf�O>^�����i!�p�{��P}8�8�L
AS�����Iv���5��Z�e��{�i��w����w[�(ݖ�6o�[��l�L"u�3ˍX��J�}�0b�Ϊ�q�S��Ҁ��K�9�%��o��	���U�9S�]�}��A8괹p��v}�{/��9������҃-o9]�@�^
�7����!{G�!h������BJ�m��������!��e�� �r���1�΢��D;����Y�I�hY�nG�:�^i���U����Kx�[��Y�7�u��L�_)�^4��B��7�l��V��n��7GI,V�X�?)֞���{��*���K�s����x1g,뢅�iEDPkk#AW�v뾴r|,�&���B/�Y��L���5��(-�A7H�Y�r
�N,�8�Y����B2�;��v�x\��MH@�Idn����6�[2���UQ��]�Ȭ[njǼW#�&)����Ӡ�������
?���uO��iS��)zfFj�VJ�G����v����$̀�8�_�{����a�Ͻjʯ;���᭺�{7�J���(!�d�r�a�� ���J5�z*jAz���x��=�Zm�BMLT����BWHQ�p�-w� �>�9�
��W{��M\Ga̗8 ��V'�"Y�;݄	m*�T���]��~u)?�A�k2	�%���Si�
���Սc�E%�h�弎�߮sĴ44�kj퉉��l���&^�A0TX��ռ�+��mƤ��e�t�8��1y��N&�u�A�h2�Ʊ��P�'<<)&�������婵5�ݑ]�������~�*s�}���J�r� b�_�Z{{����Τ���B�?pc�vi0�$���O,p���Ji��<��sNN�����B�4���}�u���r�fS~Y�w<�L�����:E~r��pc�Rspx�{�H~��WMs;F88�0=q"a;�-�%!��1����헯 �\0Z��]��x��Lɀ�%B����x�k<�߯�V�fmU>��`��ާ�ܢ7te�OS�s����`t��c��y@RD8���F���@�oҎm��hdt�:�꒹T�+�Fazm�8$�qŃᕘ���P������C	�5���S�_	��">wOe? .f6��js����V|>څ[��B@��[��b H�*�YF6���ˋ���Y��;���20�@?ߑ�4����T�G���}�a`�������0�e4�����su*�ʝs�=����u��Kd^��Q��M`:�}T�鈄�!�w40{���<����N��v�3��@N�,Um"�CXl�kB���֮����J6�;�޺�-���x�yZ�Y��VIa�Y��{`�wG����P��ϯ��c'������}��L�DO�븰�*�/ҙ��9�uR6�Ý�Q���v��y%i۬-����Dx��Z�>P$�ڨ\�t%�E��;}aI�Ϫ$��� ��oT:S�Jz���6���&}k�PbnK/5���gg;�!��D�&���x�뽊�Ĉ�FM�ߐ}BB��a���X��xB£���ج�E����c�s��I�1�F2l�'>#��-��%RR�u;G�bh�@�'�O�!.��	��¦�?��(��jē~A�qba����r��~,�#�#���Y������ɠ�H��TQQ�u��0x��ެCf�?�ͽ[�F�
�??? �-�k��O�_	�;|���Q'ɓJ�Nx�F��_߁/۔�~������6ϗ��#�҉ް����J�����c�G�:%+�/d��G)&�Y���_��q���ؾ���Ր���m�xF\��_�(�ay�oC(5��o̤�@"C(��YK�uRk9Tj� �C�	\��f����6���k�@1PnK�P*�ż��س����n�2RQDt	[sz�/�����2���G�KH�|��7:8%��!���Иsw_`+�o>Tc�,�%�a��

�<��[ 	
.��;n �f12�M�(l4�w�E7�����Nn�|҅.�C^s�I��Xg��C���D7��HK������Ȉ�&��� ��!3Sm��XJ��5�]Vp;$�"2*Sle�V#I�	�����d���XL����y3�>��7[��ԕ�%�����V���t��w���v�&l�o��\n#��wv�}q�9�fﾡ����R�F�5��i����m�1���O,LL�������ڂ:���</a���:�>Ҽ!s�ݮfW����nD�f�H�k���H�]Aʞq�_C��
3�����"�;OOo¼����T�A���M�6&�S	�Z�P���s�m�<��68�1:y����y�YT�l��c������=���"��Vt��"������(V��ͻ��iW�Hg�vm��T�70���ќ��G��F��f�fM�+�݌ŗ4TM:�Sk���<���DD=�_���,Jlh�oj���_x"זּ������z�b>U� �]"��H�l3s�������3� {0�o����vݭ~B�է�U�mn&F�����=k���R�/������w�ǵY5*g^���={o��w&�]1�s�-[h�������.�f����_�U���Z�%���Q%!/����� ���CS&�'+�JM~���}�i�=8Q(���X��j�?�Q�k ��k���������{�\�V���!Θ`�(7�t�d,zB�.K�*$������M�L/��x����nLf
�M�")�:�4��������CqZ�,�x�W�����5��!�
@VPv�s|��l��9����I�~��S��3Bq.U�f^��uYI��c���)6_�f�����~�$ى��O�'mw=�^'�͏^?��ӆ�JoC�Ǳ�ط����̏HZ���/�r���FF�������47ۖ��0Y m�*Z�_�  &���[\]�>�r��|'�OO�C� �G***Z��СuZsWp�i�6�;��Ix6������O���@���g?���8 Zw��h�hni��Ǩ�q�Ψ���Ȱ�,\�DPmr3]���X��=���me�Mi���ʥm^��y��f���C���	t���<��ϧ����v�2�����Z=�a�.pB��>q722�I�p���qk�n(F�6��Hh��WP�?��I����F�����7��J>���~W�h7O�����
貹ڒ��78SE	�ڟ�~m�w�>������:�b�� ��=@zn�9o�`H������@��8TpLN�x�C�l{w���Mf�S(_�
aQ�O]�[[gR��)@;NS�G|�_����s|�+cff��Y��+�b�ً�a�HJ*�O�̖���Ex".���&��f��{�1x��_I��{gg�u /h!)a��N���E��b�3����kZHXD�a���C��H�~�.V]K�>z�Ea���i̷��M����wA��C1Z��VS�ܒ�u2K�P���,��A��A���������z�M�9z~�3"s+���F߳�f�ÿ�oN�7�����s]Ll�+T�|o��±�2eԵ�j55���C�6���{�ڟ����0������)�jk��/�p�� �s�XX�Z<[X\'@��@"3@�.��Y�~�!��`:=�O��q,���:���5��	|ʩ���z��ٹ���υ��*
���Ω��9�������@�#�����}#��g�B��ӑ�n�`�]���U���n�缶�D>Z��>h�����dч͠�є����+���A��sү_��z����t��7����-Qzƨ�&-@sM��HT���8�уQE�WF��]�N.����qѥe}�����G��v_��c��8��*p�X{�~���A�s�}y��S�2���LAGǟӞ��N��SBZ��Ԭ,�є����A�m��jB�BN������:/ �c�=V���O��7:��l*u_@Z��-��g� ����x��,�Hj�ѵ.&���������Z����Ә����DG�_	*7��]��Q�BCI��O�L���}S�����dj���r'�6B=���a�s��BmW���{�H��4_uuW}�_�\�Y��
�ȉbd ^�9u�K�޶Q�����~�����a`*�c�T����w��s�UW4�~s�֨��eU/����\�����cWh� �4\
����b��z��Uըc�a!{��kIy����/�mbnw/�u��jFF(}Lҵ���c�0��E��$`���-%�<��&V�Y�a=��m{CY��
�����}�5��n��o��	���(b��ppp�����$뉾Ťq�\��Q���n[%�燱��1�x=x_T\lX�b��l���ۅ��bz<_����t���-�S>O_��W��Yw����`/.*z�lt�UT��/z���p,�5����5��G���wII��P�9�Lk�Ԩ��1Tn���
����[[;s�W�ͽ�{��RRy��E�n�{�����˾.nb=3�����G'v�S(!!K�ݝvG���=I)ǲ���ݯ�d�ٕ��#��y{�\K�wk������5.���O�L&��ᣤ4!���'���(�跕�����o�9s�;���ȸO���ẗ9+h�ϖpl=�\�03���4����I=:B�D����j��oI���Z���i���G��������u�n�����Ks[1�xNg93�˯i,�%��Ś׋	!�F�;���'��u� I�|Xf0�b�l؞S��i��H�[��,e��������L���;ˮB@,��?�h^���U���u��\�������
PPQP�(P5 ,u�u�9}��l��y��x����i���?,KbnNyU6���\:���n|� �w�N�ձ]����C�+6cZ軗�!A%���QN����IM���0�(c:"��KgK�m�82��d*�(���U�xyI��l��tZ�)+#�;��gL���L��4�(�;<Na�����@������Ȋ��q��̤����t�
|De2il�SD#+�gи%8@���P��qfcS�a�A�,//�ed��cµ,�'V����g|���U��g���.��
{g�*ٖ+�$:���}"��?�|�W6���';��嫯|�k���̟�L����W��Fs���R�!w�)-M���~�X7���~�q�����?a�����2�����k��O~,^��j��4jޗ;L4�&2��9�����}����[�N��Ic��/��
�)bLN�~yeY##��݄��H����#��+��[��g����i2��A��H$J9��R{���9�����t����Jjj���6Ɵ��z�/�M`5ƞ(��VJ��6�GӸ)�S���͕���U�<����R�9������5��lm�XNJ��^a���T�}V��V��y�YC�G��+h���K�<߻%�논�ޜ�<j��7 ��}��U��%�h+-�/����培��o/6�yFJ�~?ub���b�hZ0��&qΏ`��&B�-�-Sx�m=� 	�K�W�:��Cz�\`�i�ݩ�}2>�|gNZ.�&vD���-���Kh[[��^+H��{�lyyْ*ܿI o_
��[�4n+H�`i
��� %#�êX�:�"	Mtmm�o�GGQǐ��L�+�I��c��|�D�$��-�l��J9�"����㣣��Y����lВ�;�0�kRR^z?(���_���`-�����i�'JG���~��R�x$�:����a����N함�΀�>J�[yE;L�g'2,��ص��_�����S� *�n3�Ї��I�c`6jg�^"ӯ�wZx^�a(��.1��>�YԬM]�Pغ�MK�8N������rgp4�������?�0���B�PTyFB&x]Xb%���B���/9+���R`�$))�\֜'��hε�ǭ��
�
��:�� �K\b"��[�hOj�^\��O�73=���G��G�%}g*I�>�!ǎGa��YYY+�ii��ff������9��t?QI�����*lvT[��O[6eG�뜄D��Π�{W���q�%��2b����y�}t�ΔD[OC;N8����Z���FH3�����|�c���d�fݠK^ln��|T��O����W�1@���Th��3��ګ��d�x?��\>~��%���!��}<,>�ϋ�k�xp�����X����Z�p0�1q�oz|�=n�򻆞�6�/���h���B����}L^QQq���Izhlr��RL^�祫��)��po=voO���`���&""�!އ�#GC��~��q���\\�\�굽��G������c��^hDV�*ȳ�1E��v�]3YY�Y�@�^u2$�L4�r�Qc��	kE� �ĩ\��Yz��z�{L��г��M��Wz��C��81	�e�~���K<Z�c�g�G%%��M!�HF>XQO�����Yye%�P�no�jv��axdd6�Zz���/M8y���Ƴ�+�#]�&��Y�x~�c8�E���݇!}/UI�K���q�32���0�Rl�c��J�	�@�����w@)U�q�G;Z3O�鑲��!�)2�%�>���Wm$D��,�_눉�����K}���y����F�!��x�g��6�ʖ3$zUU�AKQJ�&�/���m���dDD*:�.�*�_�;���3��Jfq�̘��c��I�9~��R�__�V�n��R��(�/!J�A�d૖����5������U�����T����d߫3�s2V%$�G*��4�\�t��5d�SY��z�`'������0�G�mp��A:C�C��F'�-�)m#�"ǉ���74$����3kӌ>M��ә��=�百�F�i}�;g����?;�!�����~�}������FV����ғBz�7T�/���0ؐx��;�^���i˘)�Y�Y�{���;FkM��G�0���jEE��rS��^��Ӛ��Q,��+tP7���ܹyy}�6d4��1|�!�dW���ē͐��UU�������1�NF=�C-?��坜�i�qp�{_���)��p����Th�q%�&$�s��5wt��f7|3��m�JԬB63��G�+k���@:Q#$DL���?�����(o������ke  �����R����L.�heE�VI��L�q���o�����B}Ĝ�9�UH��2p�	�@�=��x�z��G�ܑ�T�]�r��#/�f�}��i�x�yQ���k��$[2cf��xn��Ջז�oO�@��Z��@��� �y��8�	�����e����H�ˆ�)���y�,�x}}ee[��A�Õ��H���	>����y�)�Lעt٬�؎�A!<ԯ��5tuu����⫝̸#�����@�ӤW�؏�@-�Rg��W���CRK�q���K�j�{���%�"#2BǄe�I��.�)
2�ܦ��
;ʂ5Aa[L��st@�:Q*����# �� ��3���x�HI������ݻ���������<�޿	I@i��ݐ�����6��j�4��4|�i���Ǩ����4۴�B��dk��f�L?�>�Od�j  ��H�p���ݖ�B^y2��\�L�\��1��� �@tӇ\���J\E�
9�
j��>ǹ� �Y�*Hcv�"�H� ���>�T(�n%��R���8���+�.ݮ������˗<:�*�kL�6�"uoz�x�;8]�����W�o	$M�@��L)�Miǀ1E"3a�~3
�f9R:*1�6�yE��S1����I`Q���Y�<j�}�����hh����	�oH�H6վ���BӪp%�oK��A���_�,Y���2��p(a�	0�$45目hD��6!��D0�qlXp� ���_�g]]]Vt�<rF,3�C�OO?����A�d?͢��?��`�֟�:O��tuy�w/bU4��L9b���y�/��ɰ��3���cZC����'��}�2��ܔԷ��n8ܧff0��۩�4����[=��8�1�1I�n�N7,��M��_���tu<dZ�GEk���0xw4�Ga.&�^��E�����o�C�|98>��(rx�5��˕R����^�K˓n�X�ki���*�/Ξ�1�^��R�����P��1�-Kee�+���;�C{5,R_:<_��p�vC"`7$S��,�5 A���N���\\Q��:��􇆆
�g�\��q{���.n#��(�yn b[MYI��~>,��>w޾=�϶lӅ���)\KKK��K-�١p�z���Im�T��S_�.,��蝱�˦ט��mڴo�7c��v��]CS������A�p�������n��tέ<׋fmH���_��~x��ޝ�}�:�ԋNJ�:777��r���`9C��(�p?W]v�m1�֯��J�R�@�;��`��^�\�Bs9����Mқ���: �������ftPhh��GH
�̏��e�v#���h�����-���D�డ�CD ��#��oZ�T0��@&�����o��E�hQPeIP���g%�JI���PK   ���X0jF6'� �� /   images/6462d580-1c26-43d5-8ea3-52797bde3c40.png��eX\Q�-HB� i���w	���www���5�	��h�]�}��;ofޏ��>{�U�j�:ݧ#>+I�! ������H������{!!�̌�Y�|�x� ������z�N��,+!��>��H�uw�5���9�$�TB����bdlH�<�^�H�sL]����ho)K�5�������cf����1ŐJ7=�g�OWu�χݏ��ekB����E^��Vr>L?tz�=�)F�E�!���$�yV�E�(�Ʈv��p�����2y��o��?r��|�ܿ^H� M_�H��ua�k�U�C��S���Gʃ#o�#����sa@E��}G%I3�����O���ֿ�E�/�#֑u#qaA�;�FrE��E�C���p$o>�����j&���Y��Ѹ&u�u�̀S�5;>���9 ���z��Fg��'��(�C���:�����:������@���!���{d�Ve@���
Ζa��6�謇���&q%U���"oG����H����^�ǰ�h�Hf�Mbp%�o[�������_�/�@VnU/д/��
�_��KS�g�'�?�p��2���.nR�xC���Zauc!��E��/�a�ϧ�o>��t��w'JVim�M���M�̤�Xʣ�G��:?W��a4��*����Y�yQ���������a;�z��r��@5��C��|FPh�����V�����h�?��_�r�I�["+�
��/Q����#]���DEFDN���J"�:�z�Ё���>�#R��R���*4���/��D����Th^C�aq��C�[=�_R�m���c����Ft�@�����o�Bขރ����FX��?�����̪��o!:M�p�D|��6i �u<��C��f���;.�n��zD�\D�/�D�^���w��ۗ�_ܽ���fp�^�#�E<}��+*���O�%��f��k�R���Vf�[��[U_Ym��#H�B���a�������H�C�}���|b��F%��k��}�ZG~I��wJ�}�*$6��9����ߊ8",>�������w�̗_�x6�׽"����g�U,���ț�����3�����ۿ�xȾTqd�o��q��G�_�~�x�vU�f�Q2�E)>!�hƐ��b�=�JV�_k^x���/ˇ�_Ѕ/X)Ǣ��k��+!:��;=UZ�r�Dn���y���e1����	6"�� ��u�w���T�2����P�"(F��L��l��%�)���B���q��DKM�3�cK$���*�u�?xe���(��Rm���]��e�����?�(��w9,X4��ؔ�W`U�eФ�ʕ�U
��i࿰$�uU|��y�� ��|�2�3���2�M�ݽ����O*:G��#na?���c ��u�Z�;ƿ�p��c�X��7^IO���g��׏�<>������A�]�cE���z��P��6�cˤ�.��_P���'ϡ�$���W1������ی�g�:��֝��_�+b��Ͼٛv����/x��	��������`�&�%b_���%�In"�/T3����݇��"�p����,+�V��E���������#���c^����\�SR�~��6~~iu�S�텠������OHd���[��|�U�W�^�����ֻ�?��g�1��n]s�F�^�oV[ag��N�����>|�MW8��]�_����0�9HO5w��Xg�~NU*�����6���e�Xz�*ɜ)��FV�V��`o�5�8�S\v��L�NFCH>̝;�gJ�Ն��&��:	C]�!^����I�����,|���̇�7�H_��ݢ;��G�H4פ�l52�]`�b:	"���[$ǫ8��	�����!bKd�p�8}ũ,��:�u�Rg���Y���S�ۊ��VUJ��/�<B��/()f���a���[�M��1��+2��� R����n(Z�Ò�>\�P��u�}��T�g�+��f*RC��Ck�$� ��P��eǇh����>�'�젝>~K5��UdjI�՘��T�<?[C����fk>��UfTѪJ��]������N��3�>6���i��E�66���|�6؍�5:"K�����jn�aZf��.�����gQj0�ʇ�� E��p,�R�R�$CS֍GS��dϗ��ܐ/�[�z8�-�L�|���p�ĶK$J{�g��1bE�'���r���7,,�G����В��W����5��5G������֯�_w�A6ZZL{�'C�&��,��ZG���v7
xK8�,�����'F��>�љ��yNð��LTB���x�6�듂�dcv�<�}hz���ё�eW��%rY��x�X�Y����y���$��]�#�"Y|KOr�SQ���զ��g��ll�`��*j�j�Kƍ�<N6QQg^ 䐊*������5�'�b^�!e)�M��J�Q�-7=�2�ڙ����*���#g:�0(=�S��'���+8�x��.��661?�������fm��Q�̙=��U��çD1ȒRG�V$�!�� [>{9����LC
������2�&+anj�ڼ'���t=9+��l�,���r/�N�φ�������/_���ܔ76������5!,�o��]e��6&��Eڈ4|�~���0ř��Q5���+d�E�N<�߲�4�}����&���ZD���Z�[6����x6�AJS�:AګH�E�%�g6�vF|��;ס��1̼��g�M��E��ܶ�n���ܠ�E3�ʭ:���{⦉��T4KC��W�m�?�,xN�2��F���}�C�*hX|�v=Y}+�?����,:$Wᓇ[Fn�B`�R,��*��Ϲ=5���x�������T��2aг�F��`�Ԭ�lD�e҆V|�DJ]�/��"���Y����HF�aC��S�N�@����:��/G4�u-Q{�l[�5߉f���j�N����X�/
��,�}b3�_�v��	w��"}�p�l9E�Q�ӓࢢ�>�$���V$\�%~@�����ՠE'�P�������H���Mcbc��X��`��m�w�r7Xኔ"�σ�����4<"�H�wp���R��9��"�2j�ìE����(iQ&��}� �?S��f��l.����G~+��VmA�V�D	7r�R����JE��<r��3��R���u�Q��I�| 'jG�N�H��=MC]H���'z'��i�B�o��N��Pj�w�*�(�$/�7+lB�ʤ����(�kt��6(uL�5����SF�T��r#1(\�d�,�x���vkb/]i�A���BE�J#�CW/P�����h������}#%e Z�9�#�+~3�BÝ� Y���͓��ם��Enasr��&@�zRϖA�6.���@a���Λ��?V����g�W+N�U�h|�f$�'ڴ����ue��ɀ3j��@��>��)'� ��)�=��ti��[k29tQ�O����R=ݨ�{M���8t�N�� j.�o��	ҫ������+O��nG]6 f{��=�赳O�CR�7ſ�AG�*�p��<P�>CCD8�����׊�5��<�ZVlNڀx���i�<�ޞ1 .PrZ��W5������pim��)��(�0�p����5s^�۩�(�R�+��_�&j��l1���O��1�Tc�K��8��LS@o]-è��1}+�^-1_���ƿ0%� �G(�A#�<�����$�ļ]����q������u%?H��nF6�c(�p�m�ם��Qxk���6��_�N��h�S�#��8p��~#�@�Vت~h(iR��c}��:����T�҅9g�|
�٧_+��3��⏲�� 	�&���LF�3~嘛,.x#&r"�tO��҄�O��9�`�4�6ƕ����{g����*��
����_�^�ۚ珵.������j�"�d���|��@D��1F�5�xT�:i���*��x��p�[w�����-/$#�����@4B�g&�{��w1�^����ժ�������mz������u܋��w�T�}O�7[�ښV�6�y�ε0�����+^��&ۋJ@q�~2S���|�qI'��X	�d�_2�Qm�~ѕ�H��!`�H%���
2�ҷp�<�7�`���A�1���ӊ3��M�f9�!#����"�>D��Ď|�Qo>\�ǒB���Á�A36f-8���E���SFZ�_2��/����Q��� �VhH��ZXξ��0I0�������c��b�`%��(���+��� �i�BU⪒�F���O7Ě@K{��ú��̶��͆x��'0S[x�J
��rcǄ�w8ɼO��A6�%�n���0����8��e����1K��yp�l�x��a�B��=�[M_��ۯ�B���T��&�{�>�K/�U2\>�G<3#ĉC�����UE�6Ȝz<5�+ہ�����`J��(HU�H����� �]�er�fop�5R%���0m�9[��G'�O*S�<���ۍ��*g��	Μ�i��X��Y;Ӗ���Xt�u����e�KiC+��5 ;t��^��dj>Y��+�͉��3/D\�$����(J����/�������c��#D����Ѿ*)t}�&����#�3�M����|2CO@��j"\3Ÿ !�l��V��";��p��e%cy�sFe�������F�{'l��Z��@~I�ZD�4&���,�KO��d�y/ŋ�P��B�������<�L�<!��4 �ԙ�B�)p��ؕ&_,\�n�$�d��9Q�|�Urr��Pec��덝s(�9v��|��� �Q�E ��ܠ(t�B"q�ϩS�ы�&�3e0%cC��?6���Q�cnSڈ��E�I��t��y	�,� �@���C��0W�8�Z�����ӻf����h���z�~�����`&�~Bl���J�LKX'X�/D�5B�f�4X$/���	�+W�/�Ϯ��g U�W��}yՓ���ag���Ļ�Qϻq�s���Í&���`~��*L�'����M]��d�ǌ�K�q׼���:���)�FfR�C���Ik?&A������{�����3���[�ڤ��5R��v?�>�$7௢��_a��_t�+I�|
c*8�l|,���Q��W%��WA�2Jeb�o���=Xކ&�B��çҦ��lu�L�P}��o<p��.�{�.�!r�F>����,�:�����D��n��s�[&U��)@��B^x`����0d�����Ɨ�2x�]d��z��y�ۮ��Û�0���K|,.�";b�S�|W�Ǳg���"�G|J�:l� =��|�.�x�R	��/�xE9ـB�Se�/���Ⴙ*���,�ͤ��R�w.��p�r1;�x������(Ѿ�q�Ea�}�spB��]�@L�J�����A-f���/��0z�GN��<��� l��E��d�B�����.�;c"�d��U=�a9�3�9�B�*ؒ��=����8~F��9A��ճ>P�nx
�ҳ�T��3F��ؕA���25�L�� ڠ�f4�@�~'J%�ƙH�>�*	���md�'��=��<@�G~� g,LD#���F,]QR9c�+��g��D��M"4y˅\�[�`�Yf��z�#� �`��M���PA�L��P�4� ��m�\��h�!��pFGS�w���z�D"��D�`�$l`�l�	��_�G$0̗-�����p%�:r咜("E2�ɶā�6�|��<�
� I"c���t�u�*ֵ�SH���S���4h�05��\��o:�A���K8U��ï��uf�S���T�Eᯋ���00~D_����	�!�c/
�u�bE/�T�.������]2�����
���j���r5�(�6��kt%2	�%���A,��/J��)5!"(<[�r5�����D�Gi��834�Y�/�����ip
�w�����ӂ�#�Ͱ%~�l�D���ʄz�ƗB��듟�-2��E�YbG�R�õj��Fׁ*e
l�X��P�ͪ�ԛ���%>�`�<O�����n��:�˨�
���l��2�D!�^ ����ŷ�oG�$�f/}S-�bǝ� ��_�@H�����ɉ�Y���Aa���Ҍ���{a���}�$o�	�'&��mY�t�3��O���mM�Ra����ǾQU�,9���Z�ݐj�}j'�/Wtua�v�-��v\�?:R>:V���u�T��� -D�������JR�D|(ȭ���D�4�}%�r�Cp�g�l'���t�ł�C�<��|�%���_B$��z��[@Hxl|�`�ۚE2+���)sH���^������h'[��j^��'�
c=t�Q��{>����Bl���N����0�� d�}Y�(DH.�9�"� �짡�d�q�w�Dx��� V%�n��<[�3�zk�*�,b&�1�DG�w
�r����*�	�.�K최�Ұ�z:^� ��ә���ܵ*h�Y77r�4���R���)U�Ʋs�ɖ}����)p�ɀ.��M\�~�Fk��zqN�M�M��K]7��#}�I;.e�A�����u\yo<�Z!}���~�+;iPe�w���iÃ�Og�.�����)�$�gj�@�4�+*Fe��������>���B�J�Z� ��q���p���juX5vؐ�{�\|�6���c|b�ؐ1	��%0�}�	�HUHs�,p&D��7IH�Q���c����&�_D>{��ޣ@��s��n���/�Dpix���]�v4
b��$�oV)���h�sY6��}7�+/��[�K�6���%������D��-�K�8�AM�1#�v�d�r|�=pu3V�b����iC��-��PY�Շ��+��WG��b�Y;G�x�f�1A*�����h�x���{��3n�J�y�f=n�Zj^��eJ����x5Kj:ĕ���=
�Ǎ67k�ëlRU�&N�~�������^��H�o���T�j�A����[+	1�X��̙V�v���s$��U�E+�w�b�0(����>��i�2�8��D�a�w���B��o6���O{jC�M@"c��r�&'�G��o�&�=�`�!�\UBA��X���׈Y�:ڡ�vQ����;�G�䁺N�{P��
ry���O{�����;�$饈��H��#�z���$�G?�������ܹ���phAH��Қ�^�f�(���ɡf��R����4��Ct�-p"���ثP��1w �s~nBQ�k��ay_��֍kc������MH�i�w�q��Ȓ�p������i�U�G�뎬X.~�7"<��[�i�]G�� (�]ت3����I���sT^����q@� e�{�%��I���j,"!)DK��U����H�~o��M����C�2&�Si��ǅ�VNi�J�l�P�ܲ��;_��6Y��T!��x��E�@��VՁ+��}����[Tv��?ƿWa�l,�-����X�~���^�ѱ{�<sU��᳡�d��(S �o�ڰ�_{�|+h����6���-����ui}qЏ�X���d�;����qd��S�O���_;J�u2�����H�Q��lZ�g��.��g���OJ�x.�~����(dQ �Bh@�\�S��"1	�`�奫��V�9��_lk>�Gv'-)�OB�"���FUL#%�۫<M!(�׿�l�PD��D_
/~u>��8簒�"U�#����~	by�욗����o��,���Ŋ	Z;�Sֈ���0o'�es5�]��[TD
��ؿ2�<c撌`���E�9E�����+�_uCQ�-� �Uk��i]g� N����u�C�H訅��nw!y����ԼVir�iݹ�L:A��e��e4}
5����Y-�﹵�j�h�p\�^oȵ�$���R*������Ρq	��Ø���>�b`j����S�z�?@[�L`�Gg��ͰN�(�ʽ���eS>.���<KU0��WD)p�f7W��r0 ��Vhx�(�u�3�C��J�b02��Bd�ޟ�N<Jj]IoK"lqI�jw�Έ|.J��WE9m	�t=H�`��ټ�,�J�{��׼��[f	P�;۰'���A�'��lw@���k3��b��Fr��t�R[N9M�����BD��OE��&i �������4�3_Kpi^�����3V������Vq)��sB7D��vQ)����,=�Y1�
��(��+����ʍ%�w��{,`Z	k���3��3F ���%�~�����XP5����d�(=�7&}�l�MΥ�f4Xx�9M�b���&�9!�o(�
Mw-7��B���h6&�_�o���^q#����c��_/N(P�E(
#��a�S�Z�P�����'�H���\O�;ϧ-�f�
��hh��;���w�ޔc��#���H���[=�*C2.~���v��ל�u�4~@҆{�]�N	w>�]�X�c�̟k/���=KbM��'މ�;�efTE��������D�G��̴�4�+f(��J����7��|�����s�oY�fHL�Qlˡ���U��%h��[]r�!?c� �v-���F1�&Q�)3s�����.�W���<w�ae�B�t�s�iA��J��˝Z�2\�z�4��o㜨�ۘ�t�J).Ɯk���2��s��A����Z{q?�KO��,=���"(���o�P(CA��.'�'?<C��|>ABX�A�� �;wɎ�b�j���^;�p�
����wK5C1�:~��Ge@}�;2>�?l��d������j9&��|Z1�`�F������T}F�e��c'�XPN9�[;U���}��}M6HI�,�.�*)��Ģ�
��M1��4kx�5�.����)��;�)N�AصͶ�>�p'M�aF�Z�N	��vG�����ƌIi^X�Y��كן���H�~�,b�i�6q|��C�����P�|�'�ȫ�nf�G�ֆ����4�Ȼ�0���	��tR'�$�hDp�������ťn��j$�b��xhR�8�w�~m�]K�'r���w�e������:��E)f�]�L�
�6���� �i�FT�P�]0V��yVb�i�x�Q���=������{ e
3<��;�y/|xp0�O����h����MO'R�WVU��̕�I���=���6��j�\��3 �k.����He3�^M���K)oxf�[�:��G�r�L>��Jtn\OH����Y����цZdh p_�D'P��,�m�Q��ϱ6� ;��#. a��L��h_!�H���1"r�!܋��q$;�%o�#*
P����.>�v�[̲����VQZ"ۜ�W���J觟Ȣ7K�I�b�#� �.�����X>Ohm�i���I3�-ʹ(�U���Z�b�F{`�1���R��n�HM��㌊ɹ��N*��2]3-�T��`��X�gzJ-��?R�
����s��K�&6h'l�Ӷ�2�Sl$H�=F���qo:�ǻ}��C��.kZl��C-i�ߡ[F�� �Q�/y�!���;�&=7J<�j�v�U��g�J�澦L 9���4<�tJU@LLXs�)�������H����O��[��f|����am��ݧ�ڃ�'�X_���\~� %=���*p{��<��1 Ѡy2mC�L��0q��	��װW�q��������Tͬ.��-Z�n{?{�I_J�TUV�����Hx�)g��f��=�ZWhjf&��QlD1��m�������5�2��r�z����y�h�Ay�r���6k%˴%qV��^����	+�\��i�E�ئ����1dt�(���s�,�K�(�����vfG\nvа���V��j���s����78��vڶb(ߍ3�2bi@ؚF�c����F�9`^�]��m�{��e&�O �W_
ߏPQ�P�C�x�}��g�ɅJ�F�0+����rV�"��~�F�2�Y��B0qO���b!�;3An��V�iL}/�(���ߺ����WA,�QP�ꏨ�@�Xz��Azj́���qO-������P���2�l�h*v��������Vv�CZ1_\�9£��6�5�B
�1.v�)|O��w ���J�R��RJm����+O�i��03�cz�7��#h�t����E��t��n{�h]�7�|.�[���a�aE�0�A�+��%f^JD����+B��#�2�E�j@��ۑ�� ᾵���.����~�^z��f�M��ٟH�����-�xI4n�p,�>��)]�G*��N���-0P����'&�M�k������U��w3�c���U���C-k���G�Q�)�wL��o��&�fBV?�UI��l��n^�p����K���՟Ԭ��s.�V�X�v���gC�B��̭.��/4�O?^����)w!QQ�b�t�fͱ�ƺ��S(�1��{={�!�:[�<h�ƕ�	tm0a`@p�۶�*�=ן�����W�4�2u�
~g�ޫ$l�aD�m�VK��6���Wv��5+<>�!�S�%��<5)�͔����T��� Jia��P���c�l�vF�`X���6߳���C�4l�U�C���z��O��lvt���TS�[1�I$X�H �@�ctD̏�����Z=IL0I�k�H"��o]'�;�kУ��ǋކ������u�n��BPS9��W!|�J͒�Yd��bI�4D���#n���=V|�@��zQ�i�K_���y0B�lG�p�*� �D"���[;sD�|��t��C�w��m�gw����@!��S8J�)�V�G��'���!Dr�Ȧ{�����'� g��h^^J��K��v9�<3����;��T/:'T]��@��l_	�"2u�c���3CKd��Z��
�>�~oTbq.U��U��$�_�6l�1n-�c��э�Kˌ8�z���=�"wU����AKt����5��C~��ua���|�/�ݿ FR��M`�ƣt�K?�i�_R� n�$��]f�>��:�33������?7�������S�15����|��!��pִ��W����FOY��fX��{=������<��$��y�E��[L�Ⰱv���q��t����$���aD�x~�٨�Y栭���\K�㉫�#�]L�z�&��8�=?��n�{��}�?���#�=j&���j��1D���gb1��Q�D�ɛ�$��6�[D�$�\3�{��k�����*;�k�ۦ�*���&�F�Ǩ������$���	��ai����o� ���Χ:���}a�ML�{��xA(��r�׆�����_/�1�����-�������%����a��-.��!�E��SkB[���x�V�NV�����;S����FW�i�,������f�I\� E�K�~��Y+��y@'�IhID�6@��P����K��Ħ�$k]2�����SV̕�t�������X��g�O��y�<0������8��W�Z3/�(�:#綿=��-s4�O�T�|"TTLcgY�m��y��hc*���Հ�\�*zg(����iL�L� >W��r�)Jʁ��\� ���&������J�R���������Ў��y��ΨGJ�|2��+r�y(�b(�j%��P�O'A	����Z�RfnX��� ���P\���
趃���b���v��< z���$ b뾲��x��9��o�%�������ME �	������}��<
�"D�YR�V-����0�[�`ۧVي�$��.�3���6#�	.�zc����������)/'d{�2��p�T�
���)�ɯ�߼|�3'�i��T���,VɛP�vE������s���x���	��Hne�D�{�SK��xn���S2Qˁ۠�ܘ*�͕�&����c�����	���O
8�g�
?���;k�}�R������ ^#�e.:����>�a�ꪒu���4@���G�__=YŦG@�	R����Do6��qJ�˵$2���1�_�Ȟfd���O��Uj�4V�"�(�R�ySw�_��=�n���X*U9+K+���9�Q��4_�N��\����PL��	ߖ)�hv��e#ฬՑ�]Y�ܑ	�\��$mյU�?�}�@$of��aè��j�sT��?�D�(v��X� �B��̐�^Je?kw�ƛ�%�����D6����dms��G�5 ��+��ӯL�s���1��
�p)L��K=ј}I������D�v5����؄�}x�'��q>-��D�s�N�"!�2�o�$rc"�>�`���o���Gi�I�iQ_:��G���Y�/��%��sI�GޠX��C��[�M��X''�C�e�j��)Q�M:���-~ʽ̴.˪���7��Ƿ��1������;ޓ���z���W^���Qk�1��?��!%:��^t�M���^�&���v^���\r�9��/�C���EAt���r\�B) Ǭ�,�ؗ��r��m�-JP-t)p����~�����ӵk��]f��T�1�q|��]5"���0n:��_#0��n�y���'=W�+�	�Y�o�y����ECT�uG���A��s�)ߕ��*S��5����Ub��DE��v]� ���3��3I�	c;�R�
�u:\��\[e����L-�Z� �#��T�e쏩��āUƝ��N�`� t�P���'W;�"~�%�}*�6�0�\⻾�6~��9��y��1���1�j��1��F:��V��dM�2x�c+�O�	⢶��:_�4u�+�"�� �=��o�|nJu���2ʦ2�a;e�rc��{Μ���^\&r�m}�+EL(�ƫ��)'\�`=�:�D�U��n�,����5})ǀ2��.t)]>�7��}	Ehـ4#2W�T�X���8�ӶM7w	�	��rF��p�G��A���ݮ� 33�\�-��ޫ�_�J4�o�:����z�����yl�X��nI*+*'�q�.*+���
���I���7�.���K�|r�n�$�U��������W���˒qq[i|�ٻ���4��AH����xf���^c<�k1/ז섯��<R�-�mՓrL��,G�[�_��I�Y(XK)��0NzV�# ��9m}*5;l��>��6%}�Yl�-~���z���w�7�|E����/,�>���p���"��'��Aj���#�b�1������u×VЭ~�Yˍ�)s^Ҁ4�a�u�g���D�g��2'���5�/?��	ʙ��'��Q�c�D�mT����qk��I��wDB�
Ca��0:�<olvZ.��&����21��������)��Y����n���m����|���Q߬K#$�w
�,WACŁ��da :��_(��������;)y䓯n��I��}�0ݬ1V� Z��&e_k����λX�@��(���tӭH�F�Y�5y�!H����֒��_�2��z&�)���M��4�����G��ew��6�Dk�C�+)IO	c���"���ǳ�&GE����-U����*�q�ى� ޻Wo�#ݰI�#2��| �{���	%�*V=�1�lцlvҬ�A%&����$,��VAz��Ԝ�N1di����'$5Yf���:h�of
Eյ�j�m0B�50��1"&/W0���.�Mm�S��]u�ˁx��ᬸ^���-e���L+V��tȣ^A���i����_5��++D�hw�� �R�;�K���6� �z���Y�hL��ܬ3��=����w�l5�j����oy��]ߣ��I��.:���*�C�Η�[��x����Ui= ɬ���v�԰�4j��@e�Zǯ�;tK��㚋D�+�B�7�=#�.v�4�g��'.H�R��utr�����a"(�AV�<4MK:8��L��NO��1)��o�Ni�O;�W�G��l|�gL��
=���OԞN}��H�~�qS�]L-��O���D{1j��@�~��G��l^g�{꒼�}E����W+0�]�땐��A���EE&"��v�D���XC��Q(�G���4RPR��f
u���~��G�y�/=�����iMe����G<'M��\1������jC8�����J�ů�E�D	fIF=�0iHιUjBrs�� �v��k����.BӉJ�X�^�I�cU�����e"[a��s�ɤec��0)�Gzl~2��B�C�n�a�,�|W�P�=�EK=�x�p���2,�NA���P1k)�i@/?���hv5���+�>Y2�+��q-����952��f������]���0������������2t�룿N��VA��X�)G@�Zjz\�*t�*j����� �fꌐ߆`
��( m@O�]!�:hAp���=��d����+J�k?�{�f��X���A�;j�O���<A��Q�&s�ۓ0�0t�B�0��+<[~��Q���ܵ�����[��X���P�O:��	~�
ۑܝ?�4r�y���N[cVs�Q��^Ŀ_�gl�B��7�m�og\��3Ƚ�:BԬ���Z�{L�e!:�DʇaVh�XTS��mI
.2[~q�u���eF�'w�!��+�p2�Z�Θ�9P�����Vd͚���7�;&���_��-B��F����}�:��c�o/a��Y�(M�`���Y�7�>�z�߅�U�
�xDE�5�s$+�6䢢ݛ!�nB'#a`:��z��÷ ?d�&�_d	��\���gʾG�.�9�2�o4�6�}�JY�'D.�>z>|�\�h�a�8e����<
��L����)�zڴr,�L��F6 �U#�h��9n���k�iث�q�ڈ���,!�^ v��:�ˏ���m�ٕ���%�� �n��o�'*X�ﱺ�z�@8�6���?��l��d�=��=~7�n�A��[cʜ�om��\�o�b�{���@�CA���iKl�z ����l�ՊJwP�.E�VSc�G.�e3r,S�O�����\ٝ&.�ԎEG�:Q7&t�3F��cB�[_O_�+8j.S��\���կG�6�z�˹� ��H����q�̴vE�"�R'6M<^��0�\G�uj�T��>������>�-:��~52�E��]�N��j�&��YZU�R��V���D��wPHӆ���۷l�oZu[7���J���G���D���,N���>�|�86�r/���8q�u��� ��)i�[ڽ��}�O��0�Yv\b����,��+�r�ZW��|vNs�����k�L�w���nՌ 9�Q\��Z�Ͽϵ����@����cF��}�
�Rjx	)l�*�e��:�L��T|Ud[�gn�C�]�Y:BA�Kz-.	�>��^��06�M�����3]Rs�U����N,�s3@~��^�D�a}�.���e����	���|Ҋa�kk"\�!i����;��Q�ƖM�hd����m����q���XOP�[p���`�TR[ݖ�0DQ��'�S�Z�q���["(�ӜuJ�����X��j�9�a˲����x	ի�%t��j��7+q�Ͽ�Ͼ3��ا.G��7�a�z�=K�	�?�:e��J8&�jN��o��	���2/-��?����k.�>jy��~�̸��-����x<��#ҳ����MAe2��Z�с:��!������X�nU�ڑ��Q�1;̜"���u+>[r~���:{�<��34~�|��O��-��{>��d���	���dHc�,�����(/��l��mXմ��w��cTT��� ��.�C.?���k�0�����dL�-�R��{�n���KS�؏�E1������6�?3��&���������L���x�����W���r���q�����8I�n����h�Q�=oj�=��MT�/��F����'�c%��~}X]���$"F�F�\��L)�kW�0֙�u�O�JzL��&��ጵ�����d���)�-[.�b�Xh��j]JZc��ah�Ճ�MWyw :8���Ea뮣���zn�S����)p6
X�n@�6��\�(�%�^.�raJ"�8�'�����i�]'��i�v�q��, Ի�N���`���3�������P� ���'k��������d��]��~��	�r���_p����&���zp��@��ґgi��O���}��i#{��Z�ȃ�r��;U�Ϙ�=o�=�0\WO+�]�z^+� p��`-��@D�oY�KE�aɟ��AoÚ���+d�.�do8��[2�v�~��vU����K�bd%� �qV��G7�����8���ZY�=͘?�6	v\�po�	P�&�g�����,]|��`����y|�^�1-d��1�l�&���*t>�y�~�r7C�iQ
�����B�<gbx�e":�Үg6Z���5�"1TWO����=�%�.N�Έ�A�f���L$�/�V�.ȫ)����վ�6'�l�M�M�&> ����Q�V�yyԒ��G36@���;\��'?�A��σ�[}�ԞW=-[�c� 7@ȿ�枓�[��?w����gj��$�0^�Ө��U�,z���@Պ�����w'e��I��t�U%Kc+�S���zi0�� V8�9����:7���+��|��SZ�P�r�ٹ�)��!��K����lѹ��hnzF���Ӏ��Y��^�BZ�ȵ�C�`�.ի��)<�6��g����ѠG����U���bW�b���6���o��0�5�:Ä�Ʒ��!�)-/�C7��N��+�n�K��E*�)�]�إ�>���)V�p�ld�$<Ǜ�Q�P'��p��6N�:�����d7��r-g�_�Y����Qg�E}�;�:{�2�:~wS�isB����5z�l�����E����Mwѩ3�e{ٍvW�F�YH;�k�lt��di�����%������쮫�D���0_��\d=*����>=�s��rU�8�����t��jL5em���2��D��qј�;�/��<�{=0��8���c0�%�5�����~�c?I[/[�ă�@�a�ѯ���Шզ/�~�V�fjx[��4y^��N8:��	���O�~�Ԥ��)*�;��Ex[R�R��x��O��P�F���J�\�s;t"��:��I��T����?'�q_z䙳t�ϸ9#���S�{0��z�-��y�ꁪT4<��S��ա�T�
��]�ђR)���?�tx���5s�c�)Hy�5.���Q�Xk�g�gCJd�c��aO�u��*�#�|_���������5o��{�suN:�yny^�0�xj��6����QPl�k�4;;+���HS��s�W���`�4:Hʞs�ı����ѣq�M��o�wc��q巿����3��Y5+Ӹ�^���s�GʞB}�0r۶d7	1�K���E�Ȥ��C�gW�ys��V/]ϜC�ͩ:�+5ts�b�wg���moҵk���j����v�%�����QOڑ��8�hDQ�E�ҲT��ݤ����j�ӥ�v3���y��f8�cɢmA4�_X�����!��~��eI~j� 	�M�y߻���8�|�~�z��}��Ǩ�%�3��8Y-��=%�&Ɖ}����@K���'߁@p/�|��i�k�vii��fM�QG��祀n/��|��%a.�J�n}���{������<@Ϝ:��d�^�����|�K��[Tl����:Up�ݝ���䶷�y����Yߒ��S�L�F?>��=v�q�����l���=w�1�����Oȶ�%�o���a���M�٧+�� c�D;���T졲+����8˜C��|~���K���o��F��G?BUxx>~���_�\ŵ���񿣅�A����G��u:���wx��%0��v.�f͹)����4�]�(���4�NOK�딥b�������y/?�H�r�źnx�<M2��QLa�.�jN_Z����Svp��lđ	����Q	�,�H���c?��F'9)sǜ�m9�LQ�i(K�Ö$��W�Ξm���C^*B����T$��!�t\u������Gʛev��P[
�Q8�{ڧ��5�������яR��ag�wF������'���R�����*/S�)�|�/�ȍ�de ߃a�.//����K���/_�A��o�g$��y����T���e�Cxt�cō41%�ǃA�5�td�5��Z��
Hi��1h�����Ry ��av���`A�*^�o���Û��Y�V�O^�Og��j[����A^ȉg�	T��^��pD%��yi�#�e%\�|w��hc�C����x��b�s�����Q��8}�#�H�.o��j�^��B������J!*%N��JjI����DY�#�g��a�ڑ=�Y��$W馛N�^m��7c��k�s����s��y��s.����gnY�o�bXouţ,񴤙��o��s�k���],��0�r�����a����'v�]D]�r	C�|�)����l8^��#C��A?��&�zӭ��z��!�ۭ����ʇ�/���W�Sĕ��q�<)C׽�L6�-��Yp9��ɇ�)���g����O?K�?�$���]x�1�o��>��{i�i�|�A��/P�n����K������ҵ2�{�5D�'>��η�m��ի&5�uZ=�Bm��� J.�[�A��(��q�r�xB;��3����
��4^�/�s9��/[&��h�Wd˳dq���O#;��M�y�*������ך0"� hy5Y:�1x_w6>�ݥ��maer���X̯��n�Kߚ�,S�֍�t�w����Z�D4t�wთn�\S!�J�=�Z��w��O�ԋyٚO�w��8׋ql������^x趔���p��¡?{����~�n��b��������:�t�n>qS��#O/ؖ#�v�N_�x U�lX�]��
<�Mx��^޵��M�;��{����ڻEY8�&b���!�͢^D�3��-�Cbq�@f�*�$�"�.	���&���=)�K��o.�,�+Oyc�+�A>fA��%[���^΅�M����h�ۡu�me�W���(�<�܇��A,,�u1^i�j�5��di���[�(ʕ�'eKԳ��`��\�#�z��
)����x'�
�=�!�ɦ;�b�K�\.��ބ��Q����N
!��N�*�y�5�<����m���N�]l�qAW����3��]�6[�",�웲�M(�e�ه� �5h%�ԙ�[�2�s(B��I��>h��k��m�dn���8t����l8�z.K�8Ϣ�K�8��F��$��da�0yo}C�{�$GĲ�M�m��p�s�<��8����C�"����n?q��;����#Ϻ��,���n���y!�p���ԥ�O��|U�_l��8��%���y��*�REB^nz��m�<C�ؤ���3�߀7'�
qN�N>�hЇ C/)���>r�Z�.��!-���"�1�*�s5X�Mx�<�Qr�*|YK�!G���\;G
����σ*�^	I��ԑ@�g����s1�2O�igԺ�-�`,_�����μ�
)��=#���W9���x�I&����!���)�1���h�v�.<�$�lo���r�83w�X��ٴ��X�2'W�ˀ��S#	���Yv��������򀮜�@�(-v����J^Ev�dN�xk�Td�S� ��؞$�񀹻��q}k��K����ᎌϼ֙��6Dhmc��Cx�\��;���1�dy[ϥ��6U�S�spGQL�:N����K>� ����9܏�J')V#�nq�l�p�V�5�6B�^�y��@ήb����0f���޼��-5L�`�``.��.�e��m��=-v��vgoKv�3���!�e�����[n�����������z��,e�̢��h�zE2�Ӥ�-� oT�RxG
��|3oXa�D9�1]d>��&I���벳M�b��כh�M�t��`r��ܙ�t�'�m?�N���ˏ��gOR#��7,��9�o��k�R�v}��G���"n�Nd�4��T]�=x�0.���o}��8���=�؞���L����$��p�B�|C�r\�o<�+�C��h8��%G�̍�A�.<D?�dŮ����E�l��Otyn{(e|y�Bc�/��Ju@n;6���\���8�͸L�˫�I��8a%Wy��~��\��,�w׸��L_��B�S���E~
��#NL�(�jz|�RY�O)�?0t<�"F������Rbڒc�Q���V82����܃�ӗ~��V� T�_	�rX���G#o4:�-�@�^��˫�-4h����NM����!���PE���c�Y���y��� ���/ͦ/g;��V��p�ש�����0�d�`&�G�ޥL�a KL	��E��"�.M�A���K�JF��]���]s��^*8/�k����n�w��00�R�B$<@��ޔ}��{�g�qu9\�-,�iT�֛�o�ř*a�#�-���M	�B�%Lˎs\Q/��fS���J��H�S-�`�9����Z����X7�K�\��yzT�Ҟ'��kzs���wz�B,�H��YnG�2�sd���tt���Տ���?������{�r;Ugfd_�8H�{�B$n��0�y��h��jo�^�E���p��ܕ�_��QNEu�\���Mz�.�K�<�>����Wiz�)�e����]=�]���>L����'����E�[m��F��:��iY�������\�,2?'~��r3~g�3�W�@�j%��ر�}
�@v�#ӝ����9��a �	�5x��ؖ���3��@R�Z��rbh.��%��^$����,~6Nɣ���V�l��J���+0By�U����6�R6>3��S#��,�\�0ϓq�}w�:[
>[�B�qL�+��=\��!�"�7Q$J��Q&������N0���/ﵞ�T�]�p��t0�f��}8�R��k�=z��y�̊���c����i����co��WI�~����~���U:;�2�e	Xjҗ �3e[v��%E<���`�2��׬b0c!go�C�g���xb�� ��,G��� i��'���;���b)�[3�8�\d�H2dk�b��8Ź�"i��h��$-v��0d�0�<� �J��~��q���w�����F�KB�v^,�&�MG�h ��g�f��A�����Y���{ ɮ�J�������,�U�m��i4�!A��!!z�Jq��3�ډYm��0���b%�$�DRE��@��$L$l�F�jS]ޥ��g�=�e����ٕ���G4��*+��w���sVȒ��[��v+��O?	$�^�Q��I�UT�gYocM�mI_z�udݬfJ�K��e����lk��enDl�%.WKeu�z�CH@FD��ڽ��XhH��@�n)����q��'O"(AaivV���R�������?�_�2g�G�mQ�7v.*Ś�ұ�|��IE�,G��B�ؐ`�"IPY�WG�T�����s^(����s�t[Z����ں��9�|�}��:+��Ay�C�|��|H��[x����_�-���2t��,�%1��{�B(Q�����{t*�}�'�|RK��d��5��� �A�FX]%e����N��+���*��EA�� Vd.�IlzQxL���W�K�|��������)�#�!�N�hd4��v�\���-j�f��Z����E��xT�8<W+��G���o���z�`���i��>����*�������0�0�Z��	IL�K!	3�w{>�����5*�RK�ә�؍6���>��ϬT���7OI"�L+��W��	Շb����]��0��������ƒ�/|�Ȩ,䲾�BE}�@�r�����H0����EI�l[��W�i�kf[��m̀�ŉ����٧����!w\K��L ���֦m�����ϻc��a%�T�,�m�}=�c5�ԾZ��}���j+��=�+�:��H��G!_�Y#G{�I4�M����-����7^�� 'H�B���Wx�ܚ��z�#HO���]�(�ј�����^@(�����_��h��������@?x�$10�c�L�K���/�ه�1$�>�����ԕ�D	O
���UʳTs��m{�O�ܩ#*uK��Bf��
:����:��j�04����`m5�%I�\_�iޱwJ���/�R��<�<hXW���@�}i��{���C�	i��	�Qn�ם����.��ߝ�ϭ)�T�"�������r��o|��8����1�/�ȵ��2��� �Ν����hy\<p߽(W;�91�c?����7��)��7���UU̭����A#��YF�׉	LI�SQ^�Y��O�Tz���k�4D7Olq���F���[̽�#�{�ZI�R�Cr�9c����5���hBC�[޸D�ή$h�*�Ր<��E��٪��bC�	6��Mĸ�y=A��g�q��v�h��ψ�thi��+(^���&���'er����*+5V��	��wK��jA^ӄ'D=G+!��H�9ln�ͶYr���g/��+��V�k����D�G{���S�H�m+��P4��:mQ)lb�j401֢����5R����)�a_,%�Y��y�3"q���{�{�~��F(\q����*�7}O� ��v���P
_oOU�R�(���/��[� �ǖ�5�O�u�{�EY�kغmB���yA�e����5���1Awj�����Zv�N�������T]��,1�^�",�,ݎ�/f���Cw#�k݄r#ʢ)�ʴ�<�I����d�����9hH����bppuA�g��qyfF�U�DX�D4��$_��4x�LMM!";�0ҬFG�(y�ee��P��h8�0~�Oc�SiJ���ĭc������Xki��ו�����|_�ʟ`$�恼GX;���U+�$�x�����/c0��jO�P���".]���R�a�����Ѭpv��*��v�������T���^Xͩ(L�
����y��ܪP��m	#y�(�4K�O�����S�ߖ�!h8����y�{�k�k^-�$��0,	���AA�A4$���9��_�:!s����
��D�㏄b�4�Z%`D%�Tmux���נ�Vr8��AJG�9Y�I�f�JH�3[���׊��k�4���;=]�rUX!c0ߘJ�Ϥ�o���JQ��sI�IJ���'ɐ���yރ���6�?���ii��eO�Ѣ^���QOiJ��J;�w�hIp�t��
��M:��xYw{Zn'iG8c��g��E����U9�xo����5_�A�}JR?A`8�$��p�\E������u�����X�8�19H4�A�ĽfI�bKPk�,\Dף�1U�N�L��O}?����U����9�K?~���Lb�¼��G(=Z��a|l���s+�ֆ�ҺO���U�(��5������޵c%s���SttӍ�P�V��bvq%I2�s(Kx��{����C��K/>�d:�'?�1U������� �5�>u�B'�������;LlŴ$kKy��������Sc8���(b�Ip]�-)I�#v�{eQgBkê��ZyD�^��ɹ��rH2Þ�����ݭ��-��g��L;�W~嗱<c�O~��Gp����w����*���?@8B�R��piq�`U�;�����/�ryi]xuG��(�I��WV��}J ���Xr-$A�n���ɏ�3=���vV��{w����A�[�$Ǐ��m#�N{�����u�u��x�� �@J�#�9wnߎ��.��^D�Xĭ�ޥ�==�� lI2��sa,���<��.�&aE_�}'@��\���u��C&�&(���F��ɹ7iXϬ���*����^9&�ʽ`[D�;K�67kF��9h厉�#�V�Zas�n�̀���xZݒ�iu:��!3��ue��٪�d&��[�qU��f���R���*�ᘑ���)=�)B�G�N�g<�;�lO���vك�$�5|Ɗ�o�i
�=�E�¨��=F��P��!�n_K���Q�k\�hF��nI0�5�GĠǍ�+�]S�DY�z������ᆝX\���;���Ϝ<����w���(��R��Ab���Qi�d7ڊΛ�z�;����εܬg����	VD�JQcM| ��$p�(�{mmE��#Y*I� 	�)I���<��C�	X\���p
��s9���HģN���i-�S1N��CH �huT_�\Rr��l�X�(:"��6-��7ף�e���V0h��$A�����C<HO���*5�nU��������w��8�庖~+r��QI�,5��БO���}��G�喉qIV���#ǖ� ^�]��ʪ���r3!�Q��GG��F6do�������JS�#�'����E�o�b�2���W/���}�����?�+��f@P��n�'��;���	I��럸{w߀@����k�R wN�fD�)���È�>,���^�P�Vq����Q��`X�{�:Y��ɾ����k�e�?ƒ��$G�ȃ��L�L�(���r_���{��/���gK"O���+�B_0���06��f�����t<�/����x�a�3�6L�1Ŏ����l�>��sQJ��>}�-.�,-3`rL��U���b�ŗ!K���_{N0$.��Yj�v��`��V��ݱ9-3�^���u��9fQ�Ԣ��'�7����$����V�*����lS���F��6$��[o�믿��`S�)d1����VG^ۡ���C��!A�^Sd���� ��(����Zk�8l��/5t�k�cR��`6\��@d �G��F����Q?�X�+�o3a� լ�08<����s�?���%ש%?O�%���o��k���_�i�@4���?��^����v�!���HW��C�q	Dd�۪6F�6K�gttMG�,3�l���-9W7߰[��r���ˋx��y-��9�;���=øq�0\A����k��W���p��?�o>���g��3O##�f$CJ��rAr=J%dٲm�ߺ�v����e�����uka�S^oW�	]�$���>۔�;��:yM[�o��n�CJ�:|������	u�ql�`ʘ�mI!�����=���W�9DcIc�T
��"vlI˹؂��,*��\䞌��z�����%����hYP�췇���e����ZUyN"A��׬H���j�4���W5H�^w�����΂T��M��vj�<ʳ�����<,�:M��6�t�ҋ�|����j�z��u�m��l�V�"0[����$@����;��O܃xOT��&-++kZ��߂EA%T-�iE2"�����YZgP������\zK���"1S���)a~=��kz{妱��Yf,ʣC8�A����H� �5��0��,c��2�������Ҩ�Ou��EԨB=�i'�3#G�PP�ʜզ��S�O�;��ϡ�	UÂtV���Q��s�jqڿRQ��]/g�9�� Fv���>����A�3�=#С�V9 W���|gՀ��#kLW�2AOdu��NKV.�%b_�Zܜw�q�^;r/��"�ʿK�
���99����-�S)�C���ŀ�%`�8��*�q̪�ӄL]q�<����C����j���("�5&ے�)!Y�l	�Y�>�ݿ��^=���։4�M�s�^ (�[Y/����?T9ݵ\�K�j���vI,�x凨�3J��}-����'(C�Wg3�Õ?!��0�������:&�[�,hz�1���zXb�X[�"�� ?x�ڇ�]^�{<�B~]��&�����2k���F�Lk��i�I�$#m7J��$2�����&sk��p���q����(W[Jt�`��׺ެ�}�g@	lN�L��0E����+纫����q�\���hȣjq4�aՈ
�ZMCW]�|��N�(H��Hr�\�5�$�%�E�[��n �as�n�̀~m��שUj�n��e8จ���Q�)��U#�E�E�C"�M�JY��a2���í�a\�x	����e	����L�Q^]�@b�bU ��Ȭ,�T�!�+��Ҟ�Ļ�\��h�0h��`OS�4�N9���]�轿�K��4?:���[Q�:��$����E���� ���=���oK��^�g>��:~۷n����Gq�M7a˖-J �
���Bh�>���8x伔���]�9�s�M�qus�˭U�[��^o��`�!7[K�P�u�c� �'�fg��K#a�e�dl@�O���޴�|K�����J:����z�U�H���PpG�&�#N�wVS|��,I�t2�ӎj(oA�F���FB�qw�
�� ��'�E:�`'Iff.+1k(�F.��̥Y�4u+z�6~��~_��Sr^GU+��9��o��Ɠ�h�Z��ѩ��������}�%)d�d��|���wq��C�ο�ZdLE�^ʮ���lݨ����L{��	^�\`j�}9
�>7�S�Q�&�fH����r��e�}�xq�T��I��Z�/�y��×4�%9taqN�%�f�t��ca�0�3ӳ��`�!�DM&�|V$��a
e��P.�!9�����QALl�R@�z�f<$E�5����vǚ\wz��*Gω�����&���X�+Wi!#�n��C�^F)_�[~k��u�m��h���4�A�h{��ҩ
����K�8ײ(�
9�!U�fb���E�*�hcҔ�y�5V�E����Y�� W��ᤠ�k�(�/K�%�5�P��r��U�L�P��eDc�K�Xf���)T��NU�,�0���'���=o�Xe�wM�<� )H�ԩc�
'I��=u<:x��� ��+���?��΁/��`��Yc+�mCۢ ���e�S?v�ٵ\^����- ڒs(��i�^��^�*�h�F�g��S��|e[aUc�C>a$�_��b���N"=8��zv=�b({����_�������%Y���}�XD�RC�%w��b^��XÖ�qlG�3��-o�苪�]3_��G�<}	T\�.z�����w%xxAs�`y� �I�/�V�H�5��*q���i��&��ȑcZ��::�q������9�
����T0�p~yI)�sÞ�ro�%h���V�Z���E�ufA��ي~��2Zw�����>o# ��ݪJ�+���j�Ɔ�ԊzO^]XB[���ʢ��R��N�<|��:�޹B^��<.\�$�b!A��O�@1�����
B�-	���K��<Kr�X͔�����ܯFj����:��14��)�*�۽m+>��'17Y�}#c)ad��<�V�jV�C"�|��6A�Ѡ$�Q�r�K+�g����X__�������]Y��7���
�{s����j����f"P<~
s(Z�F�ʌ6�J@��DW�GvyUe4�D�ü���қ5AI��AY�p��Y�رӅ&���ĉSjɸ��&�����Ou-���P�8
�V�� 3jY[������"t`M���T&��/t=3ck�:U��Rsq�6JEί�����uN��[o���f�����V��,-,�X���W���c+	�:�!9��+3ϟ?����`Z?�E�������=o|���	&�q�)�؂�\���>��e������Z5�H~+&���r;�U�(Y�ŋ�����J��^8���.+k/�<��,�I�w�\���&5 ��!�hrdm$J���v͆��#"2��v�˚�S��$��q.��mh_]�����G>�Q���_(,��P}��|Cл����q��Wq��2ֳyA������$���jNaxp@�����#�"��$8��*����q���O~��{_��3ht=��b���OaA�m���-#�ڨV��A�<���j�D��Ӿz�<��
ʒ�PŐ�;#I��A$F1P�"�z]�%���y��� bqy�ɫI&�5�����f<3'��1�q�%B~I�Ñ�
�6�g�@U )&�R4J��L9h�hH �J��}Ԓ�T�%�����{�MWW2�K2$Y Rr�ǩ��� !��i������q�׭k������Я�M֎�q%ӯ��hU[Q�-+},dc@��,&Y�i�19>�����j��Y��ƒ!�	K,[r!����R����)4a{,#}j4�M`0��?�n��D��k�u��|M��˕8��GF��h�q�9�b�!��!l݅%��ܹSPb�?��,����r�L_����u8]c� p�����QȬ�~��U,,,h_{bb�Z[�~��٢���I[>���43ٹa���{6�Ȭ~L1����~1 ߇%p/�k�G*%�=��٫��3�H�e���ؘz���O����=<2��/葀��^|�yMBX�'��0���֚"�G�`P����� �y�l��@���Ƶ��@lP���t,�����F�ј�\�,8Y��೟�Y���~���o���%A�^�p�v��$�uR���}zqΞ�X<ג:�5'(:#�~l(��"7���#����cl��{״FB:9��28����F��zA�p�?)�,���SN�E�K�zr��;wN���$�CL#���ae�%��?'A8�}�.9�d�{)װm[�dg�9���:Ψ�q�!u�'S$�����!��Z̢�[����^��%pg���Ϥt0{���=�� ?�<*����5c��J��}?1��}�d��S�;����IQ(7Mn�Я�m3�����Õ��[�Pu���Mr��4g�f� �.	P�+I{G!5\
�=)�I�Z���s���S!�K�#XZ�!I�*TѴ1}����a3�.�'��}�=�g�ж|��,�z4�uV�Lk��G�4��M�W{�ԧn7���h���hss^�ő_�)��m��P'����gt�r�.�+�*��,���?�a�u���;�TF-�Ab,wZ;r�������DɡXB�� z.!��mJ��H����jc_�i1c_l�wڲ��X!����+2�%�P���=�p��I��%�7�����bN�_D��[���{GI��$U�5���˗�4G^��K�����s�-�I�~ӽ��G�H��e:��Me�����̍���A����P��䭜|�k'O�	\L�r���EC��&���bqA�a��{���1I`�@#!�}c\�#�P�9~�ё+	4�F�Ц�#w��i��u��a��$7�E��n�����i�v>��.IHC������'�
y���Uچ�8���{��8K�+�kx��`�I�v�T�I��cS�	�ϯI ��cG5����z��!�Z(׊�j�e�	o��v[+Q��UV{��T
y���=����2�$�˿3��}�KO?��Q��0Q`B�NI���!x%h(�$$���a�K/�
jM�%�	ʵX��B���{��L�Jq�Ѷ����W0����j5��[�a:Q�Y�\ԁ�u�l)�p��Q�#0$����bF��h<�x"�l>�dzPf�+˚ hS�m7���vjxTQ8����F}�2}MΉ{���pU���5#P�^<�z�}.�Q����b��gdc7�2X׮7Z��W$ ���+o*��S���Z��ɒ�06����$!�� ���k�L�-�DN���eܼ/|��:�π����+��f�Y=zT+%Ac?�3��-wn�>�`z5If���6�H��kՉ���*�QF�R��k��y��֖Vd��`��%�e���{߭�|\�ctQ�|�XE�PR�M����ة3�p�}w݉	tLH�0<�����~�3.j�t˶	<��Gd��딁m�������zFLf��pM�HҲ���sH�������[gT�WM|$X��^5���}�-�QY[�%	_�.I^����rE�rr�|r/��ד.xlˬ
Jf���#�[�;�a��b��$=aE�Ͷ\�P�ȷJR:@7�VG��A�-�Y���%�`ڏ����s�}M]�IR��������GLo�����㗧/iy�U)�����A�ޒD�U*��/��kBky���]�C�Wy	�%��t����Ǟ>r�	r.�p]�R�r�xTf��U�r~x�|�*嚶���IT�%dr9�5����w؇g�� I_D�5
�soi������0�wu�8���86��f��o��o� ����۱�n�׺�^Ѯ���VS�M	*EY Ck�6	��hX�s�nP���sJfz)��Ҳ_(���<�����G02<�3�,EҘ�n^�0X�-��v�?s��ePV���� z�D�c��c��HI����6&�H`��`u�(���@�Fs��3�>QD�m�l��:S��R��v׫���g1�u��?.\���`Z�k#��s�*�{�-���W3� �
Ϗ�Sǵ�F��E�>%*���Bt��HrK�㼦��Li��HGд���^D���Ջ�ա�nj0��ռ�A�'P��w|gR�8~��I�l�,�^�kx�;�p������� #��2D��&�eA�r��.^�J���v%eEIv����r>�kw�=�4d૤�Kې�4�w�J+5tv�I����c|߉L�r�S���լ!�&���G�rޛz�%����_8�F�����&Ḓ�V
:��}�"� �H&)�s�=x��e���'	gh ��w=���U��e
.��z�l(�#�H��fe�c�Ǿ��d]u�k�7+>�4�I����X����s�R'���Q9/r�`g�YMS�'� ZSv{��L�O٣w����0X֢��ݐ����VW��Sc�x2)/�#�*/e ���"*	��p�=X^^�zn�#���x���Q����S�O��$���G����zjզ��r�����]l��m����V��ԫ5��p�k�S;I��ia��t�DK�5͈��zY�h4*AS�iٰ�O�u�x�WJ�t��C"
2�gff	*ه�Es�J�ř�&!	��xH˽6��c'��{����H	��+U�ag鑥UU�����*|vP�I���3�>$�]PAk���>?�dqnڽ*��+�y�c��]\FWQ�OY�%X��)D�i|�;�GnM�߱��߇%	�K٪.܎��d�xꛇp��U��|PV�h�Z�����(���r6����@GJ �K�Z��\�s���o��ۇ��������V4Nv}0< �R����z}o �9|��C��lԴ��`��4�VñaY����Y���s�v��E�)$�ȵ�U��e��]-�z��v?z�]�u�7$�սp�n_��s�E̲E�-N!RH>VH�n�;~�V�[��kč7ވZ1+h�v�\��ȸޣ��"��=366f�Iܞ�>����w�e4_;�� ���l]	x�s�h�KБ Vܞ����!�B�]�̱UbHs#�j"�k-��p���yo�A`T�ߠ���y�k��~�~A�*^���sP'bWqW��g��ʘ�VuO�x�c�힞G�����������j?T�%�$�HH�euA�Ч�uӍ�1����:^�8�)d
E�ΰ1D�d��V���=�����1sn���:ښM�ߪQ��/��Q��'��E�+��wzD�;u�=F셈�aɔ�\Y��3��`e=K�cjl���Kϔ�Y���#XY]Ey�+�����>�I`�s�������{0�*�u��.�.�*×�1��ⴌ����?��7�ԟ>���<�����%ᨫ�:mH;�Z����	ApLTh�ѐ�~�\0un]�_ȯc@�/^U�yY k�L�E�F��b#L.T�D{�B��(���׵m%u���)���p�յQ�k�� �a=S�TƤ$1����y�\�ëG����	�t���hJ�uP�6���kz�)����b_���"$��u�$"쩆BQ���txm����.\aI�<����=�< ��pѧ꜑�5��/f`��'2jG�2���ӗض��zlcyK�p#���a�"�/�kY>)����D��b��./�#�D�;܂��[���S	W���F2��ZV(�[Yϡ�ɫs %�VxC�b��o䰮��}/���6��%o\�}{3�g�}�}	�L���'&��F�<(���!Q9mV%Qɗzo�4��ԕk�%�6�X��*,�F*�x�B�3���$-�'?���Űw�.���Lzy���&�4���]Jb��Ys$���S��#��[��ju�FZY��&��:�6�u��m��7�_k�\	]��t1A�>u�rd�e�	G�OL��\{��c���9�6�v��`R��_TP$I��ǎɭ���d�	*)��V� �nS��}�c�h

L8��PoFP����,�!��zU�H�J���M���O�����J��tf�Uy���zEK�!��%���Ү\��0sѬIrᑤ��Vn�ݖ(D���5E`T�b���"I�U�I}UWΗ1���Q,��n-t���f6�3�=ǧ-�^��`~�S[�}%�%~���ax(����g�Q/����9ܨ��s���:tyjd��Jh����/G��@��L *����f$��^��	��!�O:�P�qB�z� G���ƨ�����|���G��:�E�:��W����{DQsm�v�!�k��3Μ?��gQ�z���wߣ�W�S�˽�;�1�����q��eA���I �~�92(����VA�6�~�~	�r����H�� ��/�K�j�uCR^k*���aϨ��_3!�����g�g����I�j����1�T��5Z딣�dE6_����-PQ;��}WD��R�]!�S[؀�Z+�iٵg/�CimK��>3@��o�\��s�R��$��+˲�X��ΚD�8+R P@��.W��r�^��܌�Ѷy1�����z4�N�,q�g6�z���˱�,@>E�0��'�2�]�5��qĆ2��@qtg��,FFFd���415���yACf[�_������P�trj+Μ:�X��p$�s�n��X�'���gm������|�c� �0�\��SZ��bH��Q^�W���}"��Zvz%��8�?�����E�?Td� Ԧ��װ�-;�\�&��O�`X�@���0 �tԲ��C��t�\Ǚ�.蘐��~�0��6�#�j��j�Ϗ\��v]�%��ৃLmyM��Қ^G�-�B�q���N�oO�Q�:������$E9�u�w4ppQ�v����;>��~/��2�x����7u���'�}���+�P1�LiG���Ư��C�T(���w?�[\� qۺ��7>���&��/<���U{��{$2r�����H�9�UĴ���%���4P����g@��K��Ԡ�(G�Ǯ}�՗�\qQ,T�ꫯc�(�S��t�hGt(^��g��=j��4GRzK�8�}���8T���*�� �v��j	[/Zu���*�Ӑy;]3��s���-��OK�D�@����I�g-��"x��%=rL9*�C�A���u �=DU>�����+�?���ܮ]�Дg�JA�I��D�YA�b�[�6t���A��ҷ���zT��k�$��=C�,�J�T�����{��o�maaa�����r��[ZZ�I�]�����W*�����*�Nέ�:�Ҟ�<�E?K]��!�w�k��U�/IPs$����D)��`Tkr�d=YlY�#h��Q��h��2s3s�f���q(�,,��I��U�j�VI��-��?�I ��Q����ϣ*����bt`gϞǥK�J���Y|�c��7����H�@�
t�]	�kj�?Q4�!��u�]fۥiLא��h�)��Q��V�Wz�K����9	���ce�O��r^�?;�S������%�����O'Pn��ڬI��V/yJ��=C
�*�y�z���~r�#V�O�S��Q� 6m�3�����*�{�my�R��^)�x�Tv4���2��Gc��Ί5�-�ft�|V�&����\�jf�9M����f[���e]S��e�Y�q`�qxz�My�����a�ה�͠9>�E�����Ѱ\��\?W�KR�����$e��~������{��':�"L��8�����V?X�� �LG˺0f�5�^ero�$i������V����*E,�����Ǿ�1�k�)�fBd4\�Eq|�5�w>h"?���A��{�ނ|����]�����mi��(��+�.�'�,��:n��<,	rS�����7�Y)=VNa���ow<�çp�/���D4�P���|	A��ca5�颠�*��>�mn�˶���[����Dn��A�@ �"�Juayy��S���,-�6+�=�;�v����=�$�Cdb����"cK���l�wV�MY�tG��\��!�T.se_Z]ҀmKp�J H8I���ںc��NW5s1���=�܎}wܦ" �F���P�nM��{�h�Ei9'�@|�G��SO�����8v�$>�O*3�����;�Wm��ELA$�PCt�:s� �^+�i�m�ODMLN8��AxkXu�~�n��,��l�[��X�}>7}e�z%�tjSN$����iT1�m��f��9A�A���3Ԫ��e�b��Z��ϹaA޷�n�Y	��lӧ�L�dn��l����
�:��Ʒ�abrR�ЗVWu��s��jG{�.y	�����?�a�}ϝ �rb���w�?�>�|�$A�V�}D���������I��2�	�F��6���7�`�1t���u\�uW�A׫�oj�Ǳ(���$=vT��2�e4klL�����O;�;��0$��2��\�ٹ%t$(�j%�u���5��=	���\�F˝v�����Y��^�^�+��;5U��^[Q5�0[#Z-�}�?�~;�-O'?Vc�b��m�Xu��������X����#X]ˡTn����k9��P>3�s#Ǣ+ϖR
��N�ɑ�d�����}��-�83�uݮOE��B�3D^,XZZ�s���&�}O]�h�ڶ�r�7��߮6Ů�f@[o�ɧ�À�����l��F	��["�� �t|P�y��P�����]׊��#>�U������;o���c{��d�f��$[�'���HX��&����ᄢrmʺF�TO�4O$�wZ�����F#c#���5M���|�%��bD4붵�� �cC�^jd�2�䊈�{�b����_���8?}N��\��p�lK@�d"��|��j)��r�����.OO����{XYZBH�î=���TEg��,/J�����*��D�|����w߮�e���ڟ?��^|Y�M�VYM%Z�$K�w����睸]� [�`z?p�k+:WM��$�>�q.�K������{�M��ɏ~ _n�W����O�����.<������m;~����2N�9�J�t`l�6q��x��]��Vn�xʖ05~&�����A����}��x�[@^�3����̼\,���b�|����jPd�C;V~]uL?�ڨΫ0M�N��O@�1�pif���Sgg�l`��=H�!(�+5�FS�3u��SչJ��bf��QԨ�p��D4�
�/(�K�p��4z$y�� �f�"	YM��q���(^��L�8�Ʃ:�I�D���t�s�}��twT�Xq�$�T��V�ZA�����$R����Rk����6<�ɩ�Iɽ[֤�M�8'�$O�-���5�L���&	���"�n	�b�Sd'"I2��=S��$��3�n���<&���A��)dH��OK����������z��0�����%sn^o�62:U��m4k[W��B�@F�?�~��h=�0�I�E��G��A�����"h�=��'b4ƽ��C1~��U�T�׭~��,������ �~z8w�Z2t�P]�eU�iʒ���R��{�Zٳ����ff/"SXƣ�<����'��/�RQ"�8~�ӟ'�t��N�ݳà���(�Fq��VLm��~�_��w��I�qL� ���-��u��/���ɷN�=��{�J</����)����XX�ǩ3՜�D�mT�x��y��x�чP�汴8���<|ﭨ���W�J b@��Ak�E�����'D����p��n��?��c���E�Q%Ku��% {wn�'?�,�c=�(�g�{n����o��� SU���RB$Β>G�$ْ�|��/!$�z��v��m�&�3��0�g�%����$bq�i�̊!�q��d<׌d)WAY�P��.a:�j�¾�	����w���gi,W L{�NW=�=�x5�����}$#��Q�d����|�#����\(��5�\����M��|�`������f���7�G�G�@����J��j�Ib��%?����un;D�	���5/W�rOw�>�� +D����?f ���U� &`u��ݴ��^��͍f[Z�
�9/�]�T@(���u _ɻs��&���	�νTlTu�R�!��|��<p��%���@ܮ���;^���}�e�m�+YT�+����g<$�°���x�8�GK����J��6��`�,���7�A�H8��; ���1�H6�S�C��4�5��sM��� ���g�E��Fj��ݾpF�kF{�:�
Е,�A�[�g���sU�R[P�؁���$DY��H�����_?��`DE4�,�F�eA)ʢ>"hwL˞��3��KZ z,=ǣ�I,�{�-�G�YE��Ù+�Jcrl�� ���]8u������pu��󧏣��@�H��;���Sx�>��_Y�#��DIŨą�iG�{�9�ٹ�uM`H��-+�`n?xƆ���G��;�s\�~�>?~J�\YR�-�¦���{w�S��+*��E7��a�	&�zXAd�9���PƮ�1����K�C�Z��ʌά��>�tBQ����R�'�kYC<P��9A����r���� ~�W��'{o�/~/f���Z�IxC~M�8��D�Zn�Ў���
�l̪���n��ykp�6�rF5�x�Ss�$=����$��#.3&+��+A��1�s;�r=wKW�%���/�4W)�{�	�.N?p�mC���3��|�@R�Jר��� ؐݻ��'r�����Yo�5����m&�����Z0����b�*'����Q0[ޯUma �֑�J�"�@]�ۣ���w�b����cR��eW9n�� 8F&���c���1�X,�#��zY�|i޳�8���q�#�o-�k2����c�V�����%��x��*j+c�V�R�Ȯ��yH�r���,6��f���R����'o:��e	$�Eͻ1:�:���PH������m{���*Yk�m�?#�����عF�a�Pٿ�Y�}�՗_5���a��@{��{5��Mp�����&�a���媐����\4�X5#R�Q��cQ��@s�NW�+NI��$���	����_�R���?��BE����pan/��J@��o��Sp+yA=��t �T �;v`ϭ���ݮ��¥/���ұۦ&� Qk�S���
�%�oEZ���\�Zc�ߺ�4.���*��J��&{[�	���.��MGc���1:4�ٕ��Ju�$��?���G
���J&0�cJ=����(!���0&%�9�+!�a0�Dv~IIpZ!�D�P��W�������~��nڒ�����=�%�����<�İ��-�����~����s��ͧ>xOg�y�\��eL{�D����y/I���d�)��kG�?w^} �CɴX9�LNu�9��I�9��+��-I����N\	��bQ^c}�k��J��BB����$T�>�%�]udM�͋8�e;m��<s��E>G�������ȵIi��,��RŊ�+����qLlݩB2���K먬W8_�N<���/=/lj���V�!Ik^�/)�y��E8aه�$�VB�$����`{��T��ڲ�����R��*Ļj����4kU8&0�X��Lŋ�ܮ��o�7���k���Bu�q�!��r�\P���۰M�r����J�w�!ǻ����]�|��I�"E�t����qAWD���.���a#��Tl�B�SE7��:f"��#S·%PUU�����N��|�)�/�Q�Ŗ(>ۨ�)�Bl(�\���RC�S򚊑�Ϥ�v&�d>��n��8��Wt�Ր�M�;b��F\���g�V�bhdTz5As���kH�����s7�pP\���Su-V!([�s� ��tJ�&VF���%�h5::GR�q�N��n�@�2.��������E	�5A�����NYQ�綏h��D"���o�R�<��q����)/J�d�O��+Q�T% f�����c��WIT�������:�$�1�`�I ��7F�5��U��mc�-�v�j�A�%l3��S1�C7~�x,UI��4��k��	�M?�%}	��pA9'�l^��mf�)����5O�5a�ο;�Ԇ���(�3�ȵ�pJ���F�A���`�����p$�z D��PD�U$�m$4D��>ɍ�,�7ku=/�|��O*2�W��<��-I�{�*�sK����" I՛���R��=gԖ��1ꂼ��~��	�����}�<���˒���/ȵҪ��l}��][�g�L�Z.���1��j��]햗t���ZΖ*[��M���h�,���������۾�q�1����ވ�9>ľ�
rQ��2�[�ۺ�	��R��� O���m颡��fK8�p��/��ԉK�ǵDh�s�$����_�箵�^M����~���f���c_��+í��?ݖ �r#�j���eԀ+l;hV��X�2�q�Oy��=��G�xX���$?)�J��"�� �{�{0�Տ��ą+��q\���}�������#���tͳZ�Q�fD,�j�Rb�"�t*f�&���G	xN��j�%񐼾�b.���I�4Jզ�Ϩ�Mo�t"��OT����y\|�j�I�F��h~xpHP�O~�#x��Y|��[=k�y��̪���0�������l۹CAx�K8zn�� �Ү�,�>O�#=9�I�����H�4�MĈZ��[���F��ڸ�r�\���LG�Y���TM���z|Zĺ}w=�fm	Ҕ��	l~���Z�Z}�]wC4�ɀe$r��'�VL��c��| �>Wk>�'6ĸ�������$��Y�TK*�R*� ����{���L��u h冤��$L�[-�E��EU@�jq�D�y����|��ךr~,'�Y^�Q� �n;C����3��'YL4�����xZ�"Μ>+�脪�B�J'5�7�Ip]���b~nZ�rUr̳�kH���lC�Ņ���!�7��Z}SX�z�6/��x�
�SSc��E���"h��l�QG���k3��T/�D9Rs�´2����lݺU_�E�3��6�kY��W�1��#�'..�]G�Պuc��n��QFW�}ג��*�_�r$Q�Ǌ�w�~��J�t�{Xʕ��k������{Ď���86�mb�Ν��59v\�."" �]�ݏ�z��>UƟ?�m\�_F���瑙�F��"�0��g�թ�&H�#V�_N��X��0:l����.�$�'03����s��M	�,v�\��8����x�AH�"�����$X���+䔩�@��A<��e�j'�Q�m�sQw�s�w�}��ތ�k_ �y���V�w�N4��ȖqB��P��~��9|�ŗ1<9)�K-�A˓_��(�B06(��E����V8��3�ݍ�M� kV�ɬ�ֹ���+�M$�8^��'�Ya& d!߀nd
��,�7�2�D���e���+#b_���-� ����r��?�h�$'<ou���-In��ro[�:��;�����R+s%I���?����-�g���@G�����gJ����X��?���jm��	ЕcuTw��|�z=��ܧ�cWHv�@Z�:cLbd�˂����>��k�!*��tU����b���
j.p��,��8S)�9�gYF��㪎�[!����jҜNiE�������SE�^�ۤA��v�l��m���t|^˱���K��5қ�)"�\�swm��ĵmnnN��Mn�_PУt���[})o��i��c_#��<��{�r�~F�q�
�tt�㢴1´1����F`/�*��iJ�4�)W0�l�����3pz^��.B�`Z�cΔ�O2Cb� � (�-�G_�:��<�8�r��>p;�s�]ؑ�������gq��q��I ��ؖ���I��n*8�귱���k�Ȼ�Ԇ�hL�hO��ְmrX�6Z�����<��eL����t088�V�>����]5�;���x�$�u��9�~2�H�115���<�yD^iT+����)$�&�Eд\�I|�(4eQg%!��Z��ӗ1�}���Q�k50�2�����@�j�3������(˩.:c���6���/�ۊ��}%5[�E�UU$i��N�]�B����3}w�Ǎ������2*�Q�>(��T)6$�YG_*H��H0$���5.q=�1�s-�s��c8 $�����`F�?t:���%��Ǳ��=*�r��i|���G^�yG�ތ]/�O=�	��'۝�������&�U�[3���D�.XA��4|�&׹��dLL@9�鉆��1�"�k�L�9�g��9�����,�$J�X!iir�չ�F��h<f<�e_X�`YXU�]*���U����]��gK"�+���Yx����G�~��u��J-����6��x�DH�
p싦"���jQ��)��W$�B˒ u�QWa	n\���Ӳ��d�/{��s�U�؆�8%%Y���q��m�g� ȶ��Z�N?��HO,�Es�H��$G��Ꝿ��g9�$� ֚���%�O�a�}��)���5AP���$�t��勂<۸��~D����2�ږ��{�=w��w<�-i?f�
B~��8z\;�:���e�V�S���<�1e���K�j�&Ms��Q-Y�bnf���سo��_=�]��R��NUݩ�Q	~,-�bj��Ӧ�W��W�˽�L�B5����gJ�ܙ�U,.O�c|���$���;/H{䆽(6e�5o����i9��\	�?v�
����c�;�߉�n���ݏ#3�J��1�}
�){n�{����S�T=�[o�@$��8`}yO����v�!9֛�����ꓱ���N���E�/2X��i(�^Lx|HȽ���D��ohxw�/锞Ǘ���%����L�%9�?<�WiZ�n���9y᷍��� 5g��}��ك[��5	V������t�=�v�ܮ��������W��'Ȯg�R���O<�m۶�3�@��[gQ(���?���O��[oA���=Y��K�qvz뗗�I"1�7��������� V3�DH����&S�FKm~��1b��Gv=���Q�kА�L{m���7PՊ���J(�R�N}�Z�#��%	Lbx�$�7�� 1��x�T,9�ܮ�m3���7�e�ΆI���*�݌���Bfm��Π�����H�>�fɍ��?�ʟh���+�7�SB4==�����ع���ײ=7U>S�L(���}�-�Ē�%���ʔ�%�Ib�!���s�<�39$�)Y��j�є�������x����`"w:��ظЅ�A4���q�<���!������Fjx �臰,��nAU��qD�d�����i�V�GI���sp�����R1ܦ:�1���/m_�sX���sA�����ʢ��3'��*n�w��������"�R��>��	`�s�;v픟ђ$ �����;��G�"�8_T)�h8(#�V���|�zձ���*�U�re�g�x�����Y`�fc���̛�PT��4G"�(MbN�w?v'�5��1a�Ά��ɓ'� ���>�S�����ݸW+�,�~��~38�~(�KFzT���Ը�B�)IV��W?��J�SҞ�aq�(�����ERG�@�z��%�I�he@�ujX��+���B�JV�񍧾%IA'��e�GI&h���AGg���vN�D���O��2��x��'$��E�=wF����q�G}�}����Ʋ<����z�8?}A[����IJ|�C⩧�V'<NILm�*�֏�W����-0%��-w݇_������M!5�M���Ĝ�	�t4�z��r���$0�k�Ʌ\���|&��i2����f%I�?|O���Lj���We%��>Lʪ�:J��%	��b�$�Kuܜ�{��u���1R�n�ڱ��u�m���&��E�3*�������е,�1��3=ꁁ-/	"�(�sA&"ZZZ«����`��i�0��@�`����gd���	8�?�����Tp����q���*ٺ\����6�;%���uHǢ���S�*��l^���Y�ɶ�c�Q-A�5	�y	�y	d˂J���O>���O~�j/�=ܶ}'�Qc�M�R����	�b4@9☖f��V%I� h	�畁�d:��k�,_P�V�BS����?��K�5���u-��*�%MR�nh�I��q%!	�ȑ#x�=��%I��lj�V�1:��Ө�*~a�`�H(h5_��1�Dgvy�|^#���`���+oԪx�/^�_}˥*�� 4N\��џ�_�et+�� �6¿���0R���w/����qC	إʂf;�2�.&�F��#G�:�@'.�C���^A�CQ���-����#��'����L�(��@�>���7� ?� ��"����;�u�j���έ�j Ԕ�D���>�(���%p�A���$��9�}�K��c���*����S!��dhH�ÉG$�L��7�Ƒ����صk���H���}X�->/��y}/^���ޮ�U����<��{O�l��P���\7��Y���m�Ƚ}zqE�U)��d�$�ȭ5��c�H"���nK�2����+��7܌j1�[#=V
UI>Qq���O���+����6����嘻�N$��$�5���a���\���{�%����:+mN+]G�f@o6e�fO��m0�7����H� ���@����"&h��<)������<*��tE�UOg��kA�=Nq-�[� ����M���7Lc
Zp��@�>��{��Ĺ��E��TjZ��G3	>�k��Y@�Bu�m�r� ��æ�6eNI �9,���Gq��i�~���������XbH��py#�/�"� (�ڪ����,�ܖ����"�)�1���s/"v���P���=r���:d����P�kRC\$�`|l3�W�/�!]���<D���a?�u%_���aDCTs�J@_��GO�NI��b'a�cYAi>���,ڧO��TDQ�ڶ�.�s��#jϚ��V` �����%Tڒ�@3�RU������:�|��RE��C1��&�JD�M�t�;*��s� sA�~O�VY���R���7���mIO�DB��*�+�u_ɮ*M5�-ޏ^��t(A���pɀ\�G�:(W
چ!\���	p�����$A$�>�t%�`a9#���s�=j�;��P�D( _{XG�3ZYY��{�Q_tP�đ��k�/{�$I~^��,_�U�g�{�Yo�~� va	�@�%�"(�$C<�u���)y�A�4 �  ��.��;�cw�k���4���Y]3��a0�����2���>��^yǎ����Y3Z&�.���_$�Dޟ%u��^G��Y]:{���NM_{h|�ܻ+h��jo��8
Ē�:>1!��8��}��N�{�abrNf�_��x�����;'q��"Ƕcmz]U��*.�}���9����������jrz�z	XW�r}��$-�d�M_����Y��i��9���h,�ygg���=�$`��9�Y�LzS��:�6��(�s��;��{�h�GP7�́�ϸ�p|M��4�P��)�+A��0	3f9~���+pOl�D2׾��S�V�U4�43����W�e��e��b@�j��]:|�?������9d�j%��4csn+@��R�2G��}�D.���P��V�nUI����P�,5�3Ʊ���>��*��e�{��W��_�,���.,���� ߎ�=�22�,S;&��Dź*˶���k}`���0�3��)����}`?��٥�j��$˲`SDMB�v�M�x�*p)O����wܢ~�d��$&�Ӻ�=�F�"A���2S['Ъ����4$�=�T�-����9���ϲ<�ש˭"'��o9��dƌ�5{m_�����K�˽b�$��f~��YL���Z��%�b�5>0 �� '�d�V�3�z��s��G�Wq����,�c�,�J�3U��X����U�ؿm������4�.kE���P6C>�� *�;>�#�o?�$`��B�1�m���_=9�Z�.+�.<����[�؟ǎ�x]��3g/*�|�(n��$�E����XԴ��M��U��w���W�ڵc��P"�FgK%)�`.��\۴wB��-p�߹�����@zj�v��Kx��_���H�2��![���} t��4�to���6ǎ�y&G�VU����~�R�Ϯ\����:-��d@G��6����
��4Z��8t~A���q�|�=��k�7��]7�&�_��%�c$@�=B�gg	T�Z�3F���������c@Y���a&`�~��Zp2cW7%�5t��s�4�ЬJ��|�Le�ֹZuز�ZV6s��VbOS�Z��ӧ�`||��x��Õ� �q{��`��EԊ\�=8I��e�r��ך0*���Y�kk�2#�2˙Y����c�����2����d�}��PiU��_XE_"�m�Gz��ЩI����^|'N]���6�dvȐ�99����8p�TkkJB�{�.�:{ߒ��}[Tz�)�AW�ŅYɢ-��=x�c�*�B�^����g����/#���E8�����(�"�q�M��G��& �T��������ѧ�uy���#�W�]eF38K�~��$�L�1�h9+�2��e7I�tRʮf���s�c�T�/�s&%%/j7���Ti5�D�^���\N��cj�Y' �>��W�&�yB2¸�����o�u�|F�ź�7m,���1�?���sl]ﵱ�1	
=<��+x����Tձ��RY^+��(�����$���7��o��pq����{	�$��q�-�̫x�ݏKP�Ēd�[h����9}Z��3���۷W�{'~�A%�-�w�8|�(.���H�k���c����%�}�� �Q���������}(�m�c�vu%�)Aɮ����s/���>���'���Z�&ǐ�.�Ԝ��d�� �X*�=pynI[W1��&� ��R�?���]%�Z����%�`IG��P���Y�j#3�U�
	��پl��u�m�5�=���`Љ�c�*FE��0#j����63(������R273reX��T�M2v�K�I��!MLR}�]-��@�i쁛�5��QV9Qᘤ�3��}}�9����-۵���[�2�A�J`P������_�����%�E5ɌG2!V"Ry�J��4�R�I�O���%]����%�!��S9�,�k�uɈb�Cߔ@����Ln��p��yS��l䘧���u�
U���XY��L,���~�H֕�̖ �edC�>ז$C��Q3���
��d��S}n����r�Ll��];��Ga f���t�4l���ڇ�����.k�X����octd�XK41+��>z�ӗ����=Ve��JV���؜�v�+�ecK�ER�q�k����Y8|I@�(��������%��?�_2��@��i���%�*�Br�J�r$2�<.
��% �X��<��)��Q֓3�����C���t#'A����ʝ %��t\��� ��xl���Qݕ�\�Ea ~�l�6.^�f[���0��n���[p��[��ur�J�Mg�9�]���m���� g���yT@��R���|����B������!�ukrO��}���q���WV�=y�&�G��S�9gC[Ƒ�ˣtyQ-~��u�yc:���R�*AX*f>ì��d��s��H�:'�% yz-��[%y?��Λ��GQ��q�k��.Fu;�R�f�z�6��F��؈�G5���C�M�h�L�������f��J>����f�NL`b��d�73��xB���e��*��]�f#�2�#��B�	�� 0�~_��:ZM�'�y͌/�ˇ���O�E'ϟGV@R
g.]��c��� -��欽����Ivӗ�7}�z�,�ZR����g$��{�j��TN�?!��Ls
��\(���TĞ�;e���G
W^���y)K tI���%�o�Q��Wp`�^=����Ӳ���sh�jX[]�6�&��땶ʹ�똜܆���w?�GJ�S>��ٺ�g&桲��,K�露�y�V+�1�]�y�rrq��r��d��*�bxf��ZF�ݬRx�9ӫ^ �-�zL@�E��V��� gq���At���bfY��z��:j��f�1'���	#�LKf�a�TՊ K�K�p�%���\�J�,�b7n>��k�*\�u��X����_�
�عs^;~
�ϝC*ׇ%	���n����.(�c��Tc�iy�+�n<��DZǳ8�>�s�Ʒ���w�F8-���T��.g��yy���������
� P1�W^��{���8#�'��c������� 񅅙�y�/�b�.A�\�E���x��Q�J�u�-��ޏ~뒕�{��r<S���b|p �x�����wݡ����K��!��T(��anf�%�x��7�P��=���4��q���t�D,�}��u�3K��g=�D`	�Ǿ[js���6��$�:^=!�E�f�� �q�R�5@�uqf���3fJ��?|B����,�3�aIr߾��j��|%�qa���	�f�m��"�=����F�,O����ńٖۦ���k�_�j��K�-�a���f��WC;2�-ه7�~'Ο���G��̱��~Yrl|g���5Lg��Ϧh8%7բ�Ҡ�d2u������
4Oq먮�	�7Q\YD�>`L�ͣ�@��������Z��AI_s�YVJ��e��,�x���eS���Icf�ǎ�O~��nK&˜4���¢ Ƃj �x�`�68���1���ɴ\������3�
�^8�o�zD�+��h��ǵ�O� ��xT��k����3>Iw�>%J�+)��t>�֟&�$v2m���y9�9l�Զ�X���=�d"+��F<g���x���k��o)�L�A'Sr G�-�5�U���1�řl{�[F�(���J����6�U���sV�stbD�����gQ�c*�DB%3sOoAs�Ʃ�֦�Qu�QJ��0�/K��Ѓ����cx���8;���q�����}D�8��>04�{�} �>��~�)�H��{$K7f��맟�@��w���/�ؑ��:t�m�c��X�&~�/����v�[9��]��s�����{M�i�8;c�p�3cI�#q>������ןP^�����du�BI��
�o��_�7�~Y�}h�ߊ�!ѕk��)�]���`����n)�xUln�Ͷ	���&��OC��n\���{���8�$�W���
�(A�2JS\������~)QN]�L��I}����o�g��1s�\E��R��-{�Ͼ9���H$���#��>}�r���Җ@�,v���ٜ�$��|�A���m_2�f�����f��?��F)dxVSK�����(D{�(����j]Vz����e����҉ �=�cY���=~O=��*��������`$����5&wm�̵�5.>��?��ʚ���=0�ɄY�N�=�/~�]��j��/}�+:2&�d&�<�x��L���s����?��df[u|���_~��+�gpa�d
򞒁R��2z�*��[�U(�AWw��Z��\<.;P�N[�6)9�t��Wem��`|x ��9��cnSK�4�I%c���>|�+_d������#׺�BA�M��'��v�	���n�b���d��+L�M$�6IΟ�T�?.��K9��*���[QE|���Cr�ݦ�)3�P��`R ߖs琣Ѭ���l�.猪K(��J@�Ů]��g�c}`l+n�`^]�󚜛U�������wI6~Q�R�S�pǝ7Kf.�K�9�\4^y���p���̙s��{�0��>:�"��y��t5�t� ���=w~E?�j�b�jU�Z,'%ש�dЇ�O�mX��G�r��J)�`�R��\?�~��3a�k�|�(�QQQ�l&��?� �x�-|����i�?��%kF��Ԏ����T��u�m�5���e���Y��Q5�b����L�۸d~(N�1��/�8�L�3�VT���7��޹��{�݌����S�4��4��}�A�=��O�p��iϝ֘�2�.##i�l]�b1�B\K�F��7^�v���Ɵ����=�;�nKB|�.�(�"��� �'O�3��Ç�b���#�+��C�eby�x̌]ql)��+�`Z�����O��S\%CY@i	)�:���i��9}�?Q}v%!�kR��0')}�Y�H$�n=��W�V�'�P�����Oq� ����2�>���R e�B�ހ�ܗX��{H�,%0��0U}��Gjke-����*��xC��q�.��@@�,�i�Hl?'A�Q1�m8��l�\�Q/��kê��!+*�'($s��x�����*��b�hYd�Q+'�VYA���s�GN̫,*�2ۼ5���@Xpu�X����hz-L�/���yT�k��7�}��Cx����˰�^�Q�u�W_V帛�k�=70�Sg�p��,�R0��`o����yL�p�ʺ&�#8tb/:��~KP��^F�n���1�55�����J����X,���g�j�Q�"mr���oK0��zM�|��u�-Z�پ5�����;��à�t.��?<��?�'���ࡇnT���_B�o�h%��-C�19v��K\e���� o�_@�7��Y�f�¨a�[W�=�/7�����tf��OLX]#�u��2\d2ٛ�uߌ��~w�͈���/���N
zks��1��R���;q۝w�̐:�3���*	p��9��s��q,,��~h��C)KU�7wR΃��*g�_����o��ݽ U@���|5�6��d���'��*
2�lBK�4?!��H�秴.�@9O?�o|ۍ�0==- G3a��-'���~�p<���sO5��"��d8���he$���FA����,�ㅬ����YM<����do��2r�YXS�d�136��l�G���	Wtf��C�[�UE27��[Q>�ƅ3��z!����ё7�1V���Ҽ2�٢`�[ S��֞m6S�ahQ��SnmX3Y	�$h�喛�n8y��+2<>?r�=@':{��V,���1��>��_�Yr2�D�|h�sI��7��N?1J���5I	��J��[G��r�&�X� �W�V����^�`-�?��|��jO��]��z�Ԅ#�+E	�y|��W���tJD��Ӭ�$���5,I OK��"�V���]�-��T唁b&�4�i�%�}|���ӿ�G(�q8I�=p+&���Lm�k�s�VLm�}��S[���K�k���L���
x�U��藀�%�ˀ_�tbs�:۾�����s��׻݊�f��G|חZ�2cd������E��@e���G�@�l�>�h��8�E���L�8���-�a�`$Y�V��.=�S��g%�چ��q���\^�Z���oq�<��fp�&�ޟ �+�K�鐖D��I͢�@dJ�0����Jl��}��H�ͱ7��%�:�N=�8U�X��B���+p^��J�i3�c�
y�[T�c	
�:��������H�z�ӷ������J��<&/熮f�r� +���
AB����V�R|1��C�KFD�B	4G7�D2-n���6���ZU02Џ��2N��kU���n~r�ZMW�O�5o3��8wa͋���6�W�Fk]�;m�x�jd�;u;�;�7�}Z�D9�
�D_�'������%qL����A�X�iJ c���᪷�ϔc�Ք�T+�.7��h����e|�ɧ�л�L6���'��+o"K a9�|^���U�̭jpƀ�"7����^���g.,h�
^k�.�g�FD\Vu���J�������������LE,�~���b�#�?8�����0�}G����x�����j0p<�gq�g�K����p}r�Ƚ�p�Ȥ8럡;���MR�u�]�%�\0ׅ��^���#�6[��f��x�5'xd��4lTF�Äe�����o�=�=�}	�ո��N�����{��Y\�⎖X9ڕ/d̸����f_-���3�C�,��e6 їFQ�#�sԍʉ�"*�#KZf�,��"ȅܲ�+�����ԙ��#>P'�ڱ��ة��^L_��} m1���f����������Y���㒡r�'�O�r�T�3�����q�R�nt��/��P�@�$�{[-�E�KY�d&3��޾��,�Ն�Չ�\�Vi]R8K�x(�b���A�L���`n�0B$��Lq��g>��D7l@>3��d�l]�ps�B�IKVI<ޙ�y��<��jn<���FU����"ᖧ"By����o?�F�%�i�hT���tcߟNu�1��8����~緱R�訥���Ȫ�9�� ��f,���a���hW�2uL ���_D��;(��x��imK4�LB2�&�e�OBg�$S����N�U�q��WD}ۑ�9���@��廎e��EF�īCϷ�#����ՌK�_���n*��6�箽���_�W��g=���A�3�$�?��Q,���?�<�����ї�##��F�D�4���w��I���Ko���_�ܾC����7K���v���&���{7����|�̚A��ۘ]D� ;�N�t�#����4��0e���z�h_��&i�T�+ԛ��M��1�E' A�
%2����1��0�w���_��H�.����:k�l�v�����Ĩ�
������M�8�&�|���w;:�C�M����ǌ��o��Ʊ�9<,��Ws<Z^�XeNUVר����;;:��|��V�]G���9�N��LM��;�3�m�C�^��`���Q��4S
�>�7��5�82�0L�qR��������*�o��$��	��~��;G�~����{�q�e����pr�"��r��y���ك�J�U,���/c��i�B9Ҏ�R2�i��fpW<����,ʕ"vc~i�$���k/��o�dms�zaf�����>,�7�[�D=_�E[
|�+枰�����/�9
�4�ldr�$sx�j-�:G&�O^ ]�<6X��աD.�wr_����iK��M�E�r�>P���{��Ghˈ�e,`��~;�^VX)by?R{Tv�]��GK�V�	��\����		l^�5%���O�S�Z���$�!���=�&G1�sT�.:�Mbvq	��t\��r�e��h��kt[^^�'��.�G}�.1�{ ��2`��`����;�٣��4���Gअ_�l���{7��`�j�0���{k*�{.��E�Re�rQ2y��ie귰kk?���q��
��ཏ?�;�G�<VK�L�Plx��S���c�H�S5�;*m�c���ʃ�4��M��0��MФ�3d��n�̀�L����r}�Ф�#0�)�B O��t��<3�XL	a*uJYN9�^x�h"��g_^�C+�lo.�,s+
����&�P�/H�c�m�Kw5 �r3�2/�x�N]�6�r��L~�5�M0t�,!�"��B^���BVԫ��}-d<��nʮq�1+���׿S����<f��d�v�D3�Ƿ_9��bY3L�uS�L��VV\L��Ƿ�7V�bn^��,}f�r�&�����ˏ��J 8��zQΡ���Km�L4p�]I�iGoܚ���Z��b��G'��N�ZE6ߧ��R����#O��v������U�hi�Fv���$�A��w�<O)��v�2:�=��7<�ZMr���� 6΀6�5��ZZ�`	>MֻC�?|2�'����*�v�佩mo�"��+�{�
@_A������K3#w��t[���M@�F7f�^���>���2���г4���(7B&@���v�{�*���pT�ޓ�%[޶c��lD��਌m�ѹ/ͦdC~^�7�@e�N�-<p����������m��î�{�J�R0_��p��[xK�M�ڧW4{�dx�PjA#0fT�%�����&���xU�=�יi.��G�K# �M)?c���� �$�q��B���R��[S��z���Y�NV��A �7-O	b|,��Y>V�z�cX�|�H��ZP!.��ҠL�B��x�)��6c[�I�Py<�Ǫ�ɎHq!jH��s�� (�1E7��I��x��ߏ�#��*�����J����v ���N��Q��{1��&���+X;uZ�+��q��q*�����g��h�{&�*3��ߤ����n���Ճ�������/����atx<��eUԈ�J�o��#B@'7�`�s�r�����0�z!9����Ui���7�'��f$��e�Nn��jж\յg��f)<�<���ܱ �v)�zb��dM��e����_~F�H�C�:���2�9yk+H�Rr>���*� ���~�'���ſ�g?��۷��Ƈ��o��3��_;�C�/��:(J�p����)���ܶ�w�&\G����{����<[�3z�������s�^��T�5*�+�([��c�m��M͔�%�u�]�+� ޛ�q���Y�3�5�S�����x�0I�\�#����$�J��-�ػR1�T&�Vic�}�K��������B* A=q�e�49�$���뵫b0?5�����<:���I����cC΁3��Y{�:��B�j�2y�i�w^���|�(鐄�ri]�sf�������YZg��$:ߐ�8ǲ8��Lŕeu/�IKP��-�e;r<���$@�s$y���4b�# JAΕ�s|��|[��i� ivZΉ����Dm2���ڲ��h��ů|�����C�
�ʢ/� �&��("��^�)u'[^��'�Da�f�f�H��P���z����,����g���߉m�>�/\FNk<�y�����V�O�k#& ��1���!>|��<���*-s��4}�=��EX=�@HΊ-e�3���z>ak�|y�/o�M?mU�*���|�G�x�cT�Fq�1�t�t���]��ȥ�� n"J�"7N?�_�"dY��/��*�sL�H�u\w��	��U/��ï��P%EG��W_z����<F�FP�[hrw?v�;����?�{Ε����;��{���r_�7������^�|���X��+�V��u�m�����%��`{�i�ۖC9S;|�6��(K�2fӃ��x�o�.���wĝ�^����n����2�ȸjf��y=#������Vc��gz���eS272�	�\h��&�zi�"v�ޯ#em��|��/ջ��{��⚖EmʏZv��F1Ύ�Gd?w�:��t��f-����Lf��<?P?�Nt�;����o�-"�>=sI�-�"�8x.�U��{�de�o�'q���*H̓�m�i�>L��ȉ�,u�9����8��8���5w�8e��Ƕ�֍ڞ��ځ�9$c�=�F�!�U
�.If^\D6}7&�꼵ۆ���@�%{�r=���..���h�Nb${��woxr��3��QG��c��pz� �߳_��K${^�B��F@`dL�d�q��4��(���f��ĶEV,^d۔�#1�0sg��rJ!+@+��#��?r/�u���������/]R�:*��}�]�22�%���@^�,ɺk������
�9���u��%��bj�l�ܦ&Ao:"Ǔ�i ��q2��u����r�9�;f�7�)�t|De-���8���aJ[�o�h{Fg�Fv�QK%��!	�Ҩ�)�$���uy�TXZ����Xby$�^�`��Z9;��,�_G�&�_�[�R���wSA�E;S���K!�ظ�ߛ8gH9Q��F�
_�W��ȸF�a�3ߑ�˅��&%_�o���i�}{�~},Y��$H�\�d(���x�-�j���w��8� ܮ��1��.��cvau*k�f��V�2����`��_ ,�e�����#ی�q�al�#z
޽|[��_=��Gy�j�����{FYڟ&rim#����P���G�U��&�����{��P3 ������'���`)�\�Pn��J�(k�s��v;��.g�mf�1]���z=�s�aj�VKK�ZҶ� �2�n��<ri���.؝���w�Q��UՑ��_��ҤO\wOlAax�o�	�nk��������%�-&�C�u;��c[&Po�h���N"���Q/z���= 8�}㭷�Ƴ�9��>f�j>ĪG+�������\��{Og�j�l��?�>�O�".�݇��^�����3�'��Ǳ������~	U�V�/�b��8�u��������J&�Ʈ����ϣO�_S��3�y:|k����Yq���p�r�h�D��tղ{�X�����y`�l5$��h��Ǟ}������� �ҩ����Z��
Y?UÜUm.徃�D+��<l��&�VU0;���t��Ae��Fr��g��m�b^�� ��i6b�uQR�@l�М+%[{ ߎƗ�A���Hp�jR]d���:�|���63r��n��M?3�k��Z*��}w%�:y��8rBU���$�ey�\��/�2Z�ѹ��,V<��ިPRL^�/��� ���Jh ����I�4�����j�����L�������bz.Ψ�4H
x��M=6������x�\���3p!@�y��uM�F�<\��XV��sn8)ϩP�N �:B�V��?�w�4�Vo�<ft�z���J�t��{�X[�wKkX^>�-�\;O�I�����1�%�c����*�v{܌� ���4V���L�p��'��p��9ͪ?��b�L��,��\���Z?#秭���m�\���ObG����S��(�ߎ١LB�+A�� �m/������p�g~��!�M.tR�O�}Vx�M�c����&�&�����n6����{n�	�C��74T�{vb)�Y)R�^�U��I�	9�q	he�F����k6���wa�?+�I�&���G����P��'=K��#H&et5��sN�~���pz�t�������-ߏ�q�t�ZAZ!Iȍ����|s�+:�ǊE2��Ź%��g�\�`�W���
bꊧ�S�L�$`j%;��]1��v���	���ƒ�,�q˾2嶰Q'0(8���	Z��u��\�D{{��k�����Þ�J���TGcp,�3#u�����5A3��𕤥$����՝N7Q������x{�|/�v��=6�G�\U�h���:��L�+�ѐL�������4[����e%9�F��+� t[����+���ƪ��t�hM#�z��Y"Kͮ�M��Xu�����!ōe���5~�D_���}l_斖�Ϛ/bpxT ��cV�^O�� ����.��7��T���u�7�Z��e�CA����$�7lirޫ*����!�,/▽����ٿd��~��:7\��6�e��Ԍ�kO��ҚjۧX1!}��R�*!�w�{�T-ah�vdcn8^i��7vN�r����Ieq��FRC�(k�g�t��wK�O�Ѩ��$_j�Z�s ׁ�F�9@E0i�����gd<���s=8Ї�d�)�����ΑG;!�:fI�V�k%��[�2%%�Q�j��~!�2Fυ�S0�tD�]ժL�^�99��Ui���
Ml�V�\pd���1e�XE��l���t��_��O�,�I�>��aT��~�9��~C��1	v�iv1���;����j��w	]l������B��ktk6���8ݙװ$������W�W�����+�կ~ܕ`�џ�z�Q�<x�gc�kŌ��>�
���b�ݪ�:g���0�M�k�dF���\��Ne�+}���p�}�k���_�+>z�,D.��x��}[O��J���x~8��ل)=��6jt�c�9<N�5�aFfØ��W��[`D^Ȉf��O��}��0���=�b2KKK(�k��̜��,-P�o���^���	��4�sT<�L�kG,�n!�h<&cYk)9Ύ��k���%���ؚʡ��E�+l�"2�����5$���-�Q�����SH:m�v�~-��K�]���8�k�*@�L��s����� ��b���J	97$b���Rf��chM{�'��������0;��*2��]3�L��j P�C��8�>���_��(�^��</�������7v����nip�]:��Id�����ԓ�T�<VU�V�� |��I���n���[r|T�;q�<N�9��7��̩S��762��/�¹A�JP3?3��o��UmE�9s�^I��j%<��C����Ϩ��G�s���%�o˹�i���a�"5�N�ŗ��M��S(��8M�?;x�;��W_}
Nz@�_�k�2��Z�'��lYxʟ�+�,��z0\_>Oh�[����^��GT�	���&�:gНh���<�tU�=�-�d}\8v	�\=K��u}0�P���|m����&��B�d��k��9e,5  aBEn�-�܀��au��>v��-��0FF��8��co�CYVK]�5��8Rpl���ߵ���r�N�'�EA��\\ ��#����p��i�e�\�H�Sp�+ڔy����Jںm�[$tq$�_�@n���w�~�T�
���۴[��q��
��角*1ږ��,�&k�����Á����g�W�����J֋;����!-�Pd~;�Qy�#��u_�bm6e� �Կ�_ĂX�j�ZS�-{����Z_N��½�ދ� �3����˕��d:��{���4����A����GG�Z��}��:�m��&�
�8���*,����s� ����]g��i��3w��K�	|��<�6<N <��������[o�ѓ�Og�3��k���` �(�іL��2���&�O�Ր������j����Npvv�/)�^'-X	Ri��o��������oӽ{�;p��q|���$P�QM�|�ϳ\G��|���T��i�C�0�OQ��X��xH����B8��NG�#i���g��h�u?���hk[����z�~ݒ���{��kt�E�X�]_-icc�$"�S��I�,۹"���^����G�zU�zg�{���&gm��GԴ U��`!4q	?�ɧ�cݬ�ڶ�cHXq�e�`e�����p�7hy��b�I�]"��lf�a_0<���)�#����/KKӄ�e	:jz���}m]s�Ph�j^�!�&&��򘘝�Yb�t�	�����l�����
���ΟI�S���v�&�$sqF��O9I�g��f73w�����0���3��I��q&��;� �!{��
n��4�)��Ouy��h[x�q<Q+�����Cg@�c�+���u4�{����j`�,�.�Q���Ͼ�W��H��u�K���S0"��a%��F�Ա¤\	WI�/fv��i�Ï��G�����o�W�Ф��4�rn�*���F,v$h!)�91Ý��I���������u��>��B����t��
���..�c��^�ub Ö�'�i1��+ G���`�(&��6�(�q�Mj���C�H�F	Q��CZ;��d:��j�lA2r_A�ӊ!%��U:nL�$������<@�?��e�7�=+gm�c��Ɔ�ru�x:~'�i�����?���s��kt#�'�	;�JXNDl��G@"kY-�}戴�#]�h.]g_����~�f�&",�m�D*��V1���0�g�=�D���P%0uvK��w��|�#�e$K�f.=��dl$������*�dԉ5d�g�125�7��M���k^tB@4=l��,�N	4�4�ӳkb�gc��#�#& c��+Q-��Fb�3�쉲������47J�R�5�͠$�2-S)�����I��_Waz��{<m�ڿZ����F���cl,��q��R�� H$%c�����d�s��ei����}�1��a��~	~2u�\��@��ѝ���ź�S�m�����C�\;0Cq*dB�'��g����	�t��H�]�\�F��D���lw����۶m��)OL(�q~��c�O�� H@�3��$Pw�hg�Ƕ��מ|G��@:2ɓF��Q�hȿ� ���8)���O�~���`x�.�~꬜Ӵf�4heՅDF'�YЛ�וbC�zI+[@��\I��me�Wj�cAB�O���nc�2��hk�f%X�J��0�{�-�G:Y�mK^�?{}�L� �cf��O����V��.�&��M��^��$�Sd/��6j�r/��A�ȠJ��Ψ;Zq�ȧjL��d�C�a��!p3ۮ���	2bT���K*q�O��O��qҙ�#�]��&�_�[C>�1�F�:��}u~�#�����[4/~5��[��(��<�z�w���3��*�E3��k�$��!�D$�pw��[��&Ȉ�h�����U�:u
��9�v��DZ-SS����Y��.+��*\�2yBF��^ތL�����3)%;���"P-�(sR2@j��,S�0C`a?]��NS���X[_�d�i��y>k�J7b��)_
�$����ʆr��_z�(�"`�s���X�,*f��������p��P�r�I/�D�]J�cM2����ڋ.K�t��CC��c�,KҘ��Pk�1�顴�)�BX�3�}6��.�����4�
IV�,���߃�P��sɓ��rv��FC�	�����xt�b�jE�����%�s|o]���ez�N��Ē�d��	 WV��+o��ލ����Z�#��îJ�*`'鳶Q�,��\��ԔL��>ݿ�����=�H0p��16<�R�װ���
ʕu4K���%�-�'K�sX��XY�iL�c�յe|���cjj;���FV��6�Ժ�{�$��t�~�~��?��`aag洍a��>+>�Q:�����Pބm2������A���M���H�5`�i_����	�V.B�:UlvZ�D�����6��<��?p#�� o �Y��+m�=o�w3��2yo��{��}#f|���lAW��
L���c.(�����my]A���M���,/�Z�L������ԭ�%@�+�1����\���u��F��qtK^�) "�.r#XO$I��P�\&t⒠�6nV4>� W����^�3�	�%0U�|Kr3��]���w�Q�Ժ�BE@���a陁G���:�^#�AmYY.�C�^��9�L�vA�#|��X�{JJ��'Y?Y�~�b�E���ϟ)�"�K�~'�܎$��� f��1;��c{'.\@�����vt��A�Z���'�b��-(ulmwX�,��Rf*��o�,?��`$0}�jccc(���R��;{��jI��M���;�?��g���K(_\2R���v�R涹�C9+d����$�&��.aj�6y��ȱ���n��ĝ6&�
��pZ����6���#��C__A����3X+�uđ����e��1�֫�R������%Yq~���c�j�L��xgϝG��������!�Y]�&ᜥ)�E�L��!Oć��3��}�y߅��D�w������k{,�X��t[���M@�F7�O�U��բ13�W*�]�W�֯$��@��pG ��"�w$#�gɹ���'�������P�������-���J�Ĵ�RB\ ��Z�jK�.}�?���-7|*�1�N�+�A�&Yr.���;u�8ٖ�]2��z~�6gf�vkOp�÷�RH��^*,�G畿�X����~����7�;��?Ԍ�2Y��<{Ϝ��<[�f�{�t�Hj�"�z���4��,c�GF�*@O����d��s_$���น��Uܴ�S�Q#g*�[-VШTQn���{hl+��~��&�gfq�-w��R�@aP�*��>�����Y[á�q�C�!72�
yZ�i��X�i{�_>�����u[���K_��>vL��BY��\aD���uɂ���7a���{�(�L���?�&:�V���q�KUdG���
43�>�	 ;AC{��|�{ߍw�u I������מ��PA��{���$������3�2-���6�K�x���%�(ʙtpp�#��߫��c��#GN�w����!�C��޳�L�ms�k����^�
#�M���ytS���2��|S����V��:tr�1FG"�2s�R�c��@�K+��km��{Sln?��&�_Û,���	�d�`���2�Lt2�ٿv�$�E?��.*�����d<�e��w�t��U��2�&�G~�Q��pމ=`��+m%�u�_��1��v�6�L�	��w��#�<�{n����o�ŗ^W@��Z�S���Fx��`���ڴ�j�ז�s�$ +t�,�1_�*�Skho�xbYF3\����3��ؗ%�[�٘��!�<>�������'eAi\�����5ˉu_��$���O,ԐwB2�:npB=��H�j�? pĵ��r=e���sv�$������d����ĩ|2'/ZE�,��:Л��#��DY�<���Kغk�����ܳ�ƊWU�h�ɔV:���*�GX������{��i���~h�u�%�# ׁr���d�1Ɋ�p�-��ν{��V2m���|%j��?<�E����-I�-��L����#�G�S��V���|xt�+�����d��d�wMb�ĸ��-#r.],̞�P~����2��%/�x���"._��?�Q����(�*����/�,�$�v�F_*���ā}{�W^����X[��B1���xmNћ���ʎ�1za�A9#=�Sv8q�A�$h����j���nxC'�蒲:fY݌݌�ZaY>�ȑm+�W&�m�%�Mln����
�?�cW����n���͠���:�[�_��{����-o�:N�7�q��f�0e���L=�kz��Q��-�cc!�9l*�%���`ou׮=ؿw��b�����7
����?^{�fqP�9�f�f:�3h�-��^�\�E���jv��f�	'�S"���-}K����T��73��"P�?�">�|��{�v�p��`�5�������F���0��c�������������n`��Z*�@3�iu$C��������u��}��*�R�6�A�`��e-ٷ��)�L�Plv�ΥKؿmF���������/��l����5e,.^@_!��ގ���%s��_Va ���ٖ2��^���ڭ".�$������_���P"�|�V��� {�V���g�'��7���� 櫦=���+й
�av�=g��˦і}��}!ߏ�����Vխ���r[4xY^Z���07���_y����������G���/aeu�r�>��GQk����v:zBv�d���=�$=����pd1Pi;_%w]Δ��L��27�aM ��1�.烥x?���cB�	�z�m-˷u�B�X%�D���$?oq\�ck?���+�o���~���=+�����f,�c7��f�z��́w����{�<:z�*�B�H���kGci
��,zf�̐5���ģ����A.F$������9*��`Î�2s����g��#���cj�Z���跪���;/��<#�JE4΍7�E�+�jpt�"�Џ��-Yȓ�,%sƗs�<��y<f;{�q_��V�N���G�;هv�a;&�����s	�|]K��̬�g[�Oy�lx��׽f���������>����I"�4܎.mK4��pp�j�L�n��ˡ�na�(��B]��e�RiL��	�r4��0�k'�����b��AZ���<r�_��)S�}X�,���A[�|N��_G���
 �����v�ju=������N�����.bfi�C㘖,��N�.x�2��E��*�����``�Q��^+�X͡7_Ã�ނ��y�N\�b,�/���c�=9��ts�X_���N���x�,,��СC��ub^{�e|�cV�>z����d�RiG}��X�>�����g�y�~����C�� �u6�2a�<����6�޳�;D�����m@O��Q}#���q���j�.����� ���Ԯ�m��~�n��⒡y�I��������u?iQ���[ԃ��������ӓ	�̟�5b��Q�2L�,gDe������E�%&��t��hŹ���cL�}%P�ٳ�l?^�uZ��.�Z��bf�H��u��tN�N�N����: ��je�.�J�!%��l;���	d�����j�����~�1}f���+ƍ.R����}�?�`J��V;$��J�#�S���zη�p�2+��-g�|�}�$p���~1�J�'�s����X�ЏX/�r�.��dǁ��&��
�+���E��ު3�
c�(I�������V8�Vc��.�TV�:$x�VO欱]�Q�Y�{��$f<��X����1��}�[�J&\RQ���*��BA����rD?q����(����\��*2���^ڒ��Gw�@GK��t\Kϻ*H�R��i+毟zBݎ;�t:i�^�y����g1��&AbRU��>��������sx�WU�����Ϝį�گar�<��3XX_��S�'�YR�4|	P2yퟻ�.��r&xn=���l,$���k�W6BP�B~@�D��~Е�.��[*�fU��I������Z�RM�:�d����/N�`~�n��~�n��4�ӻyno�Ո�$�T�2���ds���hEi}/9��`�P9����@eI�sX�;nF0S��x�$p�<�ju�'LMs&±!WK�>Gz�ь7����|�^x�K�
�T%���7��4����c~qM�Sor���Yz�:��U_L���q��)��ؾu��a��y8�*�r��;���v7A�7s��z#�����1��T�B��q7̦i��y_Vt��KVEtڮ7�~��n��#�8ǯ OB�.����L��s:s��S��KG��6W���,��� �gnnV.~�A�B����x��y�����u/$Nu��l#4Bq��_|�9��?���-9g*�+��nv0�+(k~y���rm�ٶ�Tϓ�*
���ɨ[�CJY�� ���)����}�T}T�_1��a�2��9*)`��j(c��<	������'���r�@�>����/T�$��sx���}�'���ܗYN�ҟ97��g/����9)m;� ��������G��X�^}�}���a�q�-��J#9�<�1Z�v\C���B�8�����5���rN�^Fm��k��m�@��m8���)�K�cqlS~� &��^CrR<ל�`�B�͜gש/��VHqe�a��u+,�øm�5�ɇіE��G"�4n`G=�(��Fp���j5��g��3As��DYj�������~��W*�E���ܦ�˹�p�X�.��
3�d:���ӧ�W��|��3sR�Ϩ��H2s8.G��,v�z���%;L"��g���;�U�p�������ӕ����\=yp����UiM��4��� �*��A��4�#\���S��!��-��Ĵ1}���֝��l!���V׹�oa�TX�M�$�΁��]��ss$8*bC�*��dc5��؂�ot99��O���*{Z ˝z��)#��<9ɔ�y���q�;�?��_"ɖ	eV�
�X�P ��K`c�3"F�RI��T���٬H�+0b*�;��8�e�<�X�� áʢd�NZ��O�]ӊ2sb��&iR3�OMn
�Z�rC�#qK=�}�J���r'���� �֦d��[��$jP����@89�:Oa'���*��)cP�"5�/���8%�Y=!�3�J��M8ۯa+}xK��Q	��T�،��6k��mЯ�-�J�`X�w+mW�q���Q��^x�5'c��b�_���B&uh�	'�%m�i-�r}� d��A��!���}��.�Q*ѐ�F�r�QK��~���0ffԘ�e�`�(V�8z�4.L/t�K4Sk'�y�aVAr ���%���؈`DAf/�]k;���t�TX���6F����Y��Ƶ@( �R���;���lX�^�pfض��
�X�=O�(��^7f�1���ˆd��PgF����.�d�����DcN�w�0�4�9�/A��@&�A]^ϕk�}�8n:x3�����	E	�8q�H��4#��سw/�_���U_��
˾P�{��_�\װ�I����n��v$Q���!�g?�9\8�(�I��c�|��>��N�K�X�׿�N�9/�a�J	)���_��k@����Sq��9���n+��QB�'L�,-o/V�scn�Qπ����Ub����3֒ �.u��	�j�  �IDAThȹj��:�S@o)��
��|���Jp�e�O`r�v�O��Hg�@if��k+8w��/."��J�-��+��,�Cd�l>���p�K�~�XYO��6��o�m�5�������}0�"̂�S6�2Ɉ��-��YC�c��;���u�p.��f���H0�*��6�+�8&��c��"4N2�)�����u�-�����'�Ic$J<px�G0�m��WC �+�{��IXE�yd�(�p�BE�U�ٳ��,�r8x��h.-buzƜY����V���_�����F�˨JmW��pۘ���]�+���}y
�W�B.rw��7������&G+���a,mيN����7�1�t�Q{�4M^;WK3Q�`)1��O~Ǹ�q)`�e�����|�}x��q덻�����=�������/~��
v�څ���ؾc��Ͽ��Ni�D��\���V�ZW�K�L?�ɟP���)CHg�"�v�ݎ���?���'�{�����n;8�|\[�(HB��{�/�����N�F(���A+

�jc�V�#�Uҳ�2�2�mmQ�}����BR��Q,C�C�E��,lR!�DO���ΒwL ���L�����y'غ m�=':���`ǐ�G�g�no���?����{nEN,�#|Rr6��P+�������E�uz����߶kLZ������4�UY܈Lg����j��a@�����&�_��mAu؀Y�. ���^�Z�hE�l%�t�YhnQI��@ 깇����3��&��0�7��.��#2�6ݶ���M�g�bH�á�,j,�3�����Au�{6�S)PVFGS����_��.��@��6]��P	.������ot��^F,�h�(� Q@��ŲdQv��oΗ����Ǚ����0f��$(���J�+���E�} �k�V���p뭦D[���X]���{E�O��:o��%�^o�(l�`�Q���rMW�;5�Y�e�[�%���0s��o���Myuw܍���crK��T��@͖�$>����=<��w��c����I�)@�wo��d�)�>�*D.�ok�8P+�⡇ދ���"���l�.���mjn�� ��������x�?���Bm=���琐w��� `����~��/�\�_�a��>�e2����l=������һ�V�Tx$9z�{�H�Z�5��4��}��J��j���^o�դ,p�l9)?$mڪ��L5��`Gn�f�,竃%���M� ըg|d)H[���Q?�����ѿ��?�;g.^����[!f�*ψ�xz��c�eJ=
�N��]7�&�_�� �O:3u1ǺJ ��e��#&:7��Φ��̫��ޱ߰M�U������L��aZ3���%�i��Ɍ L� �*=��P�d�Z��^���[���}�C�D�}O��XF�3i�����h9>��� 3Z���v�]�}<�]���{|���~�9�ݾWF��Mi��}b~�B��ܔ�d�!��C�ҀM�y	l8j��i"H�s�����쮉M����̲V��Pa���wɠwNM`�4��կ~/��2����O~�?��n؍��n�� H�N��E2˜�G� �jP0��q5�!x��λn�U::M�z��x��W%�p�-��@"�W��J�������?����h�/��~���9�sם�}�;!i���jCҦ���nU&��PE5�rm__���1��rl]i�I%��Ѳ56�cϿ�/A"�7hw0>:"�	�|�\	4����k����\/�����ߠ����a(yГ��-@^-���(�Qo�u�;x�ћ��/����_��ҢzУ�=�(��#yx���:c���M��
�l�����&�_�{�@���4��bsE�,Ѣ¬��)/1���=t�q�~�R��a隙s�zY�����*������I�A��1d�tʈȘRo��mޏ�x�#X��U��|�����m8{�2���� A�N�
f���Q�F�y�7nl��U����ZU$Z"a��~-$8E�-�74�"1�1��ma���?�<�Ud�h�-�G����+������FV���nY�Mn��Ԭ�d��IJC?���$[v@<�DfF�T��	���5�r9��PSz��N����Ob��D�U�o��_�C�`ny�.��/��W��ž�����#hK�e%c;��ݔ`��AF��^����8}�>�57Zk��?���d�g��X)�%��+���/|��8��謕0��`�=!sX^]��AML|�q�u-����{(=��J�V����9�� �I0�")��T\�F�-��gg��z��������^{G3^�3�5�ږd[�hRb� @�4:w�9V��~���A�g}<�LA��f7�X��������QX5�$�Y�����(�]�
�퇼��@6�ig&��`h��x�*�0Kr�Q�*�ҺQƆ�Dw�}/�ݻO�y<���R=�8���B��mfMRY��]͞$�F�:V��v m��%��׾���|=�"n��V�x�^t�"䭸�[��oވ��y�BŁ�	b�������v�U%&�/��b��P�eØ�C���&�F�J�� �щ�n.Q-�
��^D����&Ʊ]���õ����A��4M������	�q�A�sk4�g��s<�e3�c����=s�Ie�[ZZ����^8o��Ν���!|��o�C��x�DBL���vݤ`R���K����hty��L0�@}qߤ`ٷ�{.����Lɾr��u�|m�3��5�7ie� ��\��@�7��}�ɨt�'6j8�����u�O,�'+��;Hgkg
:�\��҉�R��	#�0�TYQQ���;����}�xuH�SD.�.մ/>�ͣ.F�\���`����z#I#���R�J䘤��B�z]⩸fNRb�� �"��/^�uQH������_��Lr�wc�\��+Պ��ށ>����?�!�~��t��R�|�t!�ڢe�ry1�\#m�-_ʹ��䆰�():�lW���=�O�^oE���� t�E���h��.�Δ�����Hdr��ƛp�����o�筈��Z������1dI\C�9b�3�@�$0?���33���[��g���﹝�V���Q��*1����EoZ�Qh��].�rmx�݋Ŝv�Io��\E��n�7�2�!���uZ�,ch�Ja�Q��4�K;A^�6n3���R��/	�r�&��87�U9V��ɇ�Y!{�\"a��9���L�\G��mjv�:f����v��x"ӥF=�Cےs#���m�tê�tH$�s4-��x�U��V\�'����@֎���9R,�h�������FK�p��	#���p��5-a4l���v m���P��Ip��&�����e��Ǌ�5����v?���S/���I�f;�~�)h��M�C�blز�2d4�so�`�٫S�5~��v$���U�W��[�9�
#Tn���l�,1��T͎����w�7�#J[�x����kS4WVFU�����ܢꤷ9�	ꚾf�����<ӓ�Í�V43��0�?�,I_}�N������ǖ�q\\X�����Ǐ�7�'죺fΜ����;��=�͛��:	[�!&���x��Ғ5�@!�)^�:it �0w������X
i���V2W���j0UMz`+t���u�@�`��1���-���_;}��!l��qk���`l|D�
e?�N��?-��:vLq
��`F���e�p뵻1��A*]����pߐ�I��M�Xu�`���%�X^���69�&�?�zCCh�g���!\��$k>�v�n*ߨ�_E��n�7���~���^K����
�Tlý�Ճ���1Gd0��d~*�u�>���@;�Qr��������z�^2�VP���%�j�jj��� yM1�Ů]�pn�{�wm���q7�=X�HcY6�/<�μ~��-��9�ѳ�Y�/'f2�y(q�P$F�!xN�P�%��u}\mˤ��)�jx��+ I3�������x6�����Vt}BX��o � ̵X�-�u��������v���m�QWyW���;ơR�O�Z� =ߑ?c����$"��Vvu��w�v�5�B9]��`��0$1���htH4F>����9d�&T���qrB:�奊���==*�鵺���zХ�
�f1��D�lAY��iK7������4��2r�]�k����{�{���~��˿�v���?��Ͽ�uh^�xh�U���)�궣4ġ+C�[5��
���a����4��W ��:��3��]&L��n��qi�}���R����cb��������v��{�!NgK�.p���*�s	]�X�wB��,��B~�%��6Hh?>���PX^nb�����w�/��c����n�|R�R�V1:�����_������E9����>���76R�o�v5��]�r_%>QiN�"����`}/��me����Z]S[��j3�-S�ZZ��q�NL�1�~�<*���=_)G�b�J�ʧު��l�H$�B>��.�b��ú�L�D�Yǖ�I��`�5{�L0S�hE���_TjF�A�fR�x��P���Ez�]E�jL��M�sF���Ҷ�� (#[`�k�:�D�zq�<����f�����jh<�b(���K�0{פ���R�*��ot�֧��8_��j�u�=���2F�m�h����=PyΖ"׿Kk]�f��ߙc�K�y�Q�H7!�:77�RB�Өc8��|i�w���7�Q���o~S�oU����))Z�ߟ�a�KMմ�F�&�h�U�kd�eT,��e�.��k�v��C��0��=��G�W(:�r�M���>�Z����,>����g^��� �!s1so����[gnD�&f:0!X������D\�m��Oā�J��S؎��F����v87�(?�X)W�y�aF�=>i~��M/�o�S�-|�	��<�����}9�]��h��ԓ�#)s���y,���ӟ�vmˣ#�F6d��[7e����˅=;cx���Å��%{m��m��\Ecà�I���e[WlLkG�2���#�@��mJ��o��M�l~����mѸ�-�D��#m���G�G�����9�����Zm#��S�Mv6��I����f�gh I+�k��Ħ�	d�3]���[���Ӗ���cf���8����іM��&l��x�Q��Ɯ����Ɗ��00�-Ɵ�\fÎMj��QN��zMT|F�5���)R��g�+����l��n��Y�2)ܭc1W#o�nR��+Њ���xR�)|!���f6eg��m��)���#|7�n��>9�ex=��J��(搀�{�~�x�El�{��~\]?�8�ԷQڎѡ~��n��8z���-$3Y��j�����w����������7݆�E�����ޏ��AT��(b{`�~�����/C*��O�֭[�s�~̯T���xJ������;�N�
�7��#�5ٖ�G�I�k�2�:jeժ�B^��}�}a�W�#��x?����%��{@�_U(d�k�}��UD��뼮�"�z�*s�Uy�T��N��\I;8�{��8W./"�)ஷމ�_}O<�\��d�r�m6�^q�/d�Xjh�R�c��.{x���~l��c�Nsà_Ecà�I�l*���b�9Lˌ����mZO��}`4�}��*R|_�CBߤma��ԀY~*�ȺRx���)G� �ᑗ�-b�#hmaqYH؂��Y�g}vi���~�=��|O?.]8�9�|2��SS��8{�2�^���!��:$@!Ŧeк��)3\,�ȇJbK���%T!�LЂ�Q��ҧ��&v ,AD��qʲ�x���ǉp���F��ѱ��I]^���Ж</� �y�@���z�Zm/����������5UlZ;l��V�5g/W:io@��YqY�ȣ�RA�Jr�^=z���D��;�k�M�ԏ��]1�/>uH�a|���5��!v��퀂����/`�s�5I*^��ìI��?�ؓ���wc��Mx�����iʙ����>��>3�����b�?�۶���w��~2-��CG>�s�[f³�~a@��\&r����|״�} #sXѴ�'�p�����zPȦ+�K,�RVދ�U�X�8�z�����j��~�L�%k n��T#�^���7��_��V�kwm�G��.�'rb�\�>���Ͽ�5<��A��®�֨�s�p-�Q]�`Q�F��x.����������ƆA���ĺ�n2j�1��֖��h+-�ư���E�9��#�un8���kz�a4���eQkT�iE�"�e"���\%6	�֞���8b!��&���=�'�|R"�
iX�"y"�ٳ�c��v�8�;�
R�$>���ts"݇��1<�ȷ�78��zS9qn�ls�Z�R���5���py���c�#?��� ��D��e�Uy��9Qp�򰇘+<nִ9�����(k&���º�~�*�.����W�+��iպVuW���j�q\`����fF�+5Q�fE73�����.�>��sd�9�e�d�U��w��~�?�>����@��~�/��+y���Q��ѱ�Hz1�Xǥe��]��bxx���*�C�����Y�?w<���a�Ͽ���s��?J��G�.��\���
�z����c���O��n�۬��um���%�+�W:/�]�d�|+j���_�da���jTn�s�h�Z�r��A��v�u�Sg���r����[u�>���e��q�ѭ�!.�*�e2���+�Z)������>y9��g�a��$��:���a��O�؅9��|�,͡&�
�vo����2�8���R����-6��}WzA��3�����M;�JN�pc�ͣk��`M%�E�����*x��հ�}�#�&e3h���a����� ��k��<2@�_��l>�iic��3��&�-<xP�L.�+�SC�9������I[8vvGN_�RI���^~�q�e�~����@��B{�".^�VJF)�x����(�V{�-%�zqy�)�i	Qmx���w�S��3�G�o�pl����l+B�G�����kdz�#!�@A�mQ�=lsb�B�+S�Vh�ò��Κ�u~f%�����b� F  (�H���I�[����_�Js�댓�MȒW��PizJL�v+�j���q���,����+��Q*/�^� %�j��_�?~����R����T�����ը!�̠Z+kƦ�ۇJy	�������F�Ѐ�$��L�n˪U*������7���M2n}w2�eӘ�U���$�&r�+����
�s�.F���%h�<0��~�Q1��AHd�gp�t�Q���Ƙ��'�:zS���wYj�k��]C���V3Xz�yb�#����"�-���,ŕء��=;u�2F���g�N���y���
}צ+��Q��,�L��l)um��fxe@9�NL>_�]�'��l]���bc|���:|à�IG[�@஑b`�|}m[i�-k5��*5�I%3
��W����Y��;p͎k�wd3�6�L�����`t���C$�bRz�;Tr5�����k���Hi>66��\����y����fW����"��8�������������(��K�b���N'N�u�C	$�y�ܗB�'bT�j&�-i>��r�L��mF��	�� ���\RԿk�WԠ���yhp@�5Ӷ�gnaK��\���'�:��<+�(���Qo`fnA�<vD5xq&\���8��"�eS�[X¥������ҕI��%8�!�(f@��а)�|�a���b���mhj��8Z�z��H�QjWU*4����a*ُ�*�WR�A��bvev*��fx�1ô�L��]�������2Z��v��%�J��ճy+�e9��r̜�V9Q�L�X��e�U�#K����x�g1�����o`k�*�ax��⦬���c��i#�����L�Hj)�\]���CS�o����Ǣ:;32l�dK�͆�@��)�g��r����~��~7�U�^�������l@��슏饒�'�Nbܘ�9q����:��OM�[�</�%~�㋃��x��o�~����=���
��V�^/�Db!��x�	9�D���FI��r������^C�� �ݷW�|�F��q2k1:��H�)�p��3��3�����n$%��k�{W�A�\�H0*%7����1�j5��\�H�����Qk�T��`�H1;2�>�a8p��V0�\�|�Ҡb�א�(�*�%�%{�� uɺ%�C��:M�>g��s�<'��B6�|O��o�[��{`�6����G�����'�F%�j�U���j��/��J���_����������؃/|���/}Iӿ�.ݎ�IA�;�t��O~����k�ʫ��ۿ��X.�5�m�{��c�I������S�DS"�t2���������
�҆�Ȣ$d�f�g���D?��b���R�1��xL,xr,4���à��@�35��Y���K�L_~"�g�$NDV?;����vT�M�����nr�����:W}��Ӹ:vJ��k'�/�+�q��9�%Өө�Hګ�~�tXJ���툃��Bq��S��J/��y��:�!��cC b"��XG���,���+2�w���X����w��չV'��M��:uq��J(�T�.OB�$��@L��zbtI �Зk����7ߴ+������-?5����7p|n-%Q�E@̓�"0J ��L��q�Z=#3��Tl�X�{2�Ɯcà�}��ㅶ[��ůL� Vk�
���'7ߤ�Q��~��1�}�]wi4N#O��?�����M>��j+b���O��ߺm3n��V}����^�S���i�2ijO��Z�D;+hK�Q�s��KG6oK=/y|���''����9���F~�9Կ�k�,"�L�����M�a�m�;u��&b�帺1
}��t]=:<h�<?4 ��lߡ��c<u�4����X]�kM�n���s+��(�غev�ܡ�NӻS�V>����;�Q}��֢k����
=��\�2���9T�]8=�wM��"9��3`W�XK#u�f+ [�|gC�F���wʜ�x��t�a���V��D�I���1����mӮh5�N�7\퉴���!4W1���Յ�[l]L���q���,'�%=klq���&��M�quh��{=a�I.�g�g��b]י�� �(knt��U� k���9���+�1���#@hT�
��{�
�z���y�h���D���( Ē��Z�Ő��t���ٺ��D�ܠc���E�ja�h
Uqz���O�*^�������#��ك�űJk&��r�Ɍ8{���:f�� �f�jF/�%��ԩs#3��\���?�cà�I����^/�bP��Ҩ!O���,��f���Ӏ�zY���)��iz|z�h���������O�LÈszzڤ��`0r��h:qқj�ö������`Dx��i{��a��ZL92��n�Ġ�%��0�M�p%2���A����:s�wÖ0O�ӼР#0]�Z����0����(g�[o�O~�#� b~y�<�u4�܆Q�(�s�uyq�@�i�� ��`�΅����s����W��I͆����E���y`*��r����cf88��s�!ժ���%4%j���N��Og�>�
w�Νp�\Xib��P$�l&�[XG�5@�v1�Z�f��]#�ܓ��itN�/s��T;p�r����ڥy-�xIc�Z�+� ��"�zWK���ݐ&�[�&�i3�:b�T��a^<��x�:lF��e-:��g�c���08�����L�q
��1^��2�\c����wvp���������_�������qtV�M~wɕ`��Wr�%>�Q�)�qL�w�>�\��@#zR�*�����������d�;U���j�'	%w����
�O�CC�T.���+���dI�m��^��̟��Q��d���N�:3t���a9���W���3�o�R�����J4�Z�8�Xo�i��1�[�@t�IsG��T����QT/�Ȁԓ�a:a�[�r���F��cT{��r*�>�^�M�b��GG4ҚC�(�P,b�����j��L����)*��\!�v�FRSf0:ז1�� ��W��t^4j]I���5����Kf�lt��Mu߾�q��Y\:w~ז���5��-[��TV��q�8~*���~�9v��3(ʱ�;��=^>xH6hCʾ�.��T�&���8#�֫��@O�O`�҂IM;tr�J� �xB�gϞ5�}1��y��ob+���ţ/��ɪ�J�Z�*0n}�!���W����m�.�	��:��G��)Y�Bc^�5��Y����֔֊��&y���=-?�q0�h�2f���;#��ԝ������2���r��j:�b��ℵZuMWe>q0Y��f]��63P�(����ZNqW�x('��72�Y�����-��mj!���gW�2���]#�YwB�۬Q/�}�����2���9c	��`dh�f��S���uM��vR��2zǓ��vu^�D���g�]��N��<�L���q�B��w�.(�La��8h�o4�#��s@J����V�s�W���3�?ƜCn�N��,�����`���
QҼ��uyDn���E��
��Ɵ��Fܬkk�&���Z�o	5�)-L�N���s��'��"JS��fۙ��
%�$'�8�h��5�XY.�km1IR��N�&{�؃d<�����i��ۘ�k?j7� jP���2K���+U$�Y�>uzK�Ue�#��Qt�w ��2F�7�*F��\2�����b����dd�,��tٚu�}o������Sᗴ���H�\�i���Ԁvݖ8�q��܂�J�^zE�ǖl�9�z��ԣ�g���bBJ6lFc��7o���oCK����0B3	G߯�k�
�[�bh��eMݴ��q��]w����	��^����r^<y^s��J	�n���| '��O��J��D!%�����'~C�CLw̸��DT���)oK[��r�BN��Ya���n�=o9����r��o,-h�CVe0�?h5\_z��p$���ɖ>փS鄂8UgՉ[���5�v�٬����*!��7��^$n`�S�!X���a�s�g"�rMye	�z]Q��Kg9LfC^3M��ŽnKq��G�+��U�!���(��N�ٯ���.�x��cG�)����8
�V[����
q��y;-k����A����ʖ�w?(���n����A���˲yv�΋[*=�}gۑӄpUC���
����Fh0��L�j�S�w�װ��ә�pJ���{���T�e��لF���F����߿�D(���������:���.^�A�D���M�`�T``�Tb�Vk���Ȝ�j��
�*�^%w�6e֗%�{��'�N���cfv	����ؿo76��*n�1�׎GI��d&�T�d����dC̊!���1߹cz
y��6f/^�l�x���K��O�˟�W�b�z�}bp���Kt��M�"�_*Up����)�}S"��D�#�[�H�艓����#� ���������%}/�O�A'fz�=^�hy�sg�e�y�@�c��<��|7�x#n�asUyi_o��><w�?�T�Q�f�sro�s'�~�NdS|󩗰ȹHgԠR�ִ[0Ң�<b�/�E��Nf�@渧��'~�c�2>,s�|�D�b�b�v���ki���M#����0�"�%���_�kE��+%`A��HSŃ��.�7;TI35}�����������ii\]hW��L{��V1���m5�D�S�֓c��-����5n7�&@�'�=2&Ⲇ��wH���q�����;OR(���^7��|���;G֗g��
��<1�r͔N����ct<������^·cW��{���٧�0�o�!��m�r�y�9�X}E���֧ސd�q��Ɣ�/?Dm�(���J���b��-1�I5�9M^6~�4��U5Fޮ���b�S�Ʉ����
 2bDL����>%����Pq5Z$��`�Nf:��יLNS�]�h$dk���4�j���1�=Y��Y��w;4h&,�rx�����_��O��/���e��:���%��)�1u�,.\��ё	1�i�������޾4�?�ҋ���er�~���g���Onުt�ݖA=�ܵ�g.⩧����"�o���O�:��^zI�������RU7d�Ė�h5�8|�Ҍ��i��������u�FF���������P��j`�3��Gx�ı�j`h\�M`i�����C8�X��G:��_±W�r�1�i|����ک�=;�)�b�6͈��m%��h��G�:F�$QiQ25����#����䱪̳�X��אy�U�e�� ҹ��$�,��������=��\��JȪr\�B(�յ�݌�oElq�d�����,q�`��s�|޼�|G,�o0`U㔺��we���U
2�Q��+��-�W[�脶H�2|�g���K8�O��R�kֆ�{�?t�:Oy�����:P��e�ƫ�M\Y�Y�G����F3��ѫ�d��o1~�b�h�W���y�6��t�ر�=v�%��o��Q�	��kr�~��ζ5�M--.�AgkZf󠑱5zg�Ϥ$ru�hp	`��A0��Bn�IP֠���NǂN��n��eR�Q�W��a9�hE�>:�$�\����?��,��INR�����J����l�!�e"uc�l�na4���N�s�A�w��5��4���I�XB���$zd���� D�؂���h���ʒR�Rδ��W��;���8nZ���%ȉ���Q��^B�R�Tz"m�(u�ĉY\ZA:�+�U��A&�F�������'�;G6mBeyA[9����ժjv�+ǘ����F�����<��F� ��;F�\�����1�r�qX���C_�Ï<���V#�F{��Ϟ����ǟç�S2?��3�9t��s$����
e�I��)b<�k�wT|D!p�h���� _`�[G|���<a�>2�q~|��u��V���f�LX�/�A�/��P"���Z_ZS�~��皟�XST_D���k��F�Q��=���+J_�EV��`��/x�Ƴ�#�B&Py�;r����"ɑ#���eH��i ���%��h*���>q>��Vvl߬���|Q��6�9r��
r̺Uk8z���oqY"�T��ۆ܎�Kt~��j]�WecH�~���i�9~��|à�I�l"���G���\�����ш��4#�݌52���r�Onٌ��q�~�$fg��06�L�n�ͷ�$���4S�u"�[�0=�P���.V�0����60ö%�)E"��yٺwi�ƍ^7S��:���H�H��f
��c�S�U�7���­�ߢ�f�{��-7;����l<�7R�J7̣����JȦ�4+:)����E2ߋFI"�޼l�),�Z����p�m7�y602:�J`S'N�t�6�����;9J���ضew��-M6168���\#L_�$�'��h�n]�sVAY�`w�܊{��V�f�C��f`��%�6��e�kK�($EuzQ�ھ�z�{�]����/yY����|~�)��;�rK�F��;x1:�?�:=�d�5��zM�=I9v]�?�Гw�`�6��|Sg/�ӱ��aY+6�Αp;�e���GM]�Ņ��t&Ћ{6O�_�j��|�$�}�qq�#&Ɗ�\6C}��*�\�m ���+v�뢧��zptN:��\#��8�x��}�ن@'�Ω��T&��GQe���<�4�ʾd+s�囒KF��P�%V�o�E��Z�L��ۨ�@�Xv�u��O+�NW�����j�b&J����5�9�ʝ�t�c����D��hiq"�cC�z|lod��T6�ZiAM�H-�9��q�Y�N��\�a4�ܩ��|7�q�~�(;L0]2_������@:Q�ƸjƆA�j�|�T�̤R�d!�7*Mv�����+�H�\��k�~N�Y$�Z#�k�c4�	.JgR���ڃ:Q��h����~O�С������2�zq�ʃ�hMD�)`,�pqT�%=��6c��	�%�d���iQg$�%�e���|�o�&(6��8�u�i���	r�[$Ea��;F���p#��<���T��]�z'{�)���k\���b���%������SO�ܦ��w�O��2.\�U]oIT�Jh
��l�su�m��C�:��D��{�{1u�<�=�1;�,��\Y"�y�w��oƥ3���-�^�se&��5jv�Lm;7D�un�dL�l@�>�5M�6�C�\�LC"�?�韆��7q~����Y1NqL��O?���1�iX����
9ܼ���Go�_>r
��G��+�P�e�޻o�G�{7��o1j��������~��4=OG�밤߿� ���Hq+�T�VT�t��G�i#�C�dd�a��2Ii1Y���_h@�z&����}�r�ip}�3��M�����5�2	�>����3 P�Ծ�-��j�?`XތX��3f�)I�T~�+�M�5�N���j��a� ��k�s�2҇ݛG�����C��A�i����8s���)�X+����uS��ՠ�e����'�&}�'�-��(�m�I�K�!R�&Z�ٻg[��M<:������G3��f��Gzz��8R�Ӛ��bu��Z��SFT6���lٺ	�!K���T&#e:�n��5-��i̍�sFe�ld�>�T^�2���ڏ�k��:b,�U�ϰ�͖h̴ر���v-��%"K)�J^5��I��%*a�T �Zה{`�6�Ht����t|(���%Ҏ:�}����S�fD��k����nl�ؤ__� ʵ.JՎ����z�o��"Ё��E�)��)� ��|��3Q#W�|N�)n�w�?24�ƶ�J�39�	�tV7z
ذ��d1�F0��bF^w��1��碐�"��)�ѓ- �,#E�'�`~�M,4RAD@$�(CH��ɚ��H�u�taF�獸n�6�Ҧ�����&G�����س��R��4�t�"V���W��JI�"���s�0vM��ȉ��-���ߍ�|���9e��,x�����3���� jI"�c�\��u+�#ǩ��DeY#b��ηoߎ���d֔~��H�N�3�ۮ��kb�����������3�x������Z�>L{���ro`G�t�
�ut��<C�=nJRkN��6��K;�4
ٌf��m��ක�q�M��w�d,��˥EL�x)��l*���,��ہ�:X���k�����O���j���k����8��\[�B�)��63�B��{4�>@#�.�6�m�ۏt:�]�N���Z.�Z�*�)굫��8�*�� �MtM������H�72�ٺ�'ה��+��筎�_˖���FG��:�Q�ԋ��a@Q161�z?S�O6E*�H��F=���bl(��8M�S����$!�����+h��e���G��a� ��u�;0m]}b�����'_�ɩ}�]�<����4��uE�~x�$}ٷo7����'p�գhP^���C�bVv^�dvE�fI�R^�T��Z��cb�I�����ؑ�X���w��y�nې��o����{��9$�mE�P�t+����A�ϳ��aT��������|�XڋH0�kw������{n�*�7��oڇ������%ʓ�*3u��G�xM-w��H���3����ކ][���������)� ��|���[������������?�?���iͷY�b�1'��
Rr]��"2���(�]�W��sg��z��]���3�����apq��=s^�c((�U��4%*r�TǞv֮u�D�����wD���:��q��Y`�vW�������K��KR^�N�em�%B��QY�R��F����%:/L`�5��|�f/]�p_+�zO���z�9���8�Ģ�1f���6ku�w�7��&Q-/����]�8de`�S���T7��j|��Ëg��3f���I�tF6�G=�{��{#ܠ��c:д
��d�b4�t9Ak���I��9L�ƐtXg4��
 c=�w�y�����¾wȅjm
4�\d`z�٧��=�ds�o��^�G�e�Z��J]6�NS��v��e�[�H����:�����j�G���}U�"��8��-rhT�x��g06�Wєx*� ���!�S����&�� ׹��佽}jܩ Ǎ9!�T��=����[�h�2���Up��9<����Ȟ�`�T�Z�út7.� ;�b�R��ҒFZ��ӈ�J����ߑ����I��F�-�	� ��	�_{�)y�>�vb���,��/�ʯ��~���ΛQf���H���L���m�:u�~��v�����p�:w/�x�n�Ce<�~)�R��qa�j	�ZV��|%�ZH��J���K#>�e3{ �4��TV�=��Vg�+_�*>��Oh��h��2J<u1h�3W���".3,�,Q����ɚ�<�ݱ�Vu�h�m��+Q����>�F�ĞҬG�0b#c��=>3�������Ѹw�qEEc��2��[�h�vy�4�VXc�:��L��t�Uf%��R@E"r:����R��5�2;/�3�k��6�i�o�ѹi3�\�A����?���c�f�d���u;M����k�
"RR��F�͐�V�(�Y�f�%T^��՛�i:Fj��i�GQ;7.��c!�F��(w�')��l��-!��m��4�Wђ@b�U�Z���5Yu5�LB:�ҍ��4Q�����jk���z\k�Os�Qn����'W6�{d~�v��S�֑"��F4Z�o��O}�eu��y� I�r��%��=�m�F��O�>-WZ����x���qڻ����A�9r�C��ᆛ040���y1�'q�;ށ������������h������.^����[nߏ��>��0u�v�މ�o9�щMF��}��.+�6��D��0�{��2),7�N�О�f��n����'ը����2!ml
��Z��%�3�K�dZeobT�#x葧�i���߅O���P�cO;��_Y��[�Myܶa 8@ǿ�Ź���|��q-��a�f",��)ɏ�M1^�W����c���w��oҴ2��7��,3(ɑg�;���)q�T��L�a)�!���G�uk;z�jF��WחaH\�W!_A�,�q���|�8�L�V�i��87U
�?�֤1��<7����&���(�M�^.���Yy޽�}��.[�>u��A�����JY�ܱͺ%��|�l�k���3({R�))�/,��;�4 �X����Y[���3�)�7�x� n�+y�;�ʍ��M͖�Z��H��0+!�ܨ����Q�l5Q��q��ƛ^Ig(Z�Zd�Ǽ�nE�~H�iR��U�j��f��.z� %Rj^6;"�#RF�d��f*�F�/���bT"�|*�h�x<�7��g��c�6=��:`�����f���x�7b�b`:X������O��p�;1<؇�J�|�-b�o���38~�~
�L�U_�x[&���(v����G����q�wh�5sy�=�
z�y,�M�YY\A�DH��xǽ��A;)�
�����"&�<!zU1������Y�|��O�x�;����_S�e�Q.�fe���0J����'�4j_�%Z��J�80Bk.��?8Ы�/K�=��Qd��Pj��"�:�S�\F��[w��m`naQ�q�Rhq����s_y�c��}0���!T�U���c�vl޶�b������xi~I��+����~rJŃ�ھy;f/�+��Ji	�ϟ���fff�;0����3����!�PC-� J���5�M��a�d4��C�E����V �>`2I��Ӯa�KW�8�V�V�[/�j�$l�p�ug���k��\��e��1M$��D<E�=�<��b��G����ڐ�fdNG%��cӦM�C���s>~�ͷ��_�����>�j��(�u�2{"�355���[u^�3??�;��������Hcαa���c��Ł pnq;�~dc�ѕ�J^F�ð�y������W2�4�����<��Nd��R���&v;)3M2�E}�*)n�Sw��h��۱4�3uFy]�5�3!�?�
�:�
�Д{C"�j��B���&�'��dI���U.z���s~a�uW#�P��^3�f��oY�����=���_Rk4��0�^F�G�ڡøtq���% �mNm���x���@M�Fr��d��D:���N_��61�y��LZagvE�3���\�v�eL8�����7������1
�P��b}�3�X�6�+r˖-���tq}r~˲8O�)�	��4 �(�3HQ���o��W�]#lB���+�"�7����_V�EDУ	�|&��7`��(����?�pt<:c��2�8va����|�z���˫�3?�O0(���RSiz���obvzV��.]�,�����Ϊ�,[͘qb�3*�#?��mƵ{vj�aY"ϊ8̮���<ϋG+�����n�`��� ��阯��M�e����Y�R7a������$z�
y�|�l����e��:��)R�2�/��qNf���Lʽ�&ӏ�G�=�a�\T,Uk݄�n�S���Ź�n�N	k�=���������%�5���vb02�=
����z��Og6R�WѸ��U�367W����=�����l�X��~�Z�gڭ�-�-Ѯ�v"�m[ԖN�����0ew����4����M^qF��,:jC�O�b4;���m��]�vg:��k6�͈1%Q����o홗�+S�Ÿ�T`u������&q��]��Q_Z��mQ"�q}o�1ui��!��WG�4
�~sM��(�V ��)W�����8��u�($�	u�x�y;y�8�����al���#>�n��t�os�x���˥��./.��+�⫙��?���f�CWk�3�!�=�2�8u�^��;�/�����9��}��I�+�@��Y���$�%0jmq�^;t�Uو��)�T����%'+�j�q�����E�zK�/�}����ډ��~�?�3�T���H�%�hF��,�Q����ۅ���޺	_?/NH��t�����W�//�Gxv_��0���1pg-���2.]��V��%�J�,u�V*�g���[t=��:��n�A�+^'�9��o�)N@L�f��כ��k��x<a�&�*����5yάL�����v���6��kM���������j��]5�JkaL�P�.f�� �f5�{+T�#i�q��1�up1䫎1���dq��O1Y����ik6��R���ZLLn6e
f���i�V���t&�#G�h�Zo�c',-!��Ԡ�<y;�c��-�Ŭ�J��!�r��Ϡ_Ɯ�\.b1��r�t}*�.d��������d2�����ʦ-�,��E�|;�E6�-T/#�z�bL��P\cI�SO"��3�͔'A?i��i���'Ƃ�r3���n�ʒf6�6��TN�V�k��xJ6���S�$�n��٥���̒<�b��.��:����NN��[�B�؋!�+J�B�45�G
��O:d���HY����l1G����a��Q1�+��:+�>�:f�5��@����$3���59�:����I�~��e4d�z�%L�E�&����8:N�<��S��e�l_�"����̪��31$�+ެbbl��_�9Ή��%���5�	��~GN_�������Մ	^�XҴSOL{��\�h�:��r�]ȧ�$�������妫��$I��� }*�$�e�.�#�O)���t�o�Wb~�4nؿ�������hV+8��Q�:vZ�P	���W�!ꨜl"���]��裏j9!)�[�r�f=�gf���B�8Y�i�<;-�@M{�[��P�[�bT��	�hD�+Qg��	v ��C�1��Fn^�<�`���!iL���{�N�u%������uS���Y�/)H��Qx��:���� @���I�f�=(Ƙ��T&��y4�C�شy��S]���J�J�u���%��gLLL���ǌ�#��'�TVH:9��0�f~�RZJcc\5��3�Wɐ�4&�� ��ݮ�4��B��l&����`1�8/�&l7H�=�8���s�/�mf�TKnl�w��y�q��`/�dؒ����rHw$R��'�	����i�	ƙ_XZ���WYȖʲ�^?���ƪ�ħ�Eu�=*��%-h<���y1�I탧���EK,
k�l��}ݍ(��"��6 9%���U�jN=�f&A	U���S__��z�t(xL6>���.,��lc��Y��4_"��DA���� �D̮l�M	��	��=#���ss*�a��rI����P�cF�\���r���.MN���b�f�r���;��\A�����е�vR�R?�e��sӸ��{q���(���T�/��D���N��Ш�mP+>�㇢4Vhڌ��Y��܂Dj	�[�̣.��'ԩI˼�)�ց�zI�YK�wm�إj�\W�:�El��~z���ި`A���ųX�8�s��`��8���
آX(����#��f�ӓRy��}������E��Z2��z{��8tdJ>�!�7'g�R=wO�ծQĳ".�X8z�A��D�� EZ���Q���^W��(Qo�uZz/����%����$_N~��z���F���qp`@��޵B}�fr�E��3��!�2+V�Y�k��RS٪�T;�k��@�Bʡ�KY�鴡V&Е��J�T�b�� VĩK*=���x^C��|_����6�⮢�a�ߤC^�RiT�r�s��T��Z:�~�ֱ���Q����?�x,�iS���\�^Xy��Ͻ���]��(U���m���It�pp��Iܰo?N;���i��cth\��4��i��m�vL�>��uC ��ќ�̓�"s�x����x���+>��M�{���5%����/`�=�q�@H��}���fu���F�cd�Kk$�snk��hV9�>b��}��kM�弮�?r�n�b�K��$Jn[q4s�,[Ӽ�L�֒[�� UWږ�K���Ͼ���؏���1~�.yoO�|�N�c�GG���._U���e�R�t����{
�^��<b�C.n�	��:�_~�k����(��k��^1\	<+p~���\�Ɣ��f%���ub�и]���cx��9ޑ�����b|i�o<�_�׾�jճ�q��ކ�����zԴ��?�će��}��M��%(ʽ������č{�ǧ>�1l����z����*�Z���}��i [3����O[�N�kO�ÔrO_�D�Ø������T�]�Q%15�p���YD�=����3�S6j�x��U�k�F�Fց����V5S�Z��c���M����Z�2j�1˚����p�����,������{D6o� ��|�.����3\����@��-i��8U�X�Way	Mݓ1�bG�%N�k�R�l���h�80*�Kl�s��:62\ھm�6�U36��t���5����a�����l���P�h_غuk�/e^����_?����gK�W��SjTn�K���/�Q�jb��/�I�5�ݻwk�ri���5��fг��*k��^?����('��C�my.E��jM�w�L�I��Y"���Q��ը�)��fõ���I�g��k`�ޜ��ӄ����t�q���C�ZӈߴY���L���9�%�47y�ׄ[��uϰ᱗�Ŵ��&ޛG�^���~o���ز�fLʆZG�Y�����m��eC$��t-=x����L�G�m��bnq_��1u��r���8[ �g���_����/���;%
s1#F�.b��8Zv*�����b�8<u�ۯ�v_�U�Mhֈ
?�g�{Y�{˵�t���\Dcz�:�i���h6���$p��cx��¿�����|	n���ۏ��}��/-�#Q�l���m�p^"�f'@��������������^B�� voK����~�S�8M/)��7X��Ľ����?�qt��x��0yV��OV�ߵp�C6����n��V�|�����i,�\�Ct��M\�TZ	e4C�#�Ӷ֥�-Ō�`@��5�(M��z��mXg������F��}��n��'�CB�3�ů��z�r�mʕ�m�31zZ��sI�;��T5Q�K�d%0Q�/W�o�����H��V�=����h�m�I�+g��B�Gk�ԝg��k��4����z>��D����FƋ%l��fl�7���ǎ9�/����Z����;�](xHf�\+��Ɍ�znЕ >Cˍ��PD��8�F	�s���z#�\�0��ˋ�JgڝJa��� ���~%fI�Sj�I�ʔ�(���T��n2B�˦<���/~�!\��:5(9j���H�P�Hv��N��_�Ci�&�Ĩ�a$43����3���}�b�����flT��1h�O44s�����f��6ۺ��'Ѥ�K:��͓X^Z�Eqtb��f)(��sK�u���?{��O&�ba�����i���$��l1L�@S� O@2�˥2~�9�lCB��K3ګm�cT�@eqN{�@]�D��N����x��|�����e��m��*���ga�y5Ϯ��ИzNu9��04O���d�(���VW��|�'��eK�T:���~�ٹS�~�)�	c��ޝ۔����|ᡯቃǕ�}?�:�����r�����>���S5-k�ul��S'�N!6On�����/�`Źy��q�r��JM�wRA��'�i8��ښ�1L�0t�XC��!��;98�2�N�7"���7ʲF
�ʈ���������k:mW��h:��r��R	IY�V�Q�ć�Y������
; h�e�]�p������1��%+��O�q��D�ϋ�I���X�1�����<r�]c�"����y.6�U36��|�۷�o%o�a;����RL�,q�l�L7�������zЖ��⻮�V�Ԭ�:yzUv�\��pɮ�{033��t1e-�at|Lk�*)7��玧�$5�D��O���3�4�S�$J8<ZA�v,��7[%���c��2��J4Lt��\-�2d!L�k���T;��5�k��F$!��P�����"��g^>��l�#.��5,Ht^�����f��ĵ��M�0$ZZ��|�'$"s��z�;�����e���&����!}�ŗ003�PR"�^T��6��-p�r|b�ЌA����aǕu���/v2Le�ti\�b�T1��dҔ���>��B�P��+~[����m� ������|qFU����s��O��:m�i����ѐ����Q+�pe��&p�B��o�t~<��J����8�k�8�bt�>��������`nf���(WJx���p�|�ZIB�q=�G�|;���K+˲�X��;x����j�Ǽ.�����mq���-^�>3ם�d�#.bv��z�8��hXg�-�͈�i8?��Yg����hR�j��t=S�A]�Ix�g�\�!��׊�N�:.ס!/�*P��g���mQk�
�dɌw�.O_P�>6>�NZGKX-�M�z������W_U �}Z>��x�)S�=#�*��x�w���~��~���m[~,��_%YqtHfy�8u�"
�i0
?w�<�H0���Dݽ��2�L&42R��kvv{��E����'O��@�Vb����2)u�D�.�]6_���U�2Kf�,�2� !�Ó�9�LN�6�F��.#�z�RC#�TZʵo˄��^��ei
��xN�9۷�
U��D-�j��3�ϝER�[m�ζ~�q��D5I������pef�X�r��fc�(y~݆�Ju��q]1@K�ٕ:biU������3�pz��U�w�`����w(����5DB*��!k�#�S4;��=q�;�8t�0C��NM�5��GENQ�2�m3&�'�)(�!#��=�)�1�)]R�B���>3��|^�N����b�Ӕ)�i�3�A��q~湗���o��䨯�J�k�{�6�cm���Ң�=N��8�2�PV�\��F[�mÖ� �z>t�4.]^�'�Q��5b���lUe��p�z��df��!������j�ݐ'�t�a��ו�>B7߳��tyL�{-�)��M�I��_�7{i�<����$�T^��o�G,eZ��*�N�YWyYf_x�Ƞw��ezS�B'�k�����g�9�����'Nh�3N�[�*6oݎ;wa�a(C^�/N�����6�U16�U2:��:]�璱�ckm�Z:��3�͋�?���d3�iVe㤱�زǏWիqy��Ƞnz��f
�F�����lH$���[�t%��a	��a�R�-�(eH�ΨV�[�*����3=�қջً�T�mT���.�K3���Ԁ�K1�j[�䑮n�1݈c$�!�;[�B#�P�;"�;]���<ڲ��;���ֱd��[�,WL�U)o;ګ,f�LF| ��n��1- ;؇x&��m[1wqZl�8!r�	��-��䄚U�z1�@=Yæ����&�-�|O��q%"K��7�FQ���]M',G�����P#J�M�4�lyjT��`j9&��S��NP\��'�~&a#%ש��O�,Ѫ��&�&ӎҠ��̵|�؊��m�.�uG#_�9�����D�w��e��餉��.]DQDք��V�X	����WΧ�׎��O<��ǎ�5�\ك=>�I���d�&�b��������K�����]T��c�)%�ן5k2�E�Ca�uu[u>3X
�RO�C�c�P�zt�|C՚y�r!��ق)5Y �����@!�N˰66;L��uΘ
O������uS
c�?�J��J�;��ֽ����Y�k�֨�KH�.�%/��Ѿ�qt�� s�23[4�t�q`I8����anv��y�1U**r���2��~����+K�a��*��Gaٻ��Ky�|i�e�M!+�S��\ƅ��sL*J�oclbL�W��m3��{t���}�4]�����5;v(؆��V��с֛�z�Q:��h]O�ώe�P���c�=�,=��翽��}f{��bw���@ $$��Z�,Z%[��(v�I���Ȏ�8�lɎǔUB��XE�� �ށ���>�ϝ�{�����ݻX�#[)r5?ΜY�̽����>oy��;Z���0EN��Y��'��&I�1����&�ֱ SU6��D��ᖎi�i(�R�EbcGdDK�r6��E8<ڠW��?���p���p�=�뺠�Xea����h
��/� ���!�k�V���3ʲTt��6>��ˮ��0�i������mP5�R�0bj=ˌC���
�0y�I�K`@RZ�8�ר���.Ъ�⸴��Rc(y-� ��E��/f��K��P����EE@�0$�Mpe'<g֣�$n?z��b���0(r�|!���ك�~e9?t�]��`c�y�q����_x�'�ŉ��a�-Mjf�s��/"O������`�geigΜU�ӞD�PP��^u!��vڂ*F�FQ73�g������I�ז���*-�m=��d����X1.������c���u�=�*��A��&I^��vlۦ������p�N.�i����GK .��~2]fJ�T#a��t���J�����������Je,/,�=��yO_�1H��;�{}y]�݂0y����P���5���l�����n�/ ������p@�Ed߾[����ޤ+����^(09lv�h���g��.�}AM��s�=:̺�#�<��P6+����b�z S��>99��[&�k�.�cw߃3�"��\����Q226�9ʔ-�u��h^��l�e�Ψ�Epv�r�s�6��Vvi�:qvG<�l�l�aDg�9�Lkʆ��ز��i9�VS�SZG
�5���u=yn�5�6�Y6��FQD;�0P��N���z)�!.��/��{��ˢ�׸�E
L�߭ݍ�,��|�� �� ��
߾s�0�bW��/S������Ѿ��Eu��_�e��^g�PT^��f�X���4v�v��S�}��/����ՙ���
�:-<69��]���.�,��'`�-���)�?�iH+<D��Q�����]qa�qe����4�9��19��$JE�a7��q�����k��	�#q�x"c�h�N��at�=�V�
ƶC`j��ǌ3h=�3�g�di��$�i��Φ���ѩ!�l)�w��
�d��J���O�?'��� (���km�D=�����,.�[�7�R� ��\�i��.|gsL����մN�PX��N�_Η�5	�j�Pjeq�|�K�(]O"�������z��U����1/_#��PE�����i���a<&���ӕ��v�l?���g?��M����D�v��9��Pt[�:!5�ٴFVQ.S`��`2)����!x��3ҿ����	�$�s�U]�d#ؿ��;��i�IYJ_ ��s-\�Gj�l��я�t�mz�:�꘮�<
��`r���/o�[�ho{�}oV8m2g7��]7��uԼ�\lN�_���ջ�Z�d���G�,w@�������ew��̸t�yN5�iB�`��G��XAC��@/b��j>�,A
e�zͶ��c�@�f��<��I	����y�-�m�ٞ���u�-._��4�+׎S�����s�f�X���C[0#�by���%48�H���O�ָm1�"������ ;Ӽ�(��8yeo_�V ��c(	H|������?́t4��j�(�OΕwK�|4��C�;ϡ(@h���!��A��Y\�p	A���&Jg�Ġ
{բޛ�8eP#�G�������݅�t&c�k�-Ҵn�{���Z-�عM���s��ʇ~e��7oƶm�0;;�K�.)��7䜌���,��Դ���9 �W*u;rD�����eOˊjF4]��2
���\7� ]�@�}s	H�x�w]>�P��'ޥ"H��b�ϯ�
}��>fk�z�^��nu�BI��3������0�v�V�^���~^��������դ|�6�[b��?{s�+�7a�<$��mOC@�&�T6,e$��i��E��Ȣb������w����*��٣��sػ{����G?��\�(��oh0r��mȖJ:�\�Œ��g撩
���(S4�hV���[��̹�;�R������2��uC0F+��qk����5.��Q/�]�}��<�eɾ�Ju��;ae�Q��<��m�P���b��p��J��iiֵ,B�Qr/�߶w�~h_$" U3nZ|?6�K��h�T���Mu�2(�,E�1�l��� L՘R��&<���3Ks踇:��f MY���]�/Mm<4�O��oΣ7`�"7h�#�)�P��������@�7yO�G���?���f]�'��o	pCU��.��#V��gQ�4P+0;A`�>ćzQwE�XטUo��+��|���֢̼T�z5%8ܱk'v�٦^����H�S��&�~�0g��BG��˛\�H4�ze]����?�%��������o�z��G���Ξ�o��o3�7v��g��[o��_���Z�ܢ<W1�vu�s������_ųϿ�j��zK�������ĺԾ���|��bq������{q��)d٠)�i>�U��HģC��^���9���\����\r?k0��5tK �'�*̟ͥ��-T�(�ߡ�
�.�`c�e�J@�����I�j���N��0�f�R��JG�J��vuS�.�'��g�.x%z�J�ύ� �^�p���Y����s�=�*7���M�����tat���e)���2p52@�ju@�#�ɲ�Q���"1�,�*g�����U0�r�Ʊ�
�v�L?2ɩ恛�qc�Ay�q����A����@��c�R�\X�b���zE}z�mW[MS�ow�k��TE-_B�G���ƛ�,��ĝv
��L9b6/�Y�u�bN�̴\`�5@Ѯ�w�\��S$�S����E&�����������>a���uG���Hh�"웩�F����sy���[EYZ�kW�h�˶\�>^1�@�n�]/�_�*'\��Ы�Ee@6�)�K��˹�%�;���gT[�
�� @_iY�hn��.\��%J���'���l�l7��9l���7g�Y
�ѡ�t@�=I�Q{�l�i2�Vj(����;��Ǐ#,@�ܳ�k78��͟�6mFL�}��~LO^W�=D��A�ܽ{�>G*�*��=��e�fa��>9�7�>��rZ����G}��/]3@� H3g,�|�q�/
:V�4}�{@����Q�����vr�Z7\�Z��ι�0���h0*�܃��[�az,J�2\�Y8� ����,7ȇ�rO�܁R�����W��ug�7 ���^���笠����T�*(������i�&#h!k�=�]j��Ѓ�/��R��g��ҲJP�,-ꂶe�>5aW��N,�����I�W��r����5�����w�0����teܯ�6η4S��_�*ok���>�O˹��5�|�:��[غc+��?����w0�M������"r�(P�Ym�t��<�6�:�d��h������"�j�yg���X��ff�b,hwH���� �M�s��f�v����뢩Q�� Y��:?񑏪�����&J	�0M�1$[��C@>���.'��H��/P% aS��T�Mk�LO7�	�r湮�| ��hF#	@��OXsU~T����Y�~-�m�Ȝ���鄅7 A_M�����Y8�����s�.�)���1�G��z�z040(}� �m��P�Ҹ�pړ05a�L��&q���/Eh$܈'�8&��� r�n?�/|�j��q0z�3���!�7K&�|��ѕ0�k��+������zM���i�}8r�(�>���9�uUV��ʶ�,������K��XT�G��-OɾdR�FzQ��Aԫ͓�L��xZ�6���/��s9OHk��v�}w<�Xw/�&�t�c�s�P@�]��?%�_k���fB9gc����ug�7 ���Bghl�]m���&b4:�Ŗ�E_�Jj�lk��,�>x��S�zЬ;R��]�<� ^z�,,,���̝۫M;.W٨�	�aڐ��v��2�uC�ͦc[�uN��pUOh��e���Gf&X_��1���͈�[�d!w��hWS�c�Q����	7S�v]�1��Z~��>�=�6ֲ����Jnn�oȗ��B����<�ilS�X;f�D-0�)q.�&�t>W���m���+S֎0-Հ	rn�'�nK�YKG�Xu�}�mft����rA��?v|��#�Mp��o�b4��vmFB�d�ZQ�.j��,.��Sy�b+����ԙr�(;��f۾ӣҽ��x]5%͑.�G��PJͺyY�=eK�-3�.}r4�q�z��2�{z�m������z7<ԭ�q3�H `�M@��קY$�����u���:A��𙲌f0:[�o�ݢ�˕<z{��PV	`���S�&-|&�eyFb	y�(
��TK:����ܽ<?���
ye�uF�����_^e`X�f \k
`
�����}���^�/�D.�VS�sx���P�`�Zi�!�c��p=�K__gm�n�a�,o����U[^O4$�.�(,�e{pe!��o>�����l%�;����H�#U�O������C�m �-�	[Ԟq�m��e�Z�d�rA�\.%l���D�X�[����{�:���9C�yb�<��	s���;�3���߁��]Fk�Y,�K�M�E�h��7錻e}sn��u��#��2A�&J9c\�+H���Q� .�h��]�&"��,M��-�!���7إ�0JE��~,�N˱WM��A)d�`"��=��1�YH�03���,���<�}�B"E�X��­���wN�P�#�+�b�G��mT�"��ܱ��j�][�46�<$ ������$���9����e��H���n����&�&|�Ļ:bg��T�Z_��#�i�S�.��j���7�Ȗ-H�q�f��1�n떥Z�C�v`)W�����˩�'jHMW,	ܶ�3�bf�ĸlh����zJ�r:�����'A����b���;���!76���xÉv
�",4���*��<0��q+P����JXMz��jyGK?¬k-�fu�R`����a�����4#�6�H�耗_zU�	�$򣊛ɂx�:_�x���{��'�qVJE�VV133�h,���5y.���.����8~䰎�]�2��95���%��k)J}������.t�nXj���Ϊ �믿k�,�} |��9� �沂���.����1#�Z^�Rg������hI�Ph��<208Z�����r���@��6���t��n�^K�Il�b��Ҽ���|1��������)�ʮ�#G��ɓ'd9|�=�cnn>�m�����W�E�q�.�s�
����y�M��!˰�����\kǂ�|W�ꛓ}�hO�R�ő3�lN�d1�oea���P,���cB<I�%˶ �ԥ����ܡuqvt�k��^;���UD=�s?��w1�*M�|j!�?~۶lW/�|����	e��gq�ʌ @ݤ������t9d�ڿ@����Zkf����[��# SN(U��W��S�^����D�t�uP�^�N�
����D��:��_�Ϲ��m���Q+呈�����N�	H��D�2�J���P �,�S�a��X��������67ђ��`��h��R@�����ӭ����mNb\�L���,��4֦�a�`ei3�����Eˀ?�)n����U\�`r`p��4�F7	;NkS��I}]۫�����cu�;6:v�F-�ִ;���V'N��ϳ4[r��U��`�E���>��u9�����Ё��f�_|�E��3��f���ƸمE|�[�BO?fV�z;��2��A���j��:&ђ5����~�x�m�6�� ����Q:�g�4��zߔ�s�4֖��}�a<+ϣ�="A��|�X�jZV���T���~ط@��6˱Z����mF����� �/$�P�FCl��� p���
�+$z������b�o��XFZ��P����۞ �Ֆ,>.�2EMr��>΍��7��AD�qaZMe�����x�u�T+�D7��v���edػ�Qt	=z�0��}�똼x~���G� ��^V*@��.xowD��Y?/-$A��x^,_xW�Ə�~�S(N����������ȯ- �c+�ڇW�xK�cYNeM��2J���o9w�]�uo�H7j�sd��L#7ZU�j4�(a�^a�I��K�dX�_�$�ib9���5J�ɬL!�wP�s�S;s��y�^������������:�Ȍ@�^��\_\�:���8/AA��^D����H[�	n�4�UNgt���8v��k���f4��ӌ�mR�.# d�������Q9f9�/��˫\�����.�R-Q͍���*�GE�ӊCFz�.~�9�~c� ��g�6R�ڽ71ܠ��:����*�d	+�)$��:3N����s���c?�{�:���O+S���q��e�&L�w����#ﱈ�ק4m����B�|�_����Ў����vvڦ�:u�D֞�@;.����Lyt.�e>�nf��� u�����e2�i���eK�Ww˵�j�H�\�g����n�m�o���({Zv�EyI��Z�,����3������(�g�L76�\�g�O�,��������́2�l��ld �dR���)��Ζ����%J/�Qe�EyS�7�=��֩��~�,���w�5hh��q��{vcp�GL��Ue�[7�b�;!�Y&%Ew,�x0 ����D5���0d��<�v� ��(�^�������� P[����1� ̹��DG��W��.H�@u.6h9��fg�S����H�E��yLwzK��'��,ks�ђ��}S�*¢/�>)縀��8�Ϝx/��0Gj{7tF{%�W<��~�zޙ��5��^�'0W�`Ivh&�Pr昱�P��f&�T�\�������9cb1�ti����X���4��1�W�����*��R-��_�nD�#Ȕ��pr�m�['��TJem-�}ѨH�蝪BM��4�S7S �v����iSl�9�9�W�Rrn�����Z/�PL	p���
�����S뿑`(-�ը6���}#G�A��!������\��J�o�G?�qΩ_��S��.�:2i�ҍ����/�u��l�������Nr�odJ`uZ�������o��",�����ʏn���P��
�0x��L!����6 ��M[H�,.�a�<$�ܱ��N�^����<���ʱ�y�/�}�Ҕ�dM-�*��64A�s�QI��1	&�PT�
�ж�V��8���<&ʤ`���߻ݝ4�c������C����׶�R��HЍ�ΨqI!�EhUXi�B7����E�G�V���сX$
MQ��~~�[U���[C��z���tX��(�b���<u]�� w}l�'�TQf���r���lZk�����.��d��Li꠶����;��߼���d���^I-�㢱M�CB�8���j��'p�]w������[oⳟ��
���l��'�P�1��,--�ܹs�M&�F"�����k	`faQ��}�_�rY;əf�<Z�ƌ�n�{)tL���o]Piۖ����ɳ�Ne8��3Wߴ�Ѭ�$� %͖s���]��8��=V��N�!���n�I��9̯瑓��ްu�m�
�0cМ�|�o��+h��>�c�8z�q�!��[XO}eA�����'6o��3y��-b�ZI�<ׯObumU����m�}�ԑ+T�?8�G��6�mځW_?�l����o�n����������n��ݿޭ�7��;`�N��j������Sq��Ӎ-k��wT�W�\�ܾAll�ζ���X�����W�;��uɁ�{�q4��GSz���\Y�:^�c� ���ԯ.��oK�9�2�,>��tG�6� LAa?TʢJ�����L�ݴ��D4̘�b�Rbw�k��
��	 �}��!���J!�z����O�R�_�rM���I�||�&�۪"
®Wڣc�ʻ��K5rb���RkTn�L��͎��z]}]*�I��/�8���uHn�,��W�r.�u
 (�� zT��q�i&���߃�ǫuPzTޟҞ�^l0#`���l���2���
n�}����?�.���um�Ri{ʿ
����{��4������<�ǵ�2B��&�r����>�-87 ����[v��*#���2�l�Ƕ�	-��V����6�F��j�_~�i�G}��<��¨�U	t\P�-��(��E����#_� )@ֿ��\#�ek��(Uy�N�a2��q�F�N	�ۖ-C��ߨ�xQZ^CT��T�$x���*`_��է���@�h�&AE]�!l m:^e�=}�K�;fT_�U��ݧ!�[�l����kHd��O�����f<f����?�bC���)��}��NP��tp,(s:������L��乗ϯ��P<ck߳��?����f;u�mr�&��Q�m�"�Ma$�|���S��d�^C�۸�y������D��bk��-�!���>5����/&�T	JMߺ����^U�L��9���m�c׺�;
�ܐnՙm���S?,����G��(r������%�`H������	A�b��.C�h
��<^��&!���V�����H�@@Ev��\�VW�?�����hj�����5������@'Z��9�ձ�@�����.6`��4ɚ��l�#+Ksgw|]X#�Q郭�$�&�������:#=�x_����;�K��c���<F�c��q�b�q���A��5�2�#͆>��hz���Q�S�X��>�k��U���~���s���e�m�1��{��t�x����w�A�2�gΓ���-�Y��D �g��M�Md�����N)��r�}��W�[����x��2(���r#r�黲�����d�	n�Ǒ�t.��Rjy	��%�1\�6�(5�9�2ʥz	]�s��3+��z��c�>����V�g�f��ξu�yU���R�&��8�c���rT�.X{L\��)W���r�>�(�cyU��f/ڤ�ϣY��ݲ[�ƿ��[U�n��������iY��qy����aOCܣ�V\�ZŊap���Jepu��̛ͲV�k���!9�F�P'4v�
Hx}^]pj��vpKv�UǽZ���
#��l��cT�+� �ܚ�}X�iS�hϧ��]��9�����ڤ�.P[&6ax��ΝQ�o�6�'}Z�dZ�����}�e	&�g�Vw)�W-*��ሀuY��z� e�[��`8*�9 @^����|nH밂�]	��I6$8�s<�Į t]�<93oyv�K��}�Q��m��5UN�m%�Μ9�����L�����}�]��3O��������g��櫯��� VW+ꞗ/�j{c�Qr֡��x\>��Ա�^� v��*{+�m�¦��)r^� �\��l�a�V'%�tj"��A�\'S�mЂ�Q��0JR���HR>��
��,��ۣ���ז������{ �x�ӶT�)�QF�i���#��F�Guۂ2�"fc6iyi}�M�h�S9\�x��;�=jQ+�AO2���ӂ�O[�C!��s����xƑ��~�H�G�"b��.��j����� 7,�C�Y��ؘ�����n4佧������2PU{U�lW:������z7��t�c���w�3.����HS��%]"���4��_]}c��k߾g������_aX��	�	;Ua��FA�T��4T9���J`k�3����iZ�/�&�������AKPY� �P�Bj�����|p�~�О��HYZ5U�ɂQ�U4�蓯:A�2�>���*'��M�U��N����[�!�ک����N��u����2�"��),��annF -��T 3s�:3�+��n
��Ͻ,���eq��z�C�������򇱞/#�.b WF-QӲ�zz��F���0m�^ϫ.;B~�������if(h����e9�a��%����?���*�P]k3R��\�K�:��)fq}v���x��4��ƑMq�;��Jcne�f�Q-�� c��� �麒qu�������zKK�j�":���Ԛ�eiK��M�]�l���j)�B;nz���\3-#��&@�����=a�H)Z�.�#�o,P_��
F��^��C5]����J:����ta����+�%�5��{��-���FТ�ܧ	��%�<�$8��w>���8JC8��{7̆br�|����O�:��N���}"'׍�$��}L�#_���Ջ���8��&(;2�Y����9���:�0�Ռ6t���v[���~�Y:`���3[Y��~�~��J�Z�2�ȏ&a�a@� D��QW�ef�q`P�5�SA$�7�rn�]��4���ח1�� �o��&���+�����޽ull?��F���}�+�{Z�fڝ1�B�ءx�ǑZYD@�p(�r����=�Uً�>�&����bDf��0����6�vC���������i}ur
s��x��wPNe̠�ק�i�>���
[L���u������
���&�r1/�kM��Ma��x��K�~PEY��n�uaM���l�FF��d�L�r�z�g����eA��%&��m��Tz�>��eJ9�Xsp����m�?�)�¶�y1a男�xm>��a5�F"�E���4������(V�H 쁋z�,M�L���s8V���u�{�J��jp�`����u��%�wϽj2�}�5d�\,N�� �鬎O1[16��a�3A���BY����
���q�,�@���x����$�
D��e����p�sm�\����	��.
����H���,1�Ӄ�\˨{p�$�
&9��Ҕv�Jzr�c�0�L9vU	�<�<���VA�;��OW����w%	�V��s��k/�+<J�,��HW֋9��y�A(#�~
��2�$�������OA��G��#azq�f�4��_��͛035�%$���\ӂ��O�U��y��<p���醷+��;��ą'�u��~�q���F��������g�=���e����Ł������@����۫��,��̤�8��L;-�j,�亮������WД��|N�?���m�.��]�����j���T����<�N���lC�`6��m�o���p|mk3��*2>:��^Բ+Ȥ�dq_׺m@Ť g�	+�wl-4d�f�w<��P_B/��KǨ���0?w�c�a��_��)�����0�
L���;Ǹj`���p_���=�Nm)dJ1#,�R�Y�z���X��T�Z6��h$���^�kVf{1:1���%Ν��	�IȂ+���Ay�f��j-zTA�hZ0+LO��4Q�^���c�&$z�0	X��ؽw�p�o1v�l0k,eUhf˶��v}	��]��m#���$�h�<�[�Y/� e]�_�i{��*1�M�����5eZS����K��{;7����~�n���I�-,����t��_�����җ�����t�inzN�=&�AP�#K�Wa�k���%��+��lA	D�WR�>?�V�q��yԚ�d��؇��*�K>�֯��I�~��7�n�y۾w�y}]Im�zm
�}�U��p��d3K���߻���HČ��{������g�r��0�Ƨ?�)#�IV��p��{x����|�l�����|��������{�+f
�na���ؔ���I����$z�&}�;G8�����Da	���ق|)���>D�1^Z]Y��V�"^�b�)�f�$����2��@]��u܏2Ȏ�q\�����j��y�1��^(y�N����̰as5�FA�<2Xa�GF�����e	���^�H`Pa(�
�k��Y߷��XW��BAH'2��{�\3�q��̮���@��wl�_@�h���n�,r{;s���g�p��P-dPv�tܦA�Z+3+4hД�������>N����vk�����U����.�֒��d�`�5/24������YMX<�w����7���fˤ���Y�tf]�L�~�%a�-A>�%���
���Ք�ay����Wҫ���t�����.���b�I-*K'��ZK�u鹈�=�e��j]ޯ����6�o ��ʪ72#�6_,���ZE΁�!�{��-�>���Z��L�Ak��8�m�>���זg�v�c�2�ť
������w%p��UM=���~MMgrE�"	��ߧ��D���O
@�y�bˋ+(
K&��>.�4(�Td߆���K����,�l��k�DO"�#0��u'��؂R�%L8�L���}���	"j�q����:"�#��,k�A (K<W������Gq��^$�Q�n۹I� ���.2�	����=���}�fn�ي����_��z�e��y�؃���] �����V����}$���s/���mDcA�w�=
�B��3f���2s:��-Sg'[�X\V����b���z9'˩u��[�i`znR��A,���,0@�����;�XJ��t�ӦӜ&�G�$�2��69��P#��C{|�z���`Y̭�3%	L��uͤ�%c�u�^^���mJ3~?���V��zU~�^�Lx���>���h��gJ�U�b8���E}O[�q�;ѐ{8W�m:sa򡧮:_��6����z����O�f��؜�M�;��˦�6G�ZBX��4�I��|���4��x �WfV�dtZf���鸕�ш���;���,��rI?�Q7��d�>���
rC��v��8S�4��Z� A�e���M� 0��)l��{�����D114�ɩ2z}x��{�n�<d_�C���(�@"aT�Vf	��<�ȫ�%Y]��^���7,�,�Ӓ�;�R�*�х�d����s*�q��W^�����l�$Q犭�]�;��yl&d�Ӹn	nRª� *Z�P��R.�
�$�سyBίa���#T�0d-�צ�|!-����
�28{κ-�J���G�]-�W^�����w��.&''�{�v,	(n� 1:��ͥ�u�߿wނ�Z�LO��Ia��0~��?�/|�(V\8���+]��%��ԇ�\�J	X�\���U<p�><x�.����r��2�#�1��c���o�.��؅G��0e���.f�y�kk��g~���5��#�\9��\R�ʭ�1�7���s���˓�z���!���?!���>,�;y�m	���g���ӝL�u9���� �X���%t�~fP.�C��b�k�j@��8x�W�ʑ�X&ggp��e<(ׂ���w�Ӟ��RojI�}v˥������s�y}Wg������/p�K�kK�<Vv%�r.}(�+Z�XK�i���P�g%�
�q�>���s�cg@�.�v���|�cٗ�
������
�g�-*@�ɗ԰��	����������?A�/��6�៷����7.蟵5�vȱ-���0�|�'�F�YvԆ3�NauiZ������>S��� �ɤM}�-��/2p�L�9��i�3F]�T("(��xM:�y�:�D���$�7Ч�`L{6�1/�%��6�@���& ߤ�
�j�J�Ғ�
�W��Rה>ߖW���a�1���s��?s��}I��vo&;��s/ˢ[U���0&����+3���@���߾��%6�Y+��>/̇�[5�4�%p����<3����u��q�G7V�\F���x3 �<6S�,+��zZ�=3��陚\�U�䵬�SF4(�G�N�5���J����Y��~O;���� �8(����ɂ���a~aYg�kM�N���ϸp��8q^;�)�%h	��إ*~l��E�8rh�9
�{�eM�?|߽�ilPƩ+����|��̓���|R�n	�Jx�駱4=���ߡnp+)<����ȇ�w,�mۆ��@�0Fz���'��)���K���yc��y�w�m`���SOj����}߄?���sZO���X�Z���ȑ}x��a,/�����u��7��{0}mg�.cb�W%Xhͦ��-�u��l"�I����O|3S3*[\�kO�c����|��L����y��#`%q�ꜹ[FpȾYYO�S3�љ���x��v�?f���AnJP�d?��|���(`E������=Z�����&!�'��� <��F�V�n,�Lc���:��V�?�W5+���T����R*�v�o_������k�pW�{�^��W������~H}��Y[�Y8�i�1�:G�ט���&�}Q"����ម؄H�WG�:��K+:oEu��;ޥ�ӻnY�� ���'@���4��X�Q�T"��L:;�H��z"�-=�-g���ʲ8zn4��?�Yn`evua�SK�p��ii��L@I�]�w���'�c���(+���GfeI���G�Ӻ�-��y,.�(��J�A����]{�x�������gQi�Ǆ��
&�W���?)^'N����m�49�٥U�J�k��)H2�0��.�L��t�)H�PS����ٹ%|��Ш��;���x��`f-U�,����$hbw��K��e�f��
kcP���'���^G"�0L
���=�㏞�.��w>���U,��U�,W���3X��" �B��;u+�i�_��W�g��́^A�+���+���w�[�+�Y	��_D8��ض>8ח0�F�;�s�
ұx �=qw��8wv�� ������Ŀ����j!,���:���똓�� c(ѥ�����^�V���<wD'4�Z�|�������w1>�,����Q��i�Qw������s\��^;q
���dW>��.�~�0�Ķ����Z50�i3r�rr.�$�j4��ϙs�O��!ٓT���%	V9��T�_�c&:>T�n+�����ؑ%ϐ��I��Ԃ��jo��.^��L9���D{���2�E��륚�W��3+�JP咩}ot��Ob���E��ڗ�Z�o�sN��P�׽Z�y����k��}[W�/��W��t%Bs�xo:�C+��yD4��[�����l�,1���E��c����7�?kkԛ3l,[m����0�J.� �߿ހKm%�ሰ�M������7����0���>�T���BC�9oҏ�ZF�Mq�.a�ݲ�b�nUn�5+*�e�Y	.��,��e v[`7v-��#,�iC2&!)4Br�ۿ�EM_�_0�~ғ���*�>3�(lxIP2�\:��Q��y�x|N��e[�>���d���5ho�d7��p���'�U�6.�'�_��ыB�N[3�ZtM·~����>S�5K��.����� ����ٳ��*���Fa���27�][�DS��X���nd.�-�r~�T~��b�K��3/����LM]� ��B;�wmÿ��_�K >d���l`inC##�C~ejUa��B8�g"`y%�յue�����|w��������S��-���cǵ��Y�M¼?��O�kO<!���a��'�PP�)��sV/H�8Ѓ��(J���z0<��!�*�KuԿ��󯿎�^y��#��#���{��q��;T;��6�CG�J Z��D�ZAw�c�����12>�y	��6E2�s��e,--S@pޒ�L �V@(�ǫo���M�30���vc!Wӎ�F����e�8u�2�%�Kbtb+<�.�=W�����z�ܫ��W����h}uǾ�}�۽|=OJXev�SP��o�ma�G��#��w�$$�����$$�G>`�֭�|� ��DI�=�����=�J!���=�7�P1��r2�z\�E��/ϭ�����~�w-��.E��y���p(�� Ԯ�b!��zr������}�ll�E��c�{�o��;���_�r���-ۣ��yص~G�	6����q��x�a����b�U@���-;eى�c�n��fr�s�
;��_���3!���J͖�L�G�z106�����ϣu��,r��lr4,���VT�y� ��[S?�*z��x]*��Ӻ�ܢ�M�+)�{7��\�+؏r���AZ���r��7u����,�Yu5���o 9�+�C�c������k���Ք2&FEM6��]�i��n5_�`å���\S0�ik=���!0�V�n	�������UT��m>RKk����	k=�ARE��v�`0z�q^OeA_V�i7-,.�P�����o �ݏ,{u��/�.��JZ��8qŴ��w���鵴6�5|Q4ب�FB9���[w��w�6)�"����_Cf� �B>l�������3(�w�M�ݺA˧}�ǆUB5!�˖ M�
��~�q_[/@p�H�]>��O~�r���^W0"�Żpt�mN��+���O���^}Y5	�ڎX�'�مe9v�{�$�ڵc;��ۍ�_;)��B�Ȁ��W�i5����I��� �,��Y{:�s�����RU�gS�8{u�X�Ra��+s˨��=1\��Do������b�g��LW:�A0��"ϙ+�~UK��9v簑��k+�z�,T�Q��/�ǣ�Fr�����w`hxT�<¾ r����b_����'�����{*��;u z��^e��A��ASS_ei�h]ΉO3ra���T+c��ʘ�� Q����T��K]�3���|�̶��vߋp���F=ujH�8�J�D?
�%���Ԝ#_�	0z�
r`�OU��вۜ�m�����{�vL�,�O��ELf&�cD⣏>�w�=�i캀^lh�dL["�0�.��,�AXWjمm}I���ؑ^�)�߫�j6��e��Ű2;���W�;w0�uTW�K��Y�E)O���/�
�z��Ŵ� �GdA+��hh���ER����p��&$��9q�q/�#�R����IX���F��fkQW���jo��+y�f�$ w�t��
b�D��ed��7�lt0��|&��M[)	t�����	�yV(�À��ڲPn��-���
�](�����s|��
�S����F��N�̒Eߡ�mA��� �Ǆ�S?�|�+��E�Qc��^��r]�j�ww��@�}�F����b8�g��aB��ё1��7��#��D�@B��=�<~i���LZ���~�6S��Q����;H	9t���}�p�g�.��Ó���#�pϡ��J8u���_�Z!���n�ڷ�t|���RNv�^�;�/�}Z�G���H���<���}�m.K&���S'N�����u��B�h��X��\h`I�D����k��8v�"���[�a��\_��po/6���]H��t������^�~u���J���ZHʵ�}V-�V]���έ�h�DH��l�����H��8��M�P��t����9����Z�k��{�x�?BH�/#�o��y����}U�{\]i�H)I6u2X���%h2��֐��y_�fz�KB��14��|�I`c���6 �V�&(�e�d�Gg]W!��NHH��F��˗ā=�üQ:�٤�jH����}.[��&F�I���]GO2�����0:��IG@h��]����O��Y�G~1��L
��1��11�Y�q[mR�F��u@6��l\������a>��1e�&)4"�@yN�s��ʗŜ3M��͚"���މ�.Y���
��6=�����Mt��hq_$�-�Ǆ	��e11R��BUX$uƽ�.e(p*2��2s�n�<kJ������!�tx�T7��N��hQ�f��١�
x�q��
cd��?~7a��(P���|+�+�x�2�r}�!�����ޅ-��H��ڈ����w�V�y��-�%0*sop?Qr֘Uk�c{�Θz޽Y�}d���ً�0�u�z�#.�.@yt9{�!<��k�%.�v�nW ���^,�e��_�>���[~����-�� p������=a]x�7p��4�����:t		�����r���� ����1��������c>=���J�9�k���`��J���3s3�u+v܏�����n��7�hO� ���;�nif�SW$X�����p��%a�~�s�q��痲���5	���A^����؎_��'�{S����:����+�jQ/E��D�s�� A�:�F}x��U��?���������D����=�y]r��E��u����Н�H�"A�ϭ=���ٴ�{<�H�rP���4�7=>�jE0�w�^�x�-M˳g�*׍EV�G�
f (�S�yP��j�U*�ַt�c��h��x[��]*4�)� ��@m�~m�ey�]�l�9\5o`C���5aKڭޕԿe-����$�ض�Z���6K�7�m���`��N���:��ed}��!94�O���qfn���U��aǎ�������
�KIn�h��$�ިߨ��n�o���Gq��e��q�XTe�������Pj�D����jdMG����8�s��c��QM-s��i_�����+�cvy	{����>�!��#ά� ���,N_��o>�<�|u�jYc��8��Qf����KA��2).v�aD�qa0&���^�@x=zNu�����d���K�}d�����"���z��|:������G�}5	���a���Q=.�z������GY�$���%�Q�1OP��(���P�v��;�M��K��['N������>5���hH��y�nܶ�6���o1;=����(�f�s�7�mG���s��8`D����W	Vw0��S3ڶ����,Mӗ�vy���n�Zq97�>�c��G���3�Ƿ�:R�4�wn��w��*!;�XP�B�� ��:��S�۷"�0C�Q��=[��G�b�s'q���%�bI�]`~����ӗ��Lǎ�&��q�!ݶg�Vt�; ���÷KPڭM�����$�)op,w)d���W>��b]P}b�6��N�8sI�I@�;}=h��jјF�c͏�]�ՅY��]��܈�c����)�� xwo�J��=Yc`G�>4J��͛��T��6^���"���AZ��Y0�`�U�9}���g������i�꟮/�ѐg�'ܶӰm6����Owm �-���+n��k�,��NW�P�9��vKU*�6���Y�����xYK��J%KS�S�ϟw�$��)
��+a<��z����IT]FZ5���ŗ^�:���!M�Ry�C�W
�t�R�)a�5Y��=]XJg�\����Jc�M�lr7T��n��������P������=���ɿ���b�Պ
�D"|�cGQZ��%<tｘ�G�W���ܴ��czua��z�e���aj��>�TU���X/��p#�3R��(�Ԫm�3kk(�ߐE�mH��/�5�sL} :��,lݵ��G}��tB��t�'ƽ��&1%�����#�v1��M�@C�q?viY�/,�
�45��YyM>����S�e�~�*]Ȗs8�9������ʂ��Tj٦���+��{-$F����ާ��CC�G~=]F��ܥ��K ��G��ɉW_~]���Zx���p���7	c��o����I9/K�Kؾe�N$0�[��t����������*rr�6m��q��^�����C�%���ƓOW����>5<t �>.ʭ�W&����^<�����!��X��7߻�-Ą�B�j"q�{�H �&ļ u\}�}��BB�F	�ΛG���@��:���K�D�-A2�\	:��i��� %�k���w^xEG,�r����~�#�QN��#A53A��mȽ��s\�g�� ���M�G�mlU-74`dOG(���V���[�5���D2�}���s��%.�>GP�-�1hulӍ�^��yf�<���)�w��	�r�v���K9�mw�e����m �-��|�@�qE���_}���-	QnTU��>�['�U�% ��ŀ:SxL��T���|}$d\ǒ]=�qM��W�YP�i�2�F���LA�������o`bd�bZ��8�Sk��9��߼��uP&��B���0�"�;�����P��Q��&G��TfSk�ڭ�	Mޏ�=�#�x��� �'|XY��k_�*�]���1|����p��$��2�;w���Sϼ���I�z����k|b��k(Q
W� �'�8^(�ѭ&�0�H8�Dw����0`�� ���.-@��^eh\+k͚	�p�}a9&��S���sϠ&�ç>�)���184��T>��5��g_ĥ���E����a���¤��l]Bar5��~	*��y�:s�˕��ë ������F����G iTF;{�
�NO���,v.�`|t Gn߄=��%x��=��)�ӧp���=�������k�B��,޺0���2����ož=�8x�N�(m�s�B5/�"�ӻ����ݟѬIa2��]�ߋa�'۵k�yR�#�@YNԅ�9	�丢]���Z*���s�{�^
*�{��v��źU7ݖ���OJ�>��v��O��r)"Q?�n����<N�VE �B�~��~wLa�)[1�t�x������N-�.�ɏ>� ���vџ�2�o<�,��k�
�rxQ���c �f2EN��=�A{�Z��u	t��;�<�S*�uBν�Z�i�R7v��q�T�n*4r���J���ء̓j�C �̝�;�U�@gvK��nG�z�7M��KZ�λ�;����>`5�k֪0��m�~�l�f�#Xbm�r�Q(�k�b��2h�r�䁦�����==�-Y,�V椕;��թ���U��/^��.כ�x:H��K]�<���qu{
�wN���
P�e����R���(ZeY|�ݷr�-c�d��!N��;��-
��r,��Q76�F�&���u?�i��5��p�,��*�t����2V�����>��n���\�Y�/?�]Ȧ�^��^T�R)����nR�&k�-Z��s�S�B�ˊ�ӣ.g^Y��o�[��Q��:���a�4�I���f��[��ei���R�B��K����('�ZI���vw�ח���۲`ב�]BHw֨����H��h�*���O5��ܟ��R��7�4���x��YmL<~��JYT�=�
�=�ҫ8q�"�6o�~�9|��;��s��sz	�կ����Hgh��7�z?�� 9:�-��'����ex����V�������?-Jo	��To��.��G�k�c�f� �njaMKU���Djk��3]XZ�H�!��*�sQ�{5W(!$[�c�(�ti%��������׃�FF��h�� ���Ԋ`�x���G���'>$�-�nM'7XS��\��U���=�n�B'rI�&�Uu�O��r�J��UsុB,�7���5��0��Wb�\_L�e]����ϩq�7[r�)��6��-��e���t�f�xM��38oH LfNP�3�g]��9��r%��ʣ�(z��o߶+rrD�7�U7�����VP�_��<g�\�������y]�]���~��[���)�5���h��L�̾jJNV�bQX�D��b����Lb|�=ʊ��jq��؝����Q�bw,G���`�������yY 8�6�6ꍢ�O��ZZu8�Nv�0ئ|/
�Q��H.*��
����$�Pٜǈ�Mog��Ɠ� Ǹ������2j��GI�[��?�D, ��-�@�A>7Sh`Rظ#���?��^}}}f�kbP]@��Yj�U��DP�I��ˤ"��
�m{Rk]��M�S�*�Q]@w�~�53���"s�.۰1W���:��)9���ޙ�Xv]�}��Nuk�깛�HJ�j�YEKqb'���%A�΀<�_� b ����0�؀-[��h�(1�85ɞk��<�)�[�6I��ͮ����]]]u��쳿��^���c�eL�)�Dq�~��U��~jz^���}J]����uAv�{���!5�`X��� ���V*y#����*���^��^|U��+*kV[��o�K�_���+C�(��_��Qw7-{�;*4(�R�.H���w��({���;�1o��AS�횊���*j����;�o�rb�&S�k�zV���F
�����cy��e� �w�Ή��mY]ې3˧ekmK���[=��.�gб��������D�ۿ�������6��b�������m���z.�����M��~S�¼��Y�8��ww�M�	��,���kftQ�^�����j$cLRkF�'&�v_B�f�\�Ϟ7�EјR)��3��>��P�G�"��lȜ�{I��KI�j���y�����G�o}���O?)uw�IMѝN�/:ڳ�.�82C��ʄg����Sg%7�S��`s�W�n��E����;ygE+���ī���k�?�;j�f�z{��Bo{�(���9�S�Pݵ���uQ��V���~SJ!���ejZ=�A[.]�(�/��3�.������B�KJ`�E)<K]��=�g$�� g���]�A?r�B�p2�^P�-�d����/�����ݣ�����!'�=�U�Q���C��e���<]���\]�1��R��PҮ.HIhޭ�̋/�`�4���p���S��.H��95��ђ���/���������*#�T՛����|釯�����l�\S����ٖ~f���
|Xqd�����Ң�#�vw�ߎ,U�єP�^��Xh}����"��ܦ���|σg�3?�Ko;w�aQ=�1UO���0?Q�Evji^>�ُ�y\�[M5�.]�l�Xk�=�ǽ^�Q�y�t%N��V�T�׵@���P�o�t�{4��7�ݚvw �V��n}�F��iw$����#W�]W�p(�/�����{�c��u��-�>̬��d�@�Xv�$�Hk�c誦_:��7�R^߳�#l#�s}���6���V�<�Lx��Rނ4½Q/7����ۥ�m���T�U�;{���a��K��y�p�yx��i���G�[�\��MU�b��<iƉ��sL/H�9��Vd����8�Q�7gQ�{س�J-T�F�H��*�O~���<%sU_�*�U=�g�58��&�����o�׿�e�xJ�Mg~�
$A��6���g_��?�S�i�^MVx��a d}mӪʡ�_�Z���Y�x䮋T��C[�x �Z��j]$�4����y��U ��lM�⴯s�bem��A���=7u�4$2TЏ���I���p�*6�֞����ZW��j^&�i7p���P-��b����r�Zt�A���]��%W�^Յ�gﵶ�*����e�%EA]��sj,袮�r�Z����</�kV��S�!��9<^+���`-M`��:�� q-��:șA�3����U}�f�:m� M_�s"O�wv~IzU�p��~���y�Tqq�-党z�%�W��O��y���*a*��>��<p�5�h`�SM,������̌���������yKݷ��M����gr��<y�*㕰=��=ҍ݌X'� �r������?`[����]�ޕ^|N�`hu���u��Z����o��/,�'?�!5jy����u5�*zo���@g�� 7�������H=Dgy<¨�8¶;�y6v��{��'��6r���N��ޞ^�P����7#�;�ۍ�o���Q�o�~�(�̖��X�b��&z0�p̃�(����y�<I�������k�}�,4c$uQ�еR�M���{6��2�:O��5;cn�l���h�g��P��k6�=i)T#Ro\)z�PyP�Ft0������;`���B�j9��	y�k�v��z]}��~���$d0���r�I������c0�u|1w[i5�o}۲L}�]v$q�<�ώ��rUVV6�ƍ��GS���b������'�_��6<O��x��ֆ�=g���X�;v��Qs8�� y��y)v�\?�b��J1'(�a��Bq���=A욏�f8���ԙ��ĥ^�c��8C]X���3��c��š�m
N
*�ۛ�!�UdW��"}�g��TeP��h�q�7�^Z�Vj��B	5[��a�[�Dn;*���E�`�1���夹���/��ۂ����c� �ejL���%ܒ.�%���<TK��ɔ����j��˃��ʻΞ�AcOn�֖�����ݸzE��k_��^Z�s���'M|���n���6�c5e^U���3K]�]�bۖ�n�ԃ���Vħ�baذ}�����2@�]+)[QE�Ul�(G�d۔��P���?[��@��|S.���dy�*������*W�\����\F�GEv���d��I���ep�g%R��֟x�����*�	��K����4o������Z�2��<�!0[�=5�Vȥ������8��UY��-*�4'�7�=���޸��	H,.�E��4�	n�*���	l�r��z6S\�3��M�L5�e���fVq����9	�5ٸ�%��j|t�63/}f窲|rN爨��)���|o��C]��:�����Hk�.Q�K��f(���F��sE��)�m���/^�$'Ο��i׊��Ih�;�>l�ovD^}�\�ړ��}C��s�weX\]�e�K�w� �!wO������-�;�!x㮍m�qht�w��ݙ;�������]�V�U�M���Ǥ�
feL|.C����o��8�07��HH8+��wM��ch�Q��k~�*��Z:��)�?3�;R�x�4ej���d�+I�w���(0�ܯf[�`��>!��S\t����1�߰0��ZhG�"U��#'	��,E?����<8P3>�>W�>�)�i���=�N�AU��"D�/�@�c`b��i6����#�1dx���
aR�߇#J�H��a�C���K�M^���'A&����ʛ�a��V��^FT�6Ue���B.G04ϒLW�Y��u��w�L[qb��uer�j���>A��ۼ�ә�9��a�΋H|����'`E�T!&By����w (zCc�V�F a/X(8��JG��Z}�b�zl#e�i1�Jeȣz#��`\�"���#
�� ���~53����8-3�]$�����y���{Z�v<����f�y�Z=�z/E�1�WF*��Ye-Yf��*3Jsr��S�5�'h��}n�m:M=4���m����F�*���m�?4�s���-�T��t�B��y9�92�j >�����#������.�F�K)0�]ݍt��a�୽@�O���� �L��o����.f��+��9?* [�Y%H�E��ś�C���X��	ȉeXg��Z��+<��j�E� M[?u-�,YdyVQli�Ӽ��N�>�mo���x2�hSھWQ�zW.oXn󔾽����e�ݏK�T�����SJq�Q�[�̽s��k����Jn��F%����y�)N	���=ܸ�!�f�[�>o��F��qޫ��oo�\O�\:^��"O%�Z��v����5���h̐�Cd����L��_�^!�u�;���8+N�0L���ۊ�����y�S�fV���J`�d�#��Uh�Z�5�M����-�����=�h��#��:��N�u�>���ia�ꨬa$#B����[[����o�Z�����u�W��J(M�������/d��x���X�\p��Tj�$6�_��C[Z��^�}ҵ ��9�Y��B���OC��T��:+���j��|~wg�V���|��#�	�x;�Bw
x7W��&YQOv�6�9�G�����7��Tl�������2C?�>[=�9��p�����e3��>N��KI�C��:��:4��z��t�e&p��qR���>0p}m�lߕ2�wYན���YL hm3L��II��u��|��8�9ؙBI���I>&������mC+j���k�O!����d	3�n�r5�Ϻ��`v�:����u���.�j�ɟ;_A�}�Ϧ���Y&���|O���^"�5����$���^AD8�"�&�n�����< ���0��!��5,y�n�x\l��+Rp{ɮ�\��K��|�Ԍ�g�`0)��㐼����L���5�Px=��Ic��`So2%�6�����QkX��� �t�@��9��'4`I�	7��Ow>`�6���`�yq&��4^JUUոJ����@s�̌�O���]t��ސ
��UE"��-����|�v>o��!���Z�����d�`4����=�W����p�����PD�aZK��bu���)��\��ZW���b;�R��� �ͷ��4�6����U����=�]HJ�Y�o�l_�g��r����f2ǔkk/�j��t��H��~��{�����j!F��J px�P��vq,��`���K�`2�e����[���ir&��1�Q�D;�-CSi�&P����~8,7�Vow�*2�4���i�'��tZ/��:Β��׾'37�O��g㏓��VN�7�ժ)�Oz?���u^�+웂H���yNNc�K�u�����C=5�ۜj6*����s�0l)KX�폣~,���hg����ˊ��C>��8�N�l�K<N�>K�7/�&E��y�-��&pX���o�uݟ�}�.HKK]
��ևaŦ���Kv ��*��hrwM<����ଌ?B2�U�=u�_c�#�gƣ�X�zL�e��
q����}����'{�� |A�%[h�����4&�[�ؘ�=h��J���9��[�Y���7bG2M�_��Oۉ��x��6SE�3*��Xp�c�o033���Y��d�f&���_N��5�y�q�L�7D�wP�{O{v��PNը\>\i)Az!��͑9�(m�-@	�T#_3q�RgXb�RX,B�I��o�r8?�6�H��(=F��!�3c,ɵ��"��3%�||D����9��2��a{k�BFn���T7:��j7��'U����<�3[{�_�^��CX�� @�M�Ń��;!Y`4�� ���u1;��F�Q!v��2������*��H:��<�[���!�ɚf��w��F�����Ǽ,���tN��5��d��!���\�6Te�T����5�ٔ�]>�,��)�\�y'��Y��΄�kL���4q����Z��Brn��Ʋs��E)}����ime�ɦb�줜��B[�pi<pxs�>�}�4z���P�s�Z�{p-5����N����o��[CW��~Z���6�=�W�@�x!�'O}��.ֳ��pre������>?R�9j����U�)�<���-�;��q���Q�=.W$l:��?��'�ŝ�z��������~�����NW`W9O�涛��r�h����H�M���5q�������
<��T��Ϲ�=r�bCX��Me�1�bmP��˖��^;J\�!��>���ƻ4:9iԀJ�u͙�Xc!��8U@gAr<P���M�]�}��k���k�& 9�p"	��o��"8�Z�|����]��O��7^LY:,y�<I�&���k�n�!�{�k0o�ֳ�l���ʃ���Q9{��8�{�-�KV�q\�S$;/Ǉ�C��ݸV/�QewF���¬[���.l���.0k� '�����r�Q���9�Ͱ��T���;ǐ�[�����7dr��?���{�p%�z���c>��/S�//$~h���n�3A�{Bu^�5,�6���G;�)�����#��q藪"!�jN���h�Mu~<)o%a��f�E} ;��SW�Ij���(�C�t���" {��7�(ĉYG�T��,����dA��/����ZECؤ�r��"跙 R�95f�c���s�/{�.�����ǳח�eӵ�j��I6^�n���Y�����:i���mz�%��IX��Y��١V�\���1ɷtob�$�6ܠ�Š��*�3E�gI���5�c�na"Gg%:�.k�4������N+~���I 2|��/���X��iO�.n���a�s�ɢ�-Pw��m��bV��ק�Q��;GCt�֢|
�]��"hm{{��j#+҉�����K�?�Vv+�i�QA�6�B��&F>�Ke|�;���{&��V3��$&���A���/��6Ry���-�{R*�vw�B޸xO�$�v�n|�bޝP����7��|��,2���2�*�� ,�I�{w}��jP���j�_���Y��gH����6��/.}���v�&�}��Z���0!(��.�=�8^�1 ��L�{\y��WQA�Bj�ՙh�Ȧ_6x��g�@o!�ڧ��N�V�#:ء���y�bvu~XR��ƌ�춌��B47W5��oq���@�/�ڣă����_	^o��6R��:ۘ�'ȥJ�4�v�0g�����@;�3��0o�*�>U$B|bWz��/�'�����v�G�e�֑��̨�J��uA���O�v�O�f����6��B��D'�V
�HZW[������Pv��V��h*1��(s��Ъ�%� ����������?��r-G���?��>�h���p�������C�����&�.����c��u&���C���>3��3�rD��Y_s�m!�/�����VG�S�(����M��
=F1�_2�?���::|�b���4�Z�72u�[�^�(
�N�}����C�ϕ��x:��킕!6T۟�k��#*�@�͏""���?�+�&�&6Ħ1�<[�$�h�L�M�8�N���'���b$�^�'����:B�V]#�R遛Y,��@[�Q�q���=�-�dz�5�V�X��p���\g̉\�v*�Xɜ��s�a!L74rYH$\dE.�/;��[S0��P�B����>.P�W/K ��8:���L|�����Z��ù3
(���mB-�K_�E�|g�:Z�ݓ�f�Ul;q���w5c�q,�O7km�dR�����x�5���yB� ��rN�P"������i�������S	{ü�m}��S���+��]�Rut_������h��ܽ��Ui�(�y�K����sF��z�{9��>���Ԕ�����\[k��ϽYj���q���`	�n�>}�D�O��a����0�*픪�M`%R����g��V�s�����U�&wMN��`H�P)��U`u�-p�<�I~�H�� ]4[�LF��9��f��9��~�F����j�?&������ό�]Ϭ�U_���U�~߽�R�K. B�~v��lD�Z��@x<>�+C׵�VFnٷک�Ի���W��;��0��	>��>������Q,��}�]Ƣ��������vL�8���+у���/�.�g�!����m-��R���[n�t�_ma舩�W[����/��t�:<I㘶�y1'��o]�r=��%���֓T����p��y����*�_�kI�F�ʌnfTRpG��?q�/\�϶��(= �.�(�㋳$q)O������-4]O���k�m�=N��~8�e�M���;x5�=���L���Xt�j��g<M
�+�Z��������VcF�18շ,//(�����(�W&�"VE�\;\��@����O���xX�{߱�o�[�e-�[V�a�Y���G.�+vҝӵ�o6M~��i�U��ֱ���jfi[��S%7��H�~I��	�����'A��Ǧ#�R��:�,׉��$�M�!P�zW��\�.�����/g�+J^剫M��p"�X�D��uǭ�$�9��$�^��\@A[��&.=L����6�oJku���V�r��4�F:"8�n;�����|�Gwt���"�#	�;�^kh�8}���9�@{ʲ�[KdA�x���m��?���E��&�S ;n�Y+�˥�#w�&�Ԭ���ʫ�Ʃ.�NF�-U^�yW�@�)��<��`��"�|A���Bt�`�A7��j Y��=���a$�lU�h�N%�]��V���fX����h<+�����Ǵ4_�-;Ͷ�\�k:W��2�����'��$�F'���8�����̑.��ܢ�C%�P-�@�d��!������g�xK!��b5�8�ūٻ{�ِq�w�r��,
WgH�=U��Rz�Z����Nw����	���5����|SWɒ	Ev�]�*��C�bQ����hP
��)�?c�Β�Yۺ�K��Hv���3ʻ�kD��O��x�9���55��aU˧d���У�2'?���<����v��Nk�KY:@���TaZ�50�g�2X�-^�^A����c�J�.G��o�p[��2
,VqgE�Y�L�
�mӲ@Y_�B������¢�+~wr�fz���4���~��A��j�_�qv��5ÃT��$��N�3�13��	�6)@^�2�w��rX�LE��ݔJOnA^E+�n�LٗA(�9��u�pm��r��w&G�N2���i� c�m@ʨ���q�a\���5��uz��.ߥZ |}_[�&j+��{�nQ��u�Y3k<�K,��Ƅʌ��(ş�U*��l˕/U���je*X��:S֛��͇!���X�z/Y���犒��䤻�e.|��Hg�#�Vz��9D�7�N��W��XBREYJ�-��J������J���t_�aCVS�w�#��%oeI݂��p/M�zI�[�4�)�Wޡ��q�!��@�Xq���uC���4�F�q9Èy-^�-vA	�'}��τ�WM�x�(ù�s�q�������GmqW�@�*p��@C�)ς��fB�ھV�U��[������v���U��/σ���:���
���kp��O{��C��4����8%xp�d7��i0ʁ�����B��?�Ms̤���A���oX1Q8�$ۖ�Y�&K]c�BkF a�����L�W#���G���խ2�&o�GQ_�%?�P�_˸�z&��`؆�8Yw�f�]�	l�:�X �Å��C�!�Ä���ߔ�_H�M��h���F�V�IOw�]��y9�䪨�,��� ��Sq�ɒ=���A�T4���j����i�v7BfB�(�ϸ�U�����U��9^W��䝢y�(���v�ld3H)�zU/���A�>/l;�!Į0���.`�Rl��h�re���If��i����8�DCV��<�K)n��� ��.� �bU�J ~Qk�H9Qtzo�ǊxSpx+�T��cT�|P�qJ߲I�`�L���I�M�u�Pg��X�'��T���������c*���Y�O�ih�U��7z�#�@;�=�����T�Ԕ]�̴3}G�b7*��;t��Z�"�tTw_��p-]ש���tݹ5|6U�	tΌcwh����mX��`�*tHx�ܧ��ߵG)P ��1_~&j;P"�S##�3�Wd���r��E�*d���#��E��r��=��=Z\=���1jP���59k1�2~�t#�ɢK��Y鈯Ѿ�w�Br4�`_���iAj�S9SrG�]p��!Џۥ��JZ�3�V��X޼s+�7�����^�J��+)�I]\<�p�,�3�@��q����i1�������o������s�䂌�=��~nc	C�O�_��Z����*�i�k�a�&��ޙp�#ɱ�����������y5�'���߼M��*�d�C�ĢoLQH޷�*��U�Y�w�{?6f"�<�N>��m:�bnڪ��i���(��X"�q]�T��V��eH�He���:��ޤ�+��.�	�r[����LJ��L_z4~Qq�*?/� C�P�~x��7my���
��$�EyE�c��K�Pq��]\5�%+� �t����g�lR��������ǅ�,�V�B M�.�'�y��T*�!{��v4-[�/��z!l/2ra�$�_�:��p���3�-��3�S�ݹE�[~���C�"&��ރ�K�C�~�-��ױ��7Ȭ?X
/u�LK�'o'b���D�Su"�����u����j�Hx俁 ���*��U�j���k��BC�_*�.�#�|3��e<&���ֹ�r�JdD-��D�پ�ek(��N4���͞�`Z"�hh��7�1\�~�z����8qx��j�� |F@���xn����I}�PI<a��3����m�D�H%s�y��GC�i��y�2w)��C\�s�S-Aӂ�㖣��,4�����Ox�܊$`�3@�"���G��O���a6ط��r�a!NHRu��D�bv}|��0�d�~U�;��el��e�5�^)�	f��NX���|5d��@հI	��Ǽ�ܚ��>I����Wb�mҷ��������nEW*�] ����|��g�i�K�xb?2>:�͢$����ؔT@��,2v�,!�~�H1�
��)�Ѵȝ~�+_�	˥8?����Ԥ�z�sش��g�֚��\��˻��ܚ�kܪ�	���zb�PX��(����fZZ2x��ڭ�Ai�i�3���Ɣ2�M�Ue�8��Y-Q��;IS�,�$���X��ec蝶{�,����߶�t��ӥXit�9��^��6���f��<���<dE�f��\f���}��#���&�
V�W�E�5���v��\<�rV!z����5�ʵb��dT��ި G0��f�A�.�\n{/;��r+����v��+6ӷ$��{��`gC��&�򢵓��;�W�S{2���@J�q��S�� Z6ٚ��^�; t%�PͷO�1&�!0@��-a�N�n6����-�}��ꃅzvg�9�'�����5�]D�B�z�"�لKH�&[�bfbBB�$
��� �U�n� b\g��W��TA�p϶F�+�p?�Iss��l�eQ��e�ѰEP�^��9B�m��x�E���q$��{�_�_�����f��c���Cy73�@��dth�omzv���ޥ|'��LB���ܶGTDD/������B�]�+9@��9��@a�s����Ԟ�E@G����∼�@�l��|���L�>G�}��Adl�`'��\�b�_. -6 �q��fn�Y2��e)�#D;_�-w|��<
�$H�g�VQl;���~�����5�#���{^�#>?�K�f��N�)�r�7=���9	\ҹ�k�X�3b *v۬�m�恉D^[�����SARRO����Ԧ`wB�G�Xޠ Y���4)��ƙ%
�����H	I@��2�h}�$��-u!��X�r�+�و���&���b��l�'��$ǵ9�;d������/0�{io���a;JE�ܦ �/$vĞ :�O�	Q��ݫ(��'�v
n�#pD"�����H��}eQ�q�Gr���@El�9�̏��ę�K����o��=6:(hYy�l��1(`LC���Mʏ3Ln�݊���Ҳ �.F7��+�q�?�rK�A�_��"T�aE�uf�kR�.=2-ĸ��P�����,t�>���T�{�����B)�.��;������K�l''W�99	��|�|�T[�S' a��h<DX��6ڝ R'�;"!�� �-�s�9"D��(����[w*�K?���>�b��Zud4x��X#���0�`s��=��8�vT��_����Vht����H&-����K�@LF�Pd��(n�����]c����'��67{�p2P��~\'5�D٣��<����|
����\�y�J�(���=��gI(m�']����}�����u�?J ����eX+��&BP,���DX����}�蛨�>\�pT��7�u��[4h<;����τ��~ن`;���ء��NÙ�ٯ�ѡ��uܝ�`����Ҵ�tI������ч��ƀ��2ݛ�F���7��H���<tԀlx��@~����税~Gֆ�LQ�g���Af�ݏ� �/@>8sw�;�ڥPY`��%�۲��xG��%�/6h=55h��4�r�}�`*��e|o��F�:B��ad�lq��h�T��j���_�X��h`"� ��Z�D���[��tX�x��C�6����Q��
D�+�܇�������ar��jNԲ2Y�=?^F�F~�gV�:I>�,�.��p�����A@�\�I��@l�g2�()f��6-ѐT���_b:&�n�;�n2��T'�(�H�C�H��$�Q������8ۑ9'UN�|)�����}BG�,Ў����Eް�g����k����8���_����	q�E$���bף���m�^HBa��O�(uҏO��jt�JC�Oc�����L��>t��%}!��ofH}�/J;��M��Y֟�����h숴�����?=
���ފ��!���I]�3��3|�C�K�S�o��jM:��q����`����?��3���_ ԟO�*���OZ\V�JD?�PK   �X�X�l��A Ԥ /   images/670050b8-4f2c-4603-900e-28b8075f4ca8.png�y8�k�7~��]	��%KE�N������C�Ⱦ�R�ꤐ=YZ���Rq�P��/��/�ݘ�����8�������/�u�j���z��g��Z��2�1 Xگ�� X���+�=j���U���� ��G��ϓ:��uW���cs��9�����I�OkK{�s��m��"��� � �W9�9�"ul�Y.�Ov�V�Z�d$�ί*H:�y���Ե;�_o�њ���>ض���)s{��c?�������?�#?^ia� ��Y[[��/ﮫ�ŵFFFÞD�L��gF�O�w���}I{�^�w��+���v�^3�Rj��o �зov{�������ϴG�&���*��z���E�]?N�z�Ff[2�3�͂\�$Y�\�p��v��NL�
�U�aT��?i0�&��}`���յ)��Dt�� GGG�Ș_�ҭ���y�8�X_U�hʫl?�7Bt�$�Mр�o���)+�2����G?4����%G�s�
'򟌌��?98Z�	zÆWt�	�����kk�s�r������J�ok����v�v�G6{9�ى�Ze�Vf�ޭ'��F�L�����hϴn�O����2S�'i&ȣG���"�(�i�4�"��9;�����R��Ӏ-��~�],BEF�̔�X�X��H`����Ư���{j�-ó��5
OW|]���YH����dm�j�~��uW�Y�Ke���x@�
.̒��Ʈ�����&f�&��Y����{��'F
�R����Gq�۷o�V����IƓ�Ñ��2~��b�y�D�F
�Z񚠃�UVK�&(v�_���~�M�7��~�M�7��~�M�7����0�y1��?�v�$�g�+��[�r�������D�=��DlM�ph֒H���\�����+xJ���?j���ܼὓ��?8�*D�I��x}�eT�ī�~y'Wk����H��}���G[Z�?1�7��o �fZ�/yQ��/�~���_����������T���0!ʩm�}�gf�a��R�k��ƍE���]R�)���Q �i�K� ��]o�+�+x
a&���Z��^�4X]���1d�*-Ԍ�ʳK�h7���Qu
�mKdLIG�("|�n�sj�����R��~�9[)ܞ辟��?_�-tx��e?�t?a�]�ȉD�a)� x�`�K��S��'�������1Kl�|�����aHnj� (�I����dN�g�}�R�U�e��{���?B>��м���zJ���2�g��Ϥ��!�B���sfU���Ś�c�x�����C��]kH��!���G;F\�@�Ȇa���\���{o��++{�,�C�R;I�[Ӊ��2�y��b�N��L�/�J���άV�^[Jzs����f�+y��>Ȓ�m������/m/��WFF����1��'pU)L��f�U�SJ�bH�e �NM�w��U<":��D����"!)K�.e��S0�d�-�EBD$!䋩�ܙ��H�1�e�3�� Ğ�����T-�݁��ޅ����֞�Jߎ �����!&Bk��R����qШ�9�*vU54���k�F�+!�4�A�Wv%*}N2$h�^WY ��E��e��Iņ��i����îb:]hNJ)�-��G�g[H��g @�'ݽ{�8裇&?S���V��̸1�@J�e�R�4v!XBt��1���4/ba�c��P�_q�8��J�ӡ֢t�M��`�����J{'�荘 ?�; &�OW[K /Q[	�pw��Z��Qi]���>k|�->��q��Er�| Џ�I@,��5Dn�IêI������"����e*򊮘(��>\�L+of$�M�2U�儐6g�@��t� �o{�*� ���X�W)�.�'l�GA鐪-��1bO;��`�I>��&?��,F�w������ߐȤ.�F��!*V��t0�L��|)�q�`� k>�'xM;�h�� F���q�Z�n_�����)H�+�v!ZOr8�7���	e^�4^��:k=]B�77�a2�j�_e ��/���+��[�x���51��-�.=�{6~I�(r)�,
�+vv��(E|�,�Ξo�^7;��QqQ�P���2?�]/9ޥ�[]ʗO�˼s:Eq�!�t3j����I���G�Κ�M�P ����O�cn~<65�*0R0e�?��6F�a'�[/�g؁���<�4��3��1
.S�N%�B^�*%"Ih�$��%ݶ;G��&��=��T��V��q�Kz߸Rav�٤���F3�%O�֒�/���K+��I�+���[s'T5��D�0s��QKc &�ۃoi�z4�Z�5���&�a��He���MQ�QF<a\{>��n��F�]���os�їbƿɗ'���?�e���t"�"�aAP$�H���6�ᢍ_�0#�2a�k�'��V0fm���	l���	�"c<��,�|���c�5%짞]	@���;�����k
��4,���1���z}���Lv6p����J��+M�5�C�E����NYJ���1et�r���7� Ds�خfO���Y��"���*hsq���/r��ɿ
&��b���o�H�W��5�����l��8 ��A2o�+��u�T���e�;p���b���|�zP͆h�Q1�d���w�y�I�?Vp_�i��^uV��EЁ&F[�A�fs���ҷՄ��oM����B7G� 4r��eZ�^%���?~��x���� Æ���a���φ��g�[C˜�5<�֭�F8�*w�/��nt����n��-n$�1�{Z{*�[�My��u|�K��*[��.��"�N�	�GBI��z�Ma0��t���).�u+�="���B1�d�ǬO��1��u����҉8P�(K���DV�Q����K�3�'vS,fpW`T��j�v���pފ�`CǙ��W�p�^���X�U_<��ƙZ�K4�*��l�CTe��\�
��WAJ�#�A������)-�6�"L{���}���F���M�0��`�d�j���pb	_�v�jI$�%�f��O�'��gmN��~鄦���~���fq�\�iħ�]؋.�o٠�aPT��\�� �d�������W���WV�X�mԽRz.S/'��m�(0~o��;ݟ1糖���9��SbdBH�iz��	��4�a���/q��5�c�@ ̾��CFkb��d�;��ix�aY�#�Y[�ji�ih�yC&���/���HH�q��'�a)�RV{��#�r�U�O����ceo��$�q딃$�6����l�8op��9�>�T�b�vI�������M�N���U�J:v-2�~%0����o�} P�Zt|��.�_:`���+��?����?�%� Vi���\�cz�k��\�K9=��9�a<�O���X�D�!3�ь����P6E��Z���xLo��&�a�C8ı�}{�J�@�`�4�)7��J��7k�e��%�ך	#-���`|0��6a7�׿F_�۪L���\�NN-\��#)��;6���H	���m����.�*��U�D�R�2��)�B$q%:�a��>�ХN������!�����d�{?R],���~1��	���Zv�k����Y1P�C�9�Ֆ2��^��`>��g1�<�Ki)�VC��c��px�p��5q�F��̽maJf�����x��\Z͖W#�����O�১;����A~�
��Q���l.�Z��̮���(�t��%�u�y%��2x���E��+My�'�����
����o�V`F4�ݹ�?� �(���XVd�]/rS�����ۧ�0x�#A�{2��J:r��~\y��_��.��X�ש/��I'�d��1��j�Hx�UVnZxV�?�Ue�b4�l@!O��z�?���C���3�B�g��p�'�T�Ӎ�y��o<�Ѹ�1��`9�q��|\��znQ�񯑦�Ƣ	v
��]��D=*�2a�C�x�[ͿGK��^qD����.�lױ�ֻ�����)J��|�QFy�_Qv��,��(��ϥ�H} �`H�(��th\���1B#�wV��0
<��:�nE�e��պE��0��ԭ[u����T⴬~�z;��9��c��K��$���u6#���?^��L��XO���O�JY39$z�r@�e��&�W7�+��]uV�UJ^���R����T¤�Wz�+����ldU����]�ݪtə�XѬT1���93G|�].0ʃ��jg���ү){K�=$�*��r?�G�k�ǒ����>�4��YÊ��4�JX� �$���rn�8��4K0���e'�͇d4�Ϡ��
b͐Y6����u�����/��0�i��?5�3� �oL��Z#�@~��q��l�T��Ɗ��Y��V�ϵ/��.�-ҿ���K2�Cɀ%����b�
�7���;���Dҁ^�P(��a�����sf�1��_M�,xH�
z��]�xl�� GJ)W�n���pkީ��EGC��?>>O��ű�J;�VW��w6u?��T�{��'��l9��_�{�Mn�6>�st!��,rȽ}��%����vb�G&��9���ʘ��7o`7�W�3[鰼QJ��Ӟ�!��q��GmLj�[r�]�8��H��H��� k&<��[)Ɛ^��M�?b�Co�;��e��=v�HWF��ŝ�V:Ac.z�x���J�]��|�1�;���K,%�,����6g�>$����x��y[{6�����t^D��ύ��6��
����A����U�'�6� ���.����n�wGb��ۉ5�xV:[�P�±�)u\�ݮ*�5{�[�%[	sdφ-여4D	r���g߅��*�OWKe�DCW�W5�`�)�ƴ��C��s�ó;�2�����Jp�㽻;���H���#N�t�: �����VZId�+�)U�H���k39�����"*##�X�Nh��`+6�i�/:��<8�y�-�$�CqyL��l�rl����o������X��^'����t7���e�����3��[	�F��r�p�U��3!�m�5���V ӱ��_�c�W쎬�*��7�c6��}yt2NHr�o܈�W 8��T�����N�\,��e�6��/�_����穥� ���E���6�| yY[�}��]%�y)�u�#/��`�)�r��U�W\�>lA��y}0���S���D�A�Lv �G�F	���u�J7�6�.�xm��l�\9��7D������O#�؍�����E�N#�i[i%��t��".Α��I�92	+�c=�!�C�0�Z��K�O���$m�����l|�r�G&#��ΣBt��	,Ƽ��1�./'f=g�^�i
�`�	@�a��hBQ��'����Ei�v��8fvM�<�"�s���3�Q̺�'~���O°Z�<��ԋS�
͙f�S[n]T]UTe���1SUU���h�W�3������o��gRpo�j�����<�{�[vb�9�%�^s�,����Lc'S�%�"cBA�v�%�49c�Cy�Μ�샏g�<45���1���
{�k��L淶G!Y)ݭ�8�m�3�nS�QS��3O+�m��*�0��9�{c�&��KJ��.2�H�܅�f�9-;sD���SB���tP�����{I���F3���t�P�),�����q��rT�Jw����~�$I���ْ8�?�b�d"��$)N<�3d�`��`�l�ia�w�ǅ��,�>K]�'�<
YX�0�;�j:4�A5���X���]�)�\�DeN��:���H�t�U��҂��<=���x�tz�}����hX G�ݠX�k���D�u�}o!w���Y�^����ʼ����d�+e:c�U蘣��F�2x�@f�(��m�^��EZ}ѥ�y�`atOX���Ң$����X8!�t�2�&l+D����28P|�f���s]ܹ�E�o[h�mY�@U*�߻�Zm.��5v���r�r`�	���9����9��2Zݷ_^ѣ{��lC��;c��c-��M��̗�.^4��e��ga�[��[��I9U<�eCd ȧ����G�;P3�?�f�}D��bb}'�h6���V�c��i�#�
e����3 6d�N���M?w��r����~����~�\���~��̒~��I����[����J�cѪ,�SѢN ��M��W'Y������"���@O�04^̼)#F|��	��\�'���*�d���f�p�b��da�bv��;j���-թV�� }X�N.P'�[?.�^'��#u*S�2���up�����q�Ξ'�����p���� BiT��R��"@*�����П����Ⱥ�YÓ|K��cA���,4 H�d���R���ێ�"��uq2C7>�����i�ԁ��p�)�t������+T�SKŗ���0�E���*?��,���[�z���_�m��!RB�,}�|Ϻ��<��F�}��l�2S2߬���GY��0��n�I��ʼ�>`d��g&_����n���g�brX������8t�`�p�R���V�o�L0Cë^�����-H�l�_�'�_ލ�,���xB;<r�\݂23�CW�~�z�s�K��潄�y�jŉd24&���Q�nȐJ�K���u{a�����g��xhc�����p�Ɔ��[<qn�C��T�����@M�r?n�:���&�{,�5oV1������[O�S2�	�E!�;fDX.�9���v�kh�ِ�ꛭ���g6t.үo5�U�ɻ���N�t��e�A
Y� ����:�*Է��qt�F`���{r0����HI����̄�V�/E�{;ȋBc"�I i�BԍrA}�[�������#����{[o�ԉMx�ÿ
��>�_V��E���V��}T���V
���eӰ�h�!�r8e�F�A+($m�� hN��B��U�W��(>B��x��E!�^��=��g��.-�F	h�r	���FY{A�.ǻp[���Ӽ�D�r}���������݃MM��ͷɛ��� -��'�,���z�u�Q�HMYZha�!kD>!�lI�#�U� H�5�i�8������	���o��Յ)�,hD6��Ɣ���q�� 7�K��k"w�����Nns�\U=��9�m�%�~Pn��7��[.���{#2���fr�G!��[��$ļ�v��1#i�{���/��< �Z 3y3epuj�uFn$W4��?�e֓8�:����&)�T�?uɗ*Ll*�����XG���?��T�ݼ;���b9?���塈���n/��)P�,���a��$��K`F�
�pJJ��)`w��PsL�,FQ�s��Q����#��co���J�o��px���vRe53�IԈ�W%T%����9��h@Gr��qDc��b-������aff� !����?$j8�%���xA����A�\�l���7V��ei�)͢��m�Π=��s��_�e�,�7��oQE��fV�q& al �"NND̦�=��6�<�3kzݓ�&dץ�|e�A���/��L}�t�
s��D��'�>��=1%��s���;��Y�J4�yD���6g�DF�}���J^<0��Y��t݈Ԉ��������O8p��CWi`�G©@y�v�%,���$�u�X�?cH����p
��� p��)�Y��\0�ߖ!�����3fo9fс�rH�}�" �>����Q�'�$�π	�5w�g[㰠x7���u��R"��%�/�m�q�gVK��[�B���(�)?/ ]��©�8�j/��$��2 �i�č�VF�����e����(�2�z���$���/���5�sٿ�ҥ� IC|(�^�?�l�������Ֆ �|#Z�����QGD�]Y�ls�Y�bp?NNY�?��� lފ���D!h��q#���^ |[�D"Dp�y��̼T�I=#l���M�X�6a�ƍ	��o�h��6CJw"��}�!���e��j���]��|�*�F�Kt{*tI�$O�oX}���3w��722��y�����o�{at���ϛ9Î�|�8�Cx��F�O�.l	�1�p��M�E��,��ӻJ�c�uu&���������fg�x��%� :��$o�x�����9Xa& ������;�yh��s��/:1��<�E�%{���_��eMn�w�'1 +-H�Y�KO�*c�xh�����M]��y�}N>V��8����\Hs� fq��>���>�,eee��[1�]�$��I3����pW���Sp^s��ٹ��s�Fj�,G�.h�L'T*L6UFi�r$�8�T�����<vB��bf*B۝�CKf�M�h��s��e'3e	(V�e&��J�|���2�/GI�/Gt!��Km��m�2��х8��z���sҊ$�n�0:\�zc�|���р+���g��*���:�f��43�\�Hܸ�`0�Scbη�|ĘE��0全�h����Ħ
g$Ұ#�R�[|F�9J�x��x��Gq�U���͆�YI�M�gj,]N������H�wT�?��P����Z�ј]�]1a|&>>�ݍ8�S���4z�۫���\(X��5Ki��z_�h��֋�s�����R����>�nz"�qFM�4����K���=�E=�J�o�@��?��{�Y�������l�t��fMnI�xû4�'!p^v�eϫX]�p��\��ff�h���w�oy����;ٔ�N?��y�k_񙹗�yH����q{�v�� �����\���B4�.so��|�#wދ�=�����˵��Zt�r S����3���uʥG\.м����p���hMr��I��ļ��αܻ���;\�A����.�$�q�z����b.�$��րd�*�Z�?i��$<���V1TWwv���M�m��/���O0���K੖�n2��|�U����_���k�XB�C���[���=tf3��C�l��t���:D� 8v@���z�SQ�3Y!�Px�ο
�w`�~`���N���J9�h���U��t��n]�p��m���sݞd�pd,�#���ݕ,U.�ߟ�>���$@sh<���T=3.{�o��@�I޴�g�h��SLc�ǣI�(z� ��VB��Á+���/k{.��І�j���.?uNa�=�3N�W��t���γţ�f]��f��hb5 W���ڜ�GH���xպ/��QM����)Tg���D!��&��\K*
�Qz���
m�yg��4�U��'�$\�6�iݓ����)wgC�K��;��{[�/�:m>Ro��GE�^����Ar�_�����Eu�V:����o؞ڸp 0K_�F��i��h���=(�S�,�[�u���E�W�X?��I�� T��ٔ��%���H�Z��,s>�����J��\�]��; �>�<
9f!;�8nv������N�Wu�!vr�}u�{�^��V���DC��^�ɯ?h*����B"��{Ty�h6[��^����Pa��1�<ym,?���ڌb���K���\JV8 OI�gVx�!v��b�H"����=�<u��j�"������]���5V�oh��My��ho%�B&H�~��:�$ʻ��`���q��~R���[C����n��ڂ�jP����	^��V�D�(b�M�}+�������2�F7������8Wfhr;�"'����۞�WR���Xh�QZ0A�r[{��t���1G?�!uv�}Y��: _i!��T�EB����t��ޘ�Eά��q��;�I(��[�t]��-T�L����S
^��[8�޼v�B/�,��7���?Y���B���	97�B8`��$A=�\)1��@�����+MJu[J]@�*��d}:P�P��^���V=���B&��54�n��M�[W�O[�'�V�g�Q�U���N��A�5^׷j���GԼ ��2�v�2�+��x��WvI�Z��2]�yJ-b��H��S���ș[�����ul���`^��е7����_��Ey�TC��&6���1s���EL�wo�D�tG�"�Y�r��k(�@�dd�p��1�o��=c<� D��]:E`f6J�k�)�QRqZ��Q)m��Ff�G\\rS���>G�!#��_�[�R�-��.m��/�:e�J�qs�`$QN4�_]�u����=ֺ>{UJg����bC���́��!�a^s߾�m��U��I��r+�E�s���O��ObHX�L��wr�H���!��R�^���`=0Ie˭{�KA���s��rb��W�)�6��<��`���8S�X�����ɔx�gY���"��a�')�X���J+F�V\B4�5�A�	Y��"Sχ��#豗`;�:QK
@��z_�kl0E`�MX����&?&��4r7qD�>�d�������> I9$�?�I�	����A��0+�K�����҃�qRL��`ՄoɆ)�� Ƀ�Nru��ky���8m��	��A)�ܑ��˥��!uR9�&  D��OM�q�tq��a:�8�a�B>�Tu�c,���`��ST:�T����ME%ϭ��銟!��ϋ�^�B��	/��y�ۮ&�-�a~ɷ4v�K}�Ur����:V��C�җ<�`� �I�j���P�;����Vw�߸�"+�����(�#�CH��	WV�}e����˭���X?���~��~��_`�P�3A�|���q�����r
P �����2�W�a�q�҅��en.�[wi����v�:Q�G�{�N��w:�H�%zF�T)�(9w����|dfff|Lt��T�T�n~v"#�`��"N_ܖj��M@4A�U�p�����d��Z�%��A<��)$($d\t��T�h��fG��s�����R��쀰��N L�<�>�J���w��X������C�}�3�9$�:��ۥL��:�-A��Q���!>�-Wi�j�e7�Ub��o��7�������}͢uan}*X�[R��{H�7ܥ�ԇ���\]gu�}��Vb��
6�����oz�'N�U������sH����7v���R	���8���͢	1.C�XO�'+�Vt�c�,{��q%~��{�.C}�j��*yB
E�
��0
��{�z��1qW�x�۷O;�{���-�d�.���Pe�����f�|nv�(�G�y��#� ��x�)� �k��	;� ���[SSS$3!¢!�8L	��� @��0�`LK�����yj�>'v`��9T��Ӻ�H�@���uv�܅��4>(�#��Vp��Z�*��\� 'K2��� ����W��I^�>�
4(���� �Ox���ЃD��>y�
���=��4�B^��C��(h-�Vv.�^������(wikd�2
����d�8Q�L����J��A��&<�������,~	?��Y����t؊&H�A�&r&o�v�4 ����H �?av囪�9��g4������H���H�.��a{Z�1Q��!4�ˏӴ���l��R���D���4��*a�+�>��]M3��6꤮��	s/c�lmR�m��n9��>�h^kck��l
L�/�@��́��f�$L8��.�r�~�X6��c,��:��<h'N�x��/0v��ܢ��L�<U��IU���#;h�M��ɉ98�͜�ҡ���U�QQ��I��ww�z=�SHq�">��}&pO��h��U����a̍�K�-/F����`B|G�QASk�� �*���s��A����Ș��M �bB!���h�����:�������\l��'��	���0ӑ��z1=�\|�x�4f?�6�	��HU�	5Cc6�5eZ��g�&f����Η��/dZ�[��t����"T3�t�'|���R�G��q=�{��ɼp�| 9j��(y']:��؉M��oC_�<,�D��.��<��*�K��6󫌳��:����p��1WC��k �ҭ�XPa�3�0�ј�'�C�F��A8ȚIx4�.4��5[���Bۿ3�r��qG��s�1{H�C4��?�L��oӷ�:�4h���z������������;w^Г{A�R��#�Z	��s��kj��+���l�q1��t 7q8vE,��V�(�Rl���b��Q2��K�ǿ�架]��0�4����l�r�:��j�^Pf��c�=Q ��ΜK�p�_�5���A�2�Rl������D"����GϮ�&u�&��Q]4�BB���Ք7��ڏs`��!V�a�&Ѝ��{��;~�=|5�|��d5��<�����L�x�W�5^���>�L�)e�;G�	�h//�wy�Ш�
��O쉾��ʙ���^���3�o�aT��z�rM�d��s�,��hdE�����?�է�Z�#�n"WJI_o�1*Z�3�f�q|m��-O���^z�G��oJ^��D��꼺�wT7Rt
3_[6�GC!�N��VuH's�׈Dq:2�u�H�}P�x��ڽ�g���1�A�4D���t�o��qΈ�p0��F�#������l*��3g8h�kC�2yK[X��Dm�T�{�x�V�O��{�Ֆ���GaM|$Q�M�A�rL:��
�%! ���{9ƪR�[���,�|ӟ��XN�&�><#%p�����,�	��5y�oW���nt�/Tێ���]1��z�Ldyv�1��lja�D��q�
��b��Z��|N�0��,�qe��BL�jЀs�ۺ�-�"��R��A�W![� �q�Ar}����x��:=ݱ�W��h���O�D/��ѡm�
��R6��vX��mˠ	�FB㞀�۲�dh^L�����-�����j�t$"f,�%��.Zr��ZH��ֿ�U�+���,@��^��4�H>�˭G����"=pY�m��b�,�(\��,2��f�u��)�S����ƺMٻp�a\-�*ք�<�ů�����I%{����b�-4�n��2�{ ����P9��y�������M\^*d����ɉ��!$�������p�����rك�R��Ә܅V|M5̎�#Ǳi�R��!�����g��~8�W<~.�x<	�>�;�/��k=h��ভ��!1o���=G�C�	���2��ˍ��/���c+���9j#�����:N�i%�+d{O��r��Vy
�=�VGV*ɣ�Q��SZIFD�1�2y��M���:�� �ᾦG>�|� �'�M�']���U
������K�:1�FY&'z-��*3������0�9���-��� J�;ixQ���oM%%nF�� �}E�/�L?
�,Mo"q�u�r�u�X�(��qS	�dH�"��n���q�������ST;���AU�0q���:V��P�"кb�C�}p5���h���X]D"�!T��7��5�i����{C!T�zQ�*��<B�|�$\ѝԞe]�MY�ӘG P/_�:
�#Z�Z��W�a\)�@����5�v¸:\���q}'����&9�ڐ�ut���6�FH���m�ز=������0�4X��*he�!:w�*u��ixэR!����������F ̿rj�)N�8�㍑ST�,k��a��>r����5����w���J
��Fo집�ǂ�Fߤ��ce'�[ƽuSfxL��'�C>�����mA��z7O0���K� Ǯ[N[C�Ou�GI��O��� ��gp�(1�tuu���?�YQ|:a�x	��|��lN�gcva�H�}=e����@YYY�sWi�R������+��������M�#���v�@�`D�Z(���".��eDR��RM"qFљ���.��̪��*���:��L�n3����#����]{l�[��W�x��+����;��A<�
�d+߫Z4�j�ꩴk��G���4L���qw�L}g]���c��
E9s�U��C!���'�,�����/��+�󘚚8zn�����H~���2�BfM\OW��/fP�~�f̌s�,�Hb��.?�)�`���`x,g3����j,��H��٢��E��ˤ�ǐ7N���;�����u�+=О��  ΃%P/�WN V"k+US��B_�S֗Q�{�K*�9Bc�����׎�r'?�0W �ǵ5$
�gr�_��v0�z�ZBc%�J�r��g�j�Q_9���#�����`+�ty$ڕ��vN&��/v �����S�6d�� 80��"�Oz��P�X���;��.|�����x��b}��n%�"���k"U*�Iy1&��2�0[#g��f+��������b�4��L+�F�ݭ0Q���.��q>`M����iF�J��{��I!�R��4��ݳ���31��J4`쉐W�k�c��pC7 )�E[g���J�5s��#���"�㔶�B�8��t4��\�=B�������]U��#�>�9��d�*���K��^��|p�p�n o��ID'�W��w�}Fr�#2���*݄,��Y����*M%R����\�Mh�6K5�ט��&|��Q��s�C��I�5�ū���MrM�L�Y!�t�M>�pc�g��	Z .��s=���^���v�O��ק�q�N�p��V)��O�z�����`���zPzjb� �NƸ g��om'�Ok��������h���}<&�T�=����"7�<k%�ۂ��a������R`�1S��!�k:������}�Ki��G��y��r�ouk*������g��,\2�p쪌�ښ3Ԟ<*Ο��V|}c��4@)g�j�p ,!X�O�xjLo�������g�I%����fL�0u��\�
M�u�L�ޑ��?;�5������VM1�D�G!YF�`9d��q�$�ɫ"F��k�cM`{x�X.��J����}�\a�J�z_����h�*�b"��e��T��u\�c��S�q(�������v:[c(Q�m���m�+�nk��^('���[��((�-v���e���_эr/�7��A~��Ԫ@����#C�AR�\[:<�rd���إ���E#�>2�P�ïm������pgfؼOe8d[�#�.�zB��B����sXh�2GϹ/4�'��]��l`�!����)�|1�y�܎��"��4o�@*��3��p��Ek��Gp�N�/7��6���C���[n��?S��� ���ɻ����9w�����@tƹf�n>v/eo��a"�8J}L~��d5./���X��TOؕ5�:;���������/��M�G��p!˴��q1���҆��a�k����9�����OVo,-��>ϗk��֓W�������g�h�i��E�8-W�S�S	���TE���<;*�A h���?�H�V9���H���M:B#:UJ	!�	Ӈ�pt�$�b������/���6+��]8�ñ܊��>ytI�A�S����hv���@�U��r7P��5�
�УZ�c�BѼ���r��������,���7�f�*r��-�������`�=�T��{������'��.�YP�i"CY�Y����+G*�3�}'@Z4�dR��$rL4�^|�3)��u,+�R�փ@p���,�3�9�a%:v��bO߶�vN����i�c���ȼ��[;����+�"���y2+�71��d=Bm�?\��v��v�~��r�3��̈́��Y-����:H�l/��[{�:˪�Cg��@Rt�~�Mp�惙�\_'�f!�f$��C�IA��i���E�i~�+Hfd�7ft�B��:��=���ކq��P��J%�D��!祎�\�~��F�\���@���x.��ذ�]���o�7/,�3�xu�bFձ?����N����*�(�հ��0��:T˟A5�S1�OMW�wPծ��=:s!��v�P;kʁ������!Q�8Vo�(�x�d�C�X���\XX칋�	ӟ���f���){SeiJ�Y���oȞǠt�� -��Lj��O7JS8M+0�p�~��]��t>e�Q6�0Ԙ[��|�I	� �:��C/��.�Q*u��ϵ|w��#�n�������+���u���� �J��~=�\Y���M睨���lǼ�v�6���g�ܥR-���vR�k�PI��]L�|K�=�`�e|�$�'�������H�����Ut��v@���?K���.�K���J�~-jP;�ݪP���<����,Y;u�ݧ�T��	!��	�%u|	jױ�]6Y�`:��P;:���AI%��%
�����ub-)X��{4�Ïeu����^+x*����2B@Cn���İ��n�D��D�*�� �Z���B��7�[=��������uS�Γ�$�6�#���T|��O���A��V�?��֩�.�#�6�������o3-�Fmf��άt�"e�z��+|q
J}����,����I%���?(cPu$y���z���>Ք9N�vW^i�b���B���jx�3�����ڱ���f�M��iIA�Z����o����-�Zd��ǭ��s�y��Ǝ��awf�m�?��m߇{)#�%��G~�K�1�&�/��}����}���$�Zr���μ���uB�����KJ���������%�jgtt�����\�N�@ъ���=�Վk���!7*F�,�L�K9�^W�F����dj-�#%�l�M}��֝TrJ�)t'A��R�..�S�7$\�S��vr���֤̯��Jw-N��t�:!��W_f�c��#���1ڮ�>�ü]�>N�9ڮu�e�rֺ�9ǅ���f~ܕ�$]u���v�b1��pd���+���9�rI��V-�)����O���sQ�gL3��nIyvb��U��3v�*�J
1
�*4%`�*+�,�<���h�w�q��=m�S8���atK��,UZ.����c�?3�!��;9���噦��vۚ�9����,��_	N���|F%��|9�.}1ƹW�H���&�t�+��b�����Y�&��MQڷ�u.5F4aE�N�\������֖$��Wo�l�,E|)Z[wU��b� cl�_ϫ�~ @�S�g�()�8H�h��gs�w�iC�x��m�ƶhk(���E����~������bۓx�o�=��z�c�Qͯ��=�X�zY?���_�U� �N�V�l�h'ͷ�j
������U�ۮ[82==�E���h���~�Q�[4���pM�
KL'��(M��=�%K܌����ivm�z0��0�Ж��q<�ݣ��~���W��{��d�_	�h��5��o�ភr<�CZ�:�V��+�c��L4��L�J䏖�7%T�1�{���k��S����*&QSc�Bn���<����(�?R��.���8�QJ��q/�^�<�,U �� L������Pf��j��C�b�-�^C��1���c%G���D�/�������@�����f�Z��,��*�9K�N��cӖ/[G�9�yt�	9�y��U:ctX�b�"D�"�옥�����85-�Q5z�ݤ畲ϤV���v�+��7�.�2Dyhkq���!Ǯ�C�a���Y��t�`#z�rM/����$)2:��[�O��O����n�a[D4N��,�p�3��ӧʢ�2y��͔xi�T�+����ГQ����8�y_�q����w$b�%�\�q'*:�p���w��OQ�̈߶-�AA�X�α2������/����SYB���<�����~_�+������i��AW��eI����;��A�,����	\��DBI�}~���x�_��kA��BL���D�xc,�������1�f��vVay����S�!fq�-��"��R����d�m�G\6]|��;⿅��搊��O���~�×������y��AE���'�M{s�ڃ���YE����.�%5Ǖ�^�V��4D��f䘦ޔ6���ڪԳg�������1i2���;*�G,�"�s.�XE���u1�՞n�n��-O˟�J:�x.w�T���5
���޽[���}��)a�a��o�i@��-ьǕ毾r���&�6/��U;G�;g:��I4¯wb�//�20������bf��C*_�hɬT��Qb�L�ad>[�mK/��W�"�mO�������3�������,d8�i�mo�>#�o�?}�f澭��{5o�����U����I\�϶|�`��5�3Q��F�T<�?D��ǿ�K��CH�*����ݚ??d�>�R�V"�6�2���@�Yk�q:����l�v�z�<�`���m��_��&F|9yK�G�=z��J���ѣY�;�f�D �anS�*Ź��rg��)�������9^QF�}	f���0!A�4\-09:OOڐ&GS�gSn9B��%�̝P�H�u��ɡfR�{�T�G�/�q�a�jg�mz�M���/>j�o4&�y�y8?�㪇.�2ݠ��F�������O�L\�v���膃�g��8L[f������	2��ߎ�l_Ҝ�p �yQ�C�{�CVE.CM�E^,On��h?\��p�H@���VS����\4�!v��6�A�զ,<FPr'B��!-�h�l�����؄	�qJB�,#�8�7P��L����6�怒������<4!�;���A�M۔�"�0D�6��l}g5��H�}����	��Jӆ:it[�K^��=Օ����?��ۮa�t���W�u�3\]�y�l�g�?�9�������4�B�혡\q���M
����u��gn&�|@4���c�?ÚZ��Q8��5�� �(
Xh""-`�� �t�	�{�P�n��( %�4��KhJ�KE-!�P�,�o�����r����}�/!Yk�yf�瞕�� ]>�������G�k�����ٮW��8g�o��o�u( �������D���ƾ����Do������ml�rN?���t�Yy�c�Vw���0��e�����O�	Z��ZW���'�B%oķ�'H.Vo�o�dW=�|�=�9��TPR�A�{�_m�'��D�Ir�m.li�ξ��9������%.	K��7�>[��a��[Ch�Z�m��#�K�<���J�����&�3�Y�=s+�G���k۝K|]���/4�o���N��E�ym��?�C�D?B~SR繶����&�J��Զ�e��փ544�F7+	r��� �����G|��U���K~������
��Y�5w��^{WW׿N���#��r��%a�2R�[)<t�
Ch��h�F���)��%��Pd��ERƛ�{�D`��4;j��'���X�q�SZ�MZ��g�������Y�fm����Z餹g���?챛��g[u�d6�6S����D"VW#�xc���CCCJ�NXH�㋖?#~!�U����[�
Us��n����E��х��[�s[�:�{�1>�7F��a�kK���]��[?����|�Gq���:���1�S�k��4�v���My>���2�{>kt-��]���S�H_��������u\v���38"p�O��V�4�0��?�6�9Ԩ����F���c�,uG;�wܷ����[���<�1�dLj)�׮�L-'w;z:FM�o'�<ő�?�j�?P���n�$�lvß8]����D���/ے�ʭ�V�}��L��=��tn��_���q�n�]+�q틸Y1��$n�ŝ`�M^�Y�u[!�F��4��|��y�	��\�)��l�ժ�Μz5��q.R��}_�?b���%⽂'�-..� �cpZ�o-�S�t���r���K�W~��׻ۊD�缙}Vk8�{�řQC�3ٻ}��YVh��	 o걒;ϴ�?�i��57�YK�J��h�[���Բ\wH^��*G4�P �����!���_�ۣ~���ߔD��ZY��o��
�����P��sQ8���Y��9�/��&�L��.xݍ���� z_Ǯ�ō*�^ �s��wO��P���}�<i���ߚbD�6(kg���:᯿��]�J���i���h��m�K�m�n �e�X�&	�g��[�.>� �ڿ?@�k����I���5�-�!�3^�oEW�E��W`�$�����q�|=6��֚��F^��]�A�WU�fDHz��Z\�(�N�
�Ͻ�9�E=
A����Ӣo�Z�E�,�>]���}���E����ls�TL�*5y!k"gࠎ�U�70����C�q�~u{�S,��h������ڍp����f�E�(�n;,D�7�w{A�inE����n����Bz����(�s3�x{�+4皝��w�5/X1��ٴ;�������#����W��k"9��^@8���}��5�`+T���SD����

��SȨv��8��g�l�J��Z�(ba��%vW������t���;��p?�(���e�^�CKX5{��8ב��CV7�(�v���:Ғ7���zS+�0y�o�S���s�E�dI6�,Z ��g(P�V��P����E��"O!>(0w�ϙ�΅����������-6�w��L���n�9v�O{����m9wo��ۉ���߿�K���'�.�g�?#����F�3����g�?#��F��3�P�y����ċ�'�ط�R�6��Ijut~H���	����4M�XKN+�A�U� ����i�$a�d��I���"q�諩�7^��z�:��`��m�J{��^^a�;���R���53o��8��Z��Q�2�%���I`}n�/��ל�[��*����_����{��6�}2I~ڕ�V���oa�J���H�~�_N>�)�^�ql���������O�Jb�_�NR=Y<��Ю��k&�p ������ژ����.�pv�Q�7Y���T�&Kh�Bͷͣ�����\nU8��T�ʘ���gB�.5�V�����W��j�˯GJ�r�G����������9ݹ�V3��C��ek��7����멒ٙ�D��j�P7�V�tO��&E!CJ�@���9UW����;(3y��1�\+���c ���V3<�s�b����/-+{��kT���P�J����gB���	��y�颡�7ɐ�t�
=���l�S(aSA�Z3��mfK�o\t��Q�P�c�wU(˞�y�k��FŝC��`"ݷV�d��r�:�:�F9�*]�� T=��'i�R�j�'Z����#ز^p�
�->'�#���)��se�~���g�.r�`�w��8\+�\��������b��4�:m&<U��j���O���f�\��;����{_D*rO�c+�ttu�D;-N,��`�����D�&���&��A5t�x"�����_P��aߓN�/��O�9��7�{`��I^��R�C�^�c�W�
i|vltAS�;|�����򲺑����A��y�?�3��knetyY�G^P�a�*�<�Ȅ�E�H�q�8{��b����s���e��K�rǟ�e�����p�*�҅j������SoX\k��d��ܔgG�M��c?JB��s��<����t%w}��#���v�eC���}��i���$C{�N�5ֆ������}{�L�i�b3n>�`�!�a����1A�'Mb0..<���Bݽ?���c9�����D�K#Z�w���$Sg�o���� �rhd}]Se�k�R����<=�:-:�ޣ��3@�zT�	��k�SRo�����߯�ӽ���f�%�T����ȸB-7�$�c��aӒRR�0���2�Ҕ7J_/s�\۹�0dTIT���t�c�K�f�f��]�d�)��7��K�V������X�pr�����nX�k�K��juצ��&���<r�d۴1�����9���Q�|�ԑ�Y��d�=��E4��lջ1c*XgȨ���K���Cy^E|�r0��k�a���:�P�7|r�f�ᑁ[��N�TUi�DOEjϵ�;�D_ǜh��#�Q��7�i�l�TŐe!R�9��R���<��.��V���-�e,֙X��:,�g��(�wؖ�(�ԫ,��\�RxP�8�3���'ɞ�z9�9z���TQ�P���k��. 0u����P��Z�u��j<5m��P�?�$��6s�7�H���q���My��	��Í�m0�k��>:���o���
}]]vW<��}� P<==�Ե����'Ά]�pJ���H���'�{g�U��@+iʃd�ͺ@d�NC4�~A����G\�VT���`|JM��~1�Y�-ڌt�����45D�o�F2k��-))��g�Eo�=�n����>���A^��t��6ǰ ����K�_�m=�R]E籢l��/ь�<��EIE��xui0:p�&�Z�E]���)��f�;8��H��� 5%��5��NI��{��f8��kv�N�H.��(�� �q{{�B�����L'ozKW�f� �P�D�Pg9��
j��&�����]j�~�����uN�B����W�Z�x�����9�h�Na���9V����^�.0�Kqi���Z�����]�}ֿ%oF�ɯfXv�Q��� �X���|Î�К�0�]I�	=��h�M!9=���Y[{�I�������N�n�@����|��y�^h+��^�@���V���,�rWY�Y�%�ע�C�F�ã�
��P(Z�@����W��{/@�AC�">��I��$�>'a1��qnn����E�=�<MZ�T�P>c� HN~ ��%B�6����	�2���u�ΌP|�5���l���Jo�؟�J�`�4��R�qr���B�k�����P�VK>]�r1]�q,��������	oUE���LH_����h�~U���`%<���j������'�ʿ?]�G�ru��:,t�a����J�Gǡ�O�����DI'��⌑v��y
r����п�y
T
}�<d涹�\�E[�gh�U���2ۧ���Y3&�X?ܜ�#dh�'}怉�D��I����xG7��U#L�����5����x����-aqǰ���:p��5 ���eޓd�3c(��5���`hnd29��\*'&x��e?��t�4�-�	�j u���&!B�����H�8AQ�����_i����Ʀw���X���ZC t���9��>4j�@���oo_��w��treH @�P�������
�	�b�vV�B���n9g%�t��G^"���oD4r�����q�	�QFX�3Wo��R������ߍS��\�.��wb�GC ��)Oi�6���m��cSR��|/uo�D��r���|�@ h7td���ʆ@�����G�{�!�jTݏxE���P䌋����|4�0�uLrh�&�c�El��6$Khh(�������Ƅ`���n`�9���Ŗ��ݧ����wϭ<�9eS���ܬ�s|o|
N���(��U�%a�E;�: ���h�^R�=X���W�&k�U��酼o�������
�E������?0�zI��p�^0(�%�5���䐹o�)�����������6�0�|���Q
��Í֩�	(�g�>]�>Ud[�o��_$�!�2QGC>g�)~�L��k�@:�.;!�l��a���;��j��xM��~w��̸�Ǐ��	+˔~����d�s��D�I~��CO��ϸ��f���g,l-��I��u+$$0eߑ�AX�;KO�bn��� �	��^��CqY � ��/m4y���/H�������mr[0�_��aq�ܙ�A_�F�Eg���S���G��G�y?�л�,B�:���#`CLp"����gUg�G�}qk``@s��7�i�!��`�/��ܙ���NO���t��#��mG�B�@� ��q�ٹ����[���~K���5{h����(�^3�}�7N�����>��ty��p-�L"������d:{J�:k�6�������:��7l�ۅf��.����~B2V-d�/�S�Y/f\�Hp�D�SR�12޸q�0�+ҹ��,o��r�g�5�/H��j�`C�Y�Щ4���#����a��7�wtlݽ�:B�;�j%�$��D��*R�x<M��%��Z�4��"%�~��g5W�)]V��=-J�S��dP�E#1�PQx)��t�Oޮ�`��#�0lE�z9��i�t/�C�.��&���aP*N��=(�޸wu�;LP&�m,f��~���ZT���p!���~.�-��{fv�@��u&i����O7h0褠����� ��A���E�v�(��[_��L�"ѓ��������FA��H8�i`���F�sc�3F�B{�H$:NX�H}TD�+���C �0�	�'F����@q�]���v��u��Ӣ,��ŦbPdy�9Z)�mn���m�x�����n�S�En���������g�@D��ΠZj�DTb�)E��O�D,�<Q-� k!�C��""[0O_9φ�Z�'�o�<7`�A���r��W���ߊ��M�c��
� m�����η~�f�"�#�����Q�$��ܜ0Yt���� �$m�mI��"Q��j��%m
��zbjd�� wa���4�8J;�Y����%��`{�h���X� �hP	Pq��8��ϼaeD>vx{��J�1��>��ق��~�*�AܕsV</a��PZI!\�5$�����Ċ�ZN�\T)��~����ip���qg}����Ǧ�b��"ш�1�<�P�|<���/�[�X���W^�$m�`�2��U�#�J��B��GEu;!R"8�yLƫ��8�ķ�&)���4U|Aa�:�ͩkc���kX�#"����ƢG /�Տ�i&/�K	��ꂼ�|i-++�x6 ����t�*���	�5���JR�1�DY�v�F?+BJx+�m��w���S��e��<���'�A��N�*R��,��W�����+�Z�h��Q6� ��x-940C*��7�2��3v������;�RC�a�q`�j�@��r�f��xB:�wӻxX�R�	$[r� �B�(��`��~� :\.�et�{Z,\>�|� ���/���� ���UK�V3G@L�ڰ�p�6�������Y]�:Z;ȍ����{9F�B���~������XlzŶ��uv��W�ώ���=��U���c��������J��L�.0��f�#���~��j�j��v����3��+軗	�rߤ�_Z��6+����Z��d�Q}
�0Kx��Vn?���^�o	�M�0�#�Tw���:����s��x`lG�(������f
<�z)����6��csCW<V�4FZ�ۛ�;�+
�J�� �͸��k	)`���j�O����d��?i�CW?�f���d�d�� �Rg�h:ҥ���@��h���%2�+GAL�/��L��U(Ƶc�$�eZ�K�$�t���s���b��pl�Ed~�ǫB��y�I����XVT0WʁZZZR�����P)K�;�\<��&�QR&���Uj��/���th=�ܡe%R�@2���Vd[��h(��K�u8��\�J/Z�1��L��U _35pXC����l�0�4Bb�z�MN����hM�<��)�\6<��0����Z���i[A�*R������M�1�X�m�Ԕ�E�#aV\�ΠrS��4̥��Ol��z{g;k��t�F<$7u���{[u��@t���}�j���nA<q�5��)����EG.�Z\�<�(Z8���o)��fvܝ߁n�sn�.|&���t���\1�s?�=K���bW9U~��4gi��'5G��b���3��C�HO��Ԑ�B�!tO¯�6� �9�����γ��Whm�T�SE��τO�\������cc��K6�w �� |�д��q�D��Dd���
�Ʉ%;�Lkޡ�-1�>9�Q����x�y$"��C(�H��$�Z�,��	~�P9����p����:z���!A{nJ@5��ڈ��8oYu�E�i�u�;{�aڙ8	�����-���8Ø�s? �I���CE�-���øv=�b��OY��JD(=9ɹ8칂z7���q8�����Kx�f?����
��EW�n��s���t���t:��A�;��>�)N���N9�":��\�󙌼THq��F�K ��?<.B�>����tR�!{
��Ru��4:���8z'?X�~��Q>ц=[�J��{��9�A�n�ä^��X�k��5�ǟ�1��i�*���u�aj�7��ɨ2�҃te���v�y�L%5'����e�������,y�twPO�����w��;��?K�+;��l66<��t�uw�2K���Wx��k����:wS��
�����:��.��&5c�o��9����1�=���u��KT�̘��i��f�f-��ET���ݢ8}p�BݕE���70m�Ag]�O�0�2�gs�ƢSw>UؔxB�욦�����j4��J,�1��v��XhݬK����XqO��|�q]�nY�@Bt��������h*0Pj����~ց����
�UUs�cߜ���<gϞc�5�Nv����."��8O6��|��E��K��#S��a��}d���� �P�@�P��xL�����ɜ1��򏎿5�ml`,�92���L+b$87�bNώ���u��n���I����Y��$~�F�+Is�H,���M�zGv�N���M���O}&�" �	S��W�?�x�͞�����Y_X�>�$I��q�;Ch����,O����-���M��K7��������={�¹|�b�wQ����SB�<z�-Y���grk�8�mx;�IB�zO�4}�q��!�2�tl��eS��B�	�zLSb�cPu:��R�j'��b=�Dy��꼫��DON�v�\,��Y�iK���K�����_���@_s���~�J���G
��ز���D��Y��&to=&U3�{�1����	@�<� ��N��{�=�l�a7
w�$�3O�����t�u�y��߻0My�6@M$vOs�o�Z�JZgsnME���{/.��z� fR���0jV?����������c��C&�Sɍ�Mw���>�`��o�P�J�}��Ζ*�Ň�%�����N�V�!�(r#�s-�u,��/!�MR7���h�8:w�V� lhh ���[ �,��>d��.�\�A�,e����d(��%e�����Ч�Xy;:&�e����~��������G�f�vϧ��N�^R<���`X(ђwK&_q��һ�\�x�;����`�x
;��on�<���D�d�HL�k�;��41�(�[YBH76v3�ӱ��M2�M��s��UD#�T�T]�=]�$�e���m%�A�	<��W�{�:���Z��Nv��˟�G
����j+�?�������_�>�t��By>+�7�bz��X���{"zȯ&,���K�?�Nr�d����$�lQj��G��:>�5���}�ΔXZ�\bXh�~�p7���6�8���xa�6j��B��y�˥�1ձ�c�F����V�T�����R�.M��3�z�7zsq��ۥ��yv��2_tu�N(��^(��ޔ��q?��\��/�OjHh�7���l��5yFj{��h�@X����p������}�]��g�kYj/�����~��^�{4j(�ٱ��J�A�,��A<{�x,��W ]�/��������T���k%�vQޑ��9����E���R+.���u?C�̭ŮФ��r���`�z%q����p,��C �X;�0*%�������D�K;n�����J�C���jL��^�|j���U��L�ΑM�q.x�!#�'����b�3���.��*H�~�1����l'Zߨi�xbx��}<�o{9H;�Wr�*��2\u�|��e��0'��Nٜn�y��x��w��ٸk�0rZ���т/S��ej[ZB��>�gp	)�`�ˤ��ӱD��׳���`F�(�<�"I�_}'�?@��2Z��������/�Z��w2��\m����b�S�;o�Ƹ������%�P�R��6�"gړ{��*����/�_�?��^�sC�̽H�����cB,�[���ޏ����R��Q��A��8�:kp���8D�+���]������S�Sb�)z9s�.�>���C?����uI��-�N8����]ɳyK�͞�� ����=6;�^7)�����Q%�AG�x��I��)��U�+�(l����SY�W.��|'������%�վ[�;��ݤ��cѢ0�x(V��5X�c�榀Q���ǣƙ��îlMQ����&��xO��h���̈�(�#�Æ沼�=\�g�U2��^�a�(�Rk 诗���*�dف�'�ܳ�����X突3����}s��U̐��MoPVf��F�{�W���f�%�f��d��{fΔ�S>wZ��j�w@��X�ܱ�7�Zd�_{��Y(��RV,�?��2C�r�%x�-{	d��	}�Q/�����F�-Ϯ��ZL�^�'.���qq�T�T��H��V���TO�Қ��#���������cZ�N��aѓ�]ސ�ja��x&�Hn�=(s��}Rm����!t��_�>^�����% �4�b�!�}�N��V���_�
�jM�R��Po�������D7k�` E�{f�����dzJq��|���?֒�j��`��rn�cr���p%���W�I�6��+��7�����<�y(r����ڦL���'���T��e�{h/=���5Ra��9ob.����*{L}xDȲa��A`�Q��Qq���}8�������W�(���o%r�`}Mf�`ݻuA[5��l��\B!��p����8�L����c�l�/{ْ��J�c�":���z����!���2ǵ�w%s+Lb��ar�����g��w���Mc�&��^L�lP��j�B6[\���lQp1�D��\��u���V/�Qz���%$��IR<��v���/������a��a��F��Mqa��i_<~��0s������Jؐ=����_��&�:��p��?���� ��/�����A뉟QIz�J-�/L�����U��u��^�[~/HW�$%}gn�x��}���=��� B��ݩ�/^��G_K*Ny��o���.��>�����L_����	zh�Nx�L}ޏX����9�
�xʹ�a���
a���`,讅�N�� E��o��c�y�4���hr�;,��0��z�O���6̍DV��H\�أ����/l�����P�y x���~M⫖���0C}j�� tR�T��N���Ř@WZ�[N�ck�!���o�Ի���κZ�g��0C�荎	�����i����f�ә�Th��©A�����<�/���e���;� Iヤ�z���ز��"ts�͕0�P˻�E��`E/���aW�U���[\kQE�hш��3��
>FG+X=���v��f=��k	U�Y�c-w�=��f-�0�60�6�l%=��	b4���ߠPۧz��6=åƢ@�eDN#��4�6!��T��&�d7�;�⯌��W���.������x��54���4�y+X����8���Z��:\0lU���S�#�^*���n�����g��:�>*�D's����"��h�d2,kh���Z̑�()>������{4?*r�1��$����������_x������4]�"��Gzu"��Wm}���2��#r��<}�����s
���*}��kg��c<��&� ���c��������\�Q����$��ɓ'����1����t�z����^�������ɫ�O�N̠
�*�F���d@^@0�u��Q(�k��'D�������PnII�D�z1=��ɕ7��\Ԙ܈�g���ڮ�݄]�Bk\��7�9\�q#��������fi��Z�t��%2"Jd��4F�>����έX{��z�ѽV���.�>|�ނ����z	tr@Nfltt��7�_4^�>� {�P�-�qQc؋��m��˜��&9��J{Y�8��Tܵ�WY��Yy �u:�8��o&�� :(9�VOd�]%����J�����[%2�0�3�����l�
�ʓ�S���6����:��@�bZ��Z���wQ�ǐ���Esw��苆g��嗱�
�����
d��������?�#)�Fi]Ē�욧�NB��{�}��,�ћ7��]��y��2P�Ott�t�#&"���:� Вx�����) ����VK����j�G0q���6L�݄��gpP�s 3aQz>0ۤV� 5��{fX��y�WY��L~������	'�P|AAR�D���D���#�FFw	d$�f� Ul�\�X�R�����ojiy�}DD�m{���[lj�9�,
� Kdt����h�ĕޕ�w�z��y%w��JD�4pw$ƼkQX���!��%��,�5c�<��:��ŻC�.�d?�:�_���3��`O۬���TTT������&�8����̉�K�f�����C��@�
|y�&�2��o����O�.ԶpA5���idtF�[��66<-�A�Z�δ:����|�RU�7��^�k��,���D��B��B��Kj;�=�V
x\DӘj�	��%�	�"Xj_6�<��K������/�ײ�pts�笽:�I��K1˹�}58�\U^.�O�i�r20���U?;
�Q2���n����OI? ���=��4'��Ʋ��F���,g�ҿ��T��G���c&9H=��?4��{�؊3���t�l �[,MM�7��*6��;(���.�r�D�miQ�MN�Gh H[�͗���v��|u@�l�Nw'Z*Ox�����gkk�*$�
C>nt�����k��u��<~W�|�4��%OXӘ���Xa�"�O��[z�Mo}�)'HU��#{_h��k�h���x�����ʿ\]\䎽����q,�06���]���^��72f�*�0��20##��t��%{�]����!�f��Ճk��]��ߓ�p.U�|�{{{>�2�^�zR������b
t� �"��M���h�6��=�[Yy&Kݒ@j�(4����M����B7�����x��:|FN�Xq���J�B����?����allH9��9H$�7Fk�r��(.���9P)�C����G��h��Mc���� ,'dee}�3p+ ��?���P�eM��O���2;)�@g�`��ȏ:�(�;��E������5�^�����v+�
�ȵ�m/�N���dr;�^�F�b��g2c�B{e<�*"���� �����e�Kk�נ����0)z�9>�����E7N��W�
F_[�1�t�ׯ_�S`�_��3pBF�&QjA��e�_��J~�rA���|^g9��w�ڔ�ݛ�a�2p���y���ٟ{{}������qY�s���lgg���̕_�
��}x¨<�vD�����*	�w��ǩ�8�~u~8�7���K(�Ӿ����E+m����ZZ�;[�2�M,F��g��J�(Z�E�c���ň����t�=x���-���q��1����*�%8\?�{�7@=���$�"7S``�z�r��O��'����� s�zFp'�[��iV"����r��E�Ir�WE�"��
xP�N=}}��D$D(XZ|��@�Rjز���	G��Q����)�1�q��`>��84�V_�
+�u��m�E�R�R�2x�h� ��(o��a�t�%m��(�c\Gt�ʌr�v0�D�~?L�u�^ŰὭ����Ooa��`��-+W�Q�_x�2�<�O�^%xT��=.�~67����C3v �ƚ��ʧFQh��\,`x�r����a���f�K���j$n�� ��̬�`�%�o#7�L�Vjf�)�hM�e���������4a7W�3T����-�h���א����J#��b�׾=�����GEՌNQ��֞�(�Gh$@TA����d4}��ůI'Ckk�)����Y�#��4U�&5
#�����AT�s�vϊǶh��e�6SɃd�c����G&''�n����yj�m�(�1R&�Rq�P����E������l/�jl�"Y�y�F���3�"�1:�j�'��j�R��?j�,_��~L{}��@A*ݛ�a�%�OA��ܘ�H��i*�C[�bؕ�����l̡���nh]��	�N��zq'����"�&h3K�0����� j�Z��xJ��AJ�v�?���QX�Xj#�C$����JKK��4�p�?}R���aY� ��(�e��0���,�8,��:�b٢P��g��2�:N�����z���?rM��:u��3��P/�+J��5JJ����H��Q�2��Gqqq���9�8r��cx��%��iQ�ק�������鞆�F�z%�i�<�Qp�GQu�M�>���{�{��������"���r"��C*�'�p�x�g�N�;Uz�<����}�9�΁�m�In ���f���j�F$�-0nC��z��j<p!&󰆽ZF'��63��7}�0��
��S)=����n!Y��Z�s����
v�k��FXi���/��o-rәNq?s�@�I=�aGϷͭda�u���_� +Hu�������	w���0U:��:!z9��R-���W���Y�z/����z�7�"/�ZR�e�r�
L�=b�t�L�&�&5&��@��&t�$L��eq?�r��t���E�O@�f��_X�f��	��z�����Q�q�Q�L%�o���̀���z�\�T�����0y�*�B�������̚�L��}�9��N@FQq1��6�Y>�[Ww������{��k*�a�M1���^���t���&��-��v ��4�9A�^�9`ى�>�!8�l��h3��`=@:�an	�z@qD܃�Ku���(�>8���y�����8�Ǘ.>~~9HJE�M1�w����_����;mZ,ay�{�0rO��(%'�XM=�En`p��/+�v�$A�9|ۤS�w��H4Q�B��q�8�raL�&#�L���uĦŔ;0
����/�^�����QyB�!"���9��߇\xN��,?�M9��(�oȏ�VF�5ׇ�.|��)֡t�&^p�I~�� R�"e���pH����8˫r���������r������H���]i��7VpA�"�Ks�t������(�dV�I��|D��c*�*R(��F�6���,��P�Ȃa��I���g.>�s �R���k�"ѹ���;�v��{�����j������cSL��ʜf�\���%eێ���p���1�O��QD���*Z���%�\,�4�[�8٫󳪑7.���Z�2�C�t�V�
�)�!��j�1_��ȷy�N3�_��������LL��i���D#�R��b����i�]�#�6�"88 �	�b�<+Ao�	T�����؂�o�������>*��Rc����x���X<�(�0�uX�AQ���:�Nw@�вw=rUۈ��i
��H����V��>�\�~�RŔn1�X3�R��~�v?e��Xm�tl���i��	����/������SPDدQ6ŧatP"�'�4��x�!A�}�G	�;+&=�]Ƅ�y�\fn�}�U�C�I��Y�Y�0I=�X�*����nP������ �{��r���� �2s��Ѐz{s/]����UfM��Ԛ��0+�,���h�������`��:_F��
��> �����#���������iR����'����=є��B�LB]����%�g��ć���3Y%�
zlA����j�㏠shgM�Iq��c`~U����[�(d���W~����^@O~*�$��U�c�\�� ���!Z��ܗ��#/��K}��a�ϝ@��84��aL�ҡ֦^��"���Τ?�R۱�(���9�|Ku�@]Q�zy��ep��7�
9Hua��<����
�WɏJKŨ��T(��0�� '�:��
�Q��;�:�P���i�Ն���c(��o�Z�*3�T6�{a����$/���&���}���S�V�B$é�� ���.`p�yЈi�K,����IA����}^�pcek�t��Ɇ�4��E�@6�.@���� Ef��+82��rw|\P�/��Q���,3�hy�Q��'�˓�%87�}\O"�Z���]U�/��38�f�B�V�H��ϮK�$��[��)��qd�\͠�i�.y�V}*��=�(. O(J,4��У@��`�I�W�T�d����N�l׻��;1� ����Yy�v�S:H���bD�ѣ^`�=I��i���c�=((�E.�3�_�T�avB5��r#��H����ɎyH���v��_g��mQ_|`ݞ���8�5�q��s�msk�oH�xh/}q��[( �O-���Ϣ��By��޻�����8�Ȓ}@�y���j���w�"�7�������ܿ�}Ӝ�.�%xJU��<2���r���|����N�ow~��nOX" �7�=�����������|+���6����/!q��~��S+���H3��	��w7��j����>�JlVMS��8��}��6Ҋ�Z�m�^�Z�m�W�r<��A}�AN'���3� T4)~�NKPyRx�ǧ;8Mm�$t���#�ꫡ5a��
��{u-Yy�y%�:��8:T�Q+a�)���c�<�\���-����࿏6���8tпO?�������f<������g���f�����=����e�W� S)Y���-��l����������%�b�IA��,�G� n0`��Zٓ�	�O�ޠ��F���T�Ce�a$K�%�^������oM�?��z�Y�;��Ow�ٜ:��D�g��˟<_�P��}z(�p٦�t){�ѓ6�Õ�i��>�j����8���٨uZ��+���;����Nμ��-���o>q�����?����u�#���T������[y�N��3�X�*R�c0C�&�y��tp��	�S�}K5c�ZΥLt�3��~1as�g�4Mڦ�.�X�d�$71':=������z�#����:���B����arO V6%b�ڰ�ӿ=f��1'�&d���.�Vt�乣�%/�B�e�b�Jg�Ts����J(C�ǳ(Aul�RǬgQՂ[����[\;Ժ~��N܋֌�ĭօ��N�#��`�ׇ�G�v?u}�V�~����m��_�3�Xd:�x^�! ��f���ٯۈ|���\��i�������'c�LY�ڼ%�������t��(�co��1s�i{or �s՛���\���\ǹܞ��Ѷ���C������5�m�n��������y;��[�%�wy�g~\������1�:[�}ϯ�C�
���}W�m�d]K�r�r7G`�-[ �#T�5��r��+�T�+�$��o���E�������u�
!��3gX�����8��]ժ�`
�L`�Ė�H�R��ǋ'�oȺ����8���4�w��m*�R�RG��%89/t��40<�z�3�%f���2!��m��mH6�YN5����8��'��EC���#�ċ���.��֒�|�r����@[�Ê��#�?[�1]�+3}f�E{�X.��R*³5����
��W:�u_�3�|ТŎ�o��]&�_���}x�%ޑ����"j��G'���Nh���q�W@@z�JDS����{\��Ű���枞Q���5_���P̲&�ͺ*ʲ��W6N�����3���ɗ���;�d�[�%�T��-a�2n��0���ЯCK� ��Q���:⽃�.�f�i�]��f9��>m�)r߲�K����ҝ(Z?\�gdl<vj.?����qΈ���5�A皉D�Vg��4��c��=^XmH�bE���"ThX6��K������߮ﴟh�	|�w��u���#������D��||�k�	�z��5�{ks
��;q�Z�d�M�;J�{r5B%�|��-j3��놠&G�Qj~
7{�>v��d�H���-�%�x��gs!��-F��n����ő�����*���??D~���8���N����$���^��\!q�,=�� ����}D�Ć%R�'luO��!W=|�ԕ�e�iK�	mO�R�����N7t!�5=�O_ę{�Ǒ���뜻u�w<�����]��K�Dee�$r�K�w�s�G$�oJ.�21S�_�8�,����;�&,dt��x�N��-q���~d���s++N,H��N&�%\O1���3\m��X�n���3��D=�Wc�w��gAn��ۿ�s��r�^άyJ�~c��1�rc�ͨ|BV����r����ɺ�i�H�<G0m/0[I�-!�<F�I&Nx�fo\s�7��-?溄�)�K��}��4\�r��t4A��W�V?���H�	l�� A���m��)�3��
�6e�)%��G���u|6�����g2)J��mtZ; a�_!�"]V�:/;K5������m���An)��&21��>��Z촃{���pQ�"S��{��������Mj�HZ�����������Q�A��PPRB�i)�J����z�nIi��Q:���c���眽?�}]x)�g��b�uϲ�]��9�Y��$���v���1����7P�_���`���F7c	+�F���ʾk>���V���"��t�/y�-!�[˹�K�ġ���D�Б��cU�t�V�l�Cz}Sl��1��2��;o�"�p�|����7��{�Z�<֢乯�n��[��Ю�f0����tTğܸ���Q�5D�i�U@�\N(w��;h�
���0�@!��1�~a�B�8ϗp���B%�ت�5<M��5���]��h�D�(Z�`�Ax��P��zck��g��Ci�G�ই��Q �:���?�&�䓶<!�P�����Vb�F!�����x667W'ˠ�ȾH������7��X�ma�^-�#zP����2�Z�lޓ��lbMA�!n�oi#{3����f��6k�D?��_f	`}%�c	L��~sr�lx=P�F���NJ��u|��?�{�W��3���VҽfN-����=;CW*3��^���a+yw�:�\��̹��i��H���6>�!�6Èچ죛��e��M+�7�\�\D��V#DWb2�f>7�����C�#��~؁��p����(�.����SlF�
'F�`^������v�Y�3G�:��m�^��S����Ϩa�y}�0����Lk����k;�`�I����{��&%A��An���:w��^�c6&�\�"(���l֜�|w�l�����!�B<MRP�/�DK<nZa��vx6j�"�������,���v�t�J޹?��۽����@����2b�ҽ[����s1���'s?�+��5d��P�+�Wp�)8J���<�;�����e��xE~����@�&&�M>��B�:l,FU���v�w��}��M>�pd-�����.3#��ejb\�H��Yo/�RY��`�M��t�+��8\u�7h:�+�sh�r�_�1���-��e��j[����A.iB�q`�
}�X��f=Q���Lm���S�p�?���du��/�/:%���-q;�:��ݞM�lV`��T�]�k��Ih��®!�k<e��̷�t��U�[ڸ�È��9�a\�u�#A�݄Z�v	ͧu=A�Z=w~���$�i�H��@* �ӯ:/�~��O���!�?a���w-����69�u��J;>�0�8)�u����Vϟ��(I@o��8S����Ч�&�������3;%��q��^}0φ��f��]�$T��{�o���9/jj��k�())D���_��0� d���۫��p�1�kep�a�D�qZu3�G��и��h3oiE�~_���a�N��
E��������?�[����"q�N҃-�Ӄ����u��:��L��z�s��]U�6�>`�-�@7j:���w
��{>��C9��IHZ�h>�N~I�>�)���ֹ����{dx��*)�:��4A�=�l��"r�4����O��w^��i^)����h�{{�#$Z(�!�5qIkE݉���(.X�����#�*�H�]�堙�hҦi�\ۊ��2(�c��-�<�<�m��GE��҄;c�OBׅo��{�A�c�F���|����E�h'�ɬ�H�5ٙ���_&�)B�Q��j!]Kb��н^('��
��}��& z��o�v�Y�c����R#�ת�̨��F��Bd��{������g����w+�}��*�4���+�b楏��A������*��*�n�f��DRX�Û7oV@�|%�����R./�Vk�v5�=w�
��e�3����^F!"O+��ج�����yN �z���#}��ÓvZ�I�n'�<��T����z �:�Co�r�
R�mD˩&0���IH~��S�����Oޠ6w�re�E��x�D�q����^Z���h�u�8 �Q��[�B'l��F�$(�K����OS#��DV���b�#��!��c��<#|��%�g�c��/wL����(��u]B��q+��_5��Et���t;�,Qz3���t�غ�w��:��ֈ)�K_N2w�I�j�o�)qCg�u�2"�,[m� ���'�7�`��:{53���a��Wm�������f{�҈Av<�i�4	�b��mippG�� �[AF��\���jI��y� ����.��&4�(��ݨ�n�@>8��}��)z��p\���#�k�r������0�Ƴ�-�J�{蘙���m³ȱ˕���$+q�����[�2�i��]�ZO��-l��­���0��wKzԡv���D�����4m��D��V�]�w���)�?Ox����H��y�AY�B�n�#��Ɣ�SJ\O�5������;�������c��c�/�D��(�������8�/�=�c����8&�F̭bn«$^�����͕<f��;N[����I����������{{��dA_I��Г���Zb�=�ݐ-����K�U&G�A��%� ~�D\m�/��,����_��߱���<f�_*جK��~��VR��y	�.B^���&i&v��#W���#N�9ی��MlX��g�13��'��ʬmYxm�yIT��ʢ�a��eǴ�����q�8�~�sLݑ?���B��6~��d^\��;�>D�L�����Kq��@�#"��=溴�����w��:��na�X���)�]+��z�a�j:��]��Q���L��-�%s<�j�a[̓?.>��ò�_i�ѫ����FP��+�+Mn���"��l:�"@���H��q�su��JKBQ3�Ej�A"��OՄc�C�ĝNs���P�,��0	����������lbĠ��0A�V�T7 %�M�%�pK�]��2��z%��!.���������|�g܎��i[��R�~�u�gU>D8y[�C塗WS $�%X+[ѻ� zݮ��(}��s0����Vt�ʡ���q|Y=��������Ev���Ν�#��mF�Wq�� ��quM�M��t{���>V�y̻�ٳ������o��E_Eb����W�ם��0d�ꔒC���i��xeT',�J+��_U>fI���T�����c��%koE��o�aj�-%_q1�8�+�>�f�j�Z��V���0�z�7�sAB�� {���޸��q�ֵ�>�CE��E���o0a,ikɌh`���U�m�3���V�'�M8Z��6�_렏�Г�?Z//��*j�:�z�������i�Ԣ��Q� *��H��|]\'5���#z61����C����	��K����5�¡Ew�y�����Ԋ����=��]��։��e��7a����=��;�7����|��=6E��'��f��ry����Q������1zo��/��a���9���4	(S�ZοJ�K��_�2rom���*|S����?_\�'�{����"Ӵ��'{!P#���h��8W�G�k�r�zMe�>{�_�!���XZ%����.vb%�mb�e�����K�-��,zuJ��+����a�E�jڡ�%�����d����a���%�P�ŨaY7�wdߋVB�F��N��q����+�� ������mѴJXNu�#�U"��tӎf��>������`7V�yq\v��\����'��3sֲ/a���bx�D�A~���Fv��~��Qat$����ɓ8t��p�<�k~e��߯V���;����%�B)��^s=YE^��&���Q\�����9�A�,1R[�{o�l�0|��gK{�����ی�g�T���_`7�sssu��~�*k���1����<�6��9��2=�C����>����f�!�R=es�������2��-�����ׄ�\����������D�=���)���Y���N��Oג�~�����2����9�9�(+.�B�!�V�=Ά[�'m�X2�n� �ռ�EI2,;�Ƿup,z��F��H�*�����ltgR__Oi��ڷy�=�>c�vٚ�ڳ�n�c3uQ�[���^�]Y�����X ���Z��������-��e�bc_t�����k����a�yX(G��XOUhw���/��ǫ��Lu�U��b7�������U.˟֞�}�]a�.�I�7�🟬��p�8��Ǜ�X:�}a"p�e;(v�naj��t�"��w�kH8�pq�?��������krrK��$?X��=�8���6
7f�Q�Z3���
��0A����'�J��ݝZ�U��=倪X�<~��Q!��.���v�j(�H��m��.���߿)ݼWz�?ji&'ӄ����_�����|TW�/�D�8:�]��
8sMȗr�_�'��Z����¼��j[A�p��N����6�D�k��>C$>�mBG����Zr"�^�}�����i���4M̀��+	���Vq==��{߶0�P��������ү߿!��S�ȼ*�\%|�����|����	=c1p_p�ND&�56>�c��}<?oP�[u||��]nbѲ�R9uu
�����,~v��@.��N�������O>/}���N���|�A�_c��Jo�&6A���Ȩʂ(�0 ��DST���&)�/����`z9yy��tX�T4���o`�����/8��Dh�A�nB��cՏÖ����x���*\���B�>!5HR[SC�{j�/�4�k����M������E	BDJ�?�-t̶���@#�mi�=mi짯���4�G
Khw5b��2Yr`��\�JH�^K_�� �P�+z�����ǭ��efe1Y�Y4��A�=,���?���t����9�M��	�t\	�"b��>��ro���a~1��W�on��*keU((.�QS#
Z�]g ���T�W5�Ret�Nh�u�o��ʓ�V���s�������D�ůr�
�2��gVt���9���|��9Xh<n>����*bU�RP�S�q��!�[�D��C����U(���U÷����Ͻ�ELv��z���{��p`����MMt�׬��Z�qj_8к��AX�N���C�A�f+�
b�}�J�n�^�)�SdGގ�����5x�����nf^�F?��i��\R���6���_��ӊȸh���+��·�_���x�A�H&�hV����n�(�/l�ud�)ſ?�� Ȣc��Sj��j��zzz�[����uLѼ��]��)���nd�k<S�ۓ�߻7�3�&���
�VmX6>�-�J�Y��C��ׯξ��M	�����w������zG�Z͋hv~�Pggp���
�{����)*m�9�πp>��� ���Ѿ�׹������K�%�p92���on�L���D�K}�C*����ecÇa.a���ޙ�F���.?�Y\�Y����ĝ����UR�zʗ��d��>8��׻�g�R�-ΒX��l��OW� x몝�U�v~F'a���(p5�*tl�d�x����y��+�ߨ��N"��M��֠���FJd�d�>cv6�VUdnKZ�q�{�X	�LѽB����'�:�����Գ�����S���m,9���C ��f 8�7��0�o�\>���-������ǌ�\�B���a�{%a�۾�a��Թ� �4ek�V]D*�7?LLN>O�^$��s���=�i�u��sJ�����ۖ�7f�J��{�Q��(0�-��n<2��i(eyJ�|q#��.�xy:�Uf����$;�y���O�����m��s�.Ð��y��>���JVcz�3b'����>+fudz8��xD�<:�?��D�@���F�b�����:��s��ݰ�A�+\�f4r�D����������s��%8���s��-Yn>�]��L��E�{�yL�2��GbM����瑃��h�G�~GI�?�  \�ݐM��eVN�

|�0��z@AA����g�(�DQ���9������cc�F�Z�Ω�)NK�)�E@E/ha�
��k��#��?�D_B.g�O��Ij��WwOJ��@�|7d��S���}U���Q7tt�����C��T�A�*�ۋ��}a��:�2	�i4�v+��Տx�V�T�3�#e�	�εi�����q�ړ���z�����\��nS`�v�㠤�D�������Ų�-x�w��N�lA�������|K�������<��;����W5���`��}�������s�qf2eeecGGҴ�4a�B`�o<X	 9�(<�����X�un��l�e�gs��wu��>��J5�����\%��w�J����`���T�MhM������w�gff���ni�MOw��N���rȃ�������]�n�U �K4��<HT�=��#���(����ebb���:_�G!#��n���X�)=#cg�4M�$�?��w��ڄ�����x�ܷ���	��cvV7.��G��K��F��r��-,����]�XYY���RV���tc��0�K{u��������-B�A�ju���x�3쩲���GY�����d�]��:|���sWCv��S�TѮ�+ dzzyc�&x٣�7�*��YӺW�I���h\t�&%� R~�}6���B/c�}� `�����4���?E�54zc�r^�����j����l�:D��S�� �pg�m�Ǐc�=:���y���O%�NT��SS��X�ˁ�RRQ�j�m�}��|�3����Zٛ��Hy������"|4F� 5I��֦-�Ť�6M�6p����>��6� �B<Bm�b	��k�U������P�x(���L\\(���n��2�+a�F���
�mi�۳��]J	7����as����Jh�5UyPhZޘV�?�= @8�G��3�yJ����ذYD~�:����>��2�|�V����5�;~m��z=z�jQ�܋��6_�!d��~�c�:::�؞����y���\;�ֆ�UfM.m�p2��T�I�����w���&������3����b�ى�����R��y��v8�>^�+��۶$bG8-�w&(���2���:��;� Z|�>}��'��pp��
`�%--و�E�'%QS>~����&���M���! ߳~+,<�2�+�K��4��@VR�h�s���_���'b��|� ��Ϡ`�����|�z���hd*)�����aC� ���mJDӊ�===+�g���[&.��OU%ߎs{d�)�}���-������8�����?lz�%��D�A�`��`�XT���O���{�BAQQ�L��j������mfFۤ��3�p����w��B��fL�|�9���
?���K$h�H���x�eT�b�� F�FEE�B���<e`�sw�`H�8/�a�z���m���5|�ry�JLKϰ��nq�\�o�a�+�4�7sqvj�����w����FB@ �?1��!6NG��C@W����+�|�����N��"��e�A�������=F*c]�o]sZ�4���-b�1��4��,@Yz�v+��׌�����ү	~��L7�x-F���2�䦨� ����� Vf��t8_��Y88p�����1�t�8���"Ъ�m�em`��ڹ�x������Ռu9h�UCم/ꍘ��Ϊ[h���V���3��mYs ����t�Q[�����N	��H!Y�wM���U�+͚ &`��3�^ž5�y�!�!��lC��Y��בm���V+C%)��*��ͩ��������l��n< �^	Y	���~�|d�^_�VYE��.��R��\�B��B�Þ���?�l�<�Zn��\�E�@Zt?��6��
{��~��to,7NM�~
ȳj (�x�0OOO�"{o[A������H�M��
���m׭������W~�[]3�<q^���ZDD�h�;�/�F)v>�.����h��"�SB��@�@�$i�\�u����qg��k>>rX�ĺSVa!����r5�]�=Nv������s���\��R��%E���� �D֖ȫwrD�e��J���nB����E�TN�w���5��Q?�|���z�/��������P*�7BF,�A�u�,��wS�o�_@�t���E ZZ_Omy?������4p�zUx����fǆ�m��%#���6f>9�B2=|X�Y�MKn\ ����P�����Ƽ�==r�FT���~�*l�l������`h/�/_�6~�w5σgي���WM$���.}����H�b}����mR����m�,��E��f�6X���|��[��k�	W370=����(���`�tX���3@Հ~=�NII�0��� ʤ��ɝ���v���R���}�=a5�$O[�NՖ4�����؛�+l&_�j�:5!O���OGgf����B��Ê�lj'g�/�%�/ĪG��� �D�:�(�U h�dǌ�)�ix��{��C��ͩ`'�p8l�
2�"��BK �T(�|����*3{b���"3���?ggg�|�I}����䫊����u�4#�)�/~"3�48b@��.�NJ�7f8�k���ܶ�
#昱�b��u�h4�r�^^��I?�gSӎX��=uu���tm��i��/v�Ps_NU��o�Ke��S�|�6�4&˄&nmoWl��,��=���kB��8c��1���6�6�y��2��~�_��̏	��x�+*j��\�L���¢'�B���-��w7���8��v���
w#<�
YNЄ.3��f\�K]	P<�7���ϑ⁴u��4�5��^of�,29�=���T�}55_R�=��av �F� D�w�����8кh��`����؉��5�eX)��ͬ0v(;��#�����c�C��-��{�xR
�H���k(|Fnjc�w��;������Ņۼۮ�ʛdmtMKIn\�(���;��6�)l��Z��L[��zl�x����� 1:v_ |�]3-hY��){Dw�Sϸ�<�큚���t��M���lKE������5Y�+��v�uTb��I.^���0�_��bWztjҀq���N,Ֆ�PFmڂ��֡� ��3`26���k���R��?�Jn&==x����L��b����.�ݲ^#ԤAA�VG��N��\
�+itcc��\m?�&66�+����������N�b~ʕ>�j�L��@Vs�
�S��WDTT�ɡ�Vw�2�}!�6��T$n��b9��?�7{ ɀ�}?Q�
�$�*������LE �����?���G]���$�'�yҖ���WQS#k9M;l�w{T�#��ˋFZZ:�����P�$��C]�Q:��
�`yy|����(#����s�s��}�(�/���0(���LF�Ջ���b�h�+.�eok�]\�]}��c�DF��Ur����L����"�����+.&$��z��H<�Pa�}G��gb"�b�%�f��#2�=�"�d|�3��aκ��U�:|Ř�j�h"�c���Ғ���'ZH���y�˅���+4��X�z�_=�X:v�:���׿|�O�q����&�����F�A_�PR.a�&j�(��A����.?��&���[;�-�ڹ/�*B��:� ����%�.���EX,�l����]惏xƘW����s/1��Qŭ��� �G�sE��m�BZ���>xD�ś� u6������|������.\���s�l�9/���T�����c�o=~hʂ�yj���V��U�jݪ���d@�4˛�t�y��qqqaMmĠo�"��Е�g為�vfCg�}��=0A�1CF0Թ�٨�=��E�C77��Y�2�p9.����ُ::OA��^���a�z�R�(�B������s�Z<�\\�?l��'�}���}P�ψ��;��ի�%�m�Q���b�������+m<h��h04v�5qW"�Mt3#d��k�����VQ���C�C���p��r!���!O3��p���0]�v^�q���ݳJ��`�ط	�r��^��6.�����.�}tw�4�Y��}��̆7�?�5ޥ���!�aC�mhH��df��φ{���{׹�#�����ռ��-~�L�I�_��B�l��R�]�����t�@� }~�Uv�� )a����oM�j�P���s.�����^@�b�f^�I��͞�{��T�ik�i��`�؅cC#*0���KUӛ��Z�hVԮ���������b��7x�݃AZ{8��uˁ��C .����y���ye�烒�O���f�wx���r;>#�G2p(ej�\__'�%i;Tu���{�������(*���*�-������"�Y�H�������� ;bs����6\�W{�0��L�Os���b%�'f5�}��gu�����Lll�p;/��L������_�z��	U�j��֟�hˤBY��v���zVr��%�}n|8��Ҩ�>H�L�g����n�X���+��)_��S~�����߂���!6�^�q�+�Plz1T�	���
��Y~��H�QSS�cj���\���#��� ?�-|_��{&6��`Á<��"�뛺M�<���b�)͋�u�����\~�N�f:���a�임��Ą)9�?�nt?��D�˨�	jJ�6Ͽ�RH\\�rK$�=!v�n0YS�{�0�Jj�O�"&���0�~���ӯ�l�CL)[a�g�����,�p5�ә��^^��E� ����Ιæ$�@=c묘'�4ika����T�o�̌������[#@�]5�s��$�!�=M���fV����T���Q�ئ�W�ܹ���狰eض�H�-��w^)��D6ꇈΗq?	���ee1-o(yz��^BIb����#�_�2��T:��Ԫ;��K��zɕ�;uxH�'��:rNUij�����"�e\���wf�Ó���y��k<8�ɬ������p�!_��St;n��UG�����Ӈ���A,&)q�Ra��b�l�2�!�Y�#`��/��⾸�r�'��3�x�r�����H��)- īE��ؙ��<����LO�ۡ�2KJ��s���0ޟ�>^��B�1/�$p]��A1��n��M�(~lHu���?z�s���p9�eJ�3�t�`��n<� Q$访$�m~
`���)))�W{?珇D�����}/�W����|C�C.����VYY٫K	��� bz���~J9[Q���R�GmMMǶKO$��\K#6�y��W���+����Ҩ�>���ڔR��S����wUz��=PK�D`ve%9 ,�3�%��R���tL}����;�sp�spp@����V�>��M�G�����UY�` ۨih�f���JCC��١KV�J��f����@��5,~i\sJ��i����O�Wq��/�P"9`��pq�������� �+�W�-_;;�o#�g<���/g�4Tç�_�
�*��;."^�J�߱�����AZ2�=����WoOK�1K�k�/���o[��>�g�ڟ��ي}g>]��}��$��ud�>^��ު��p�M?*;��Y�|�軐���<�� �1F��B�џ�ѳ�²����r���G� ]��*HM]x5KM�h�ZM��mᥲ


Ⱥ�
2�ī�F��ws>"	�ˤ��h�ܣ!�}���V2'rwE�����]w��vyJw�.�k���I%�Ǒ,�aB�!�
�?彼�,d�2�~@�]��1�;d.�gO`��D�I��ĕ�4�L�,9՗>���9����\�N�&��h=�<> ��\����ޗ*4��MB����>Ϥ��XZzfa�m��C>V��+uM��!&��������
�����y��A�o�~������A,@r���KJJ���t9�2+�tbƒ\����%�pq'�"��^1�~PUe!_.�Xq]8�� ��� �>5e�;U���Y����̈́�TҌ;8��!؁s�G"jٳ�`,���"�'#"��B4��;n����Q!��{}d�7�_3�;a��&��3+�����ʈS{N�hϒu���d������H4�:;�<�3�g�ѯ�Sn9>t�,r�Ӌ�}!V}l~���x[ś�w�,�!KWǫR�VUZ1Q��ײ�`C�����?H��*�;
xF.�P��[R��Հ��fMKKc�E$�iሄ�5m�ޙMDD�F���� 
 u|d\BBNe%�����N����m�i��;��]ۈ��g ��[V6|&��]	����$�>,W@���z �-�M���Hi����o�2�Ű*dloo���$�}�����Ҍ�4=��E�҇,�m�}�@�w���s4��_	Y��&ؓ��:|�g#���M����}#�u*1�rP3�t#�n{}$KZ
BsQ��������$��u�ܤ�r�O�oA�go�R�ckZ�8�ଚ Pd��&ओ�����rm�k	qت[���;V�q���u�����7ge��-q�6������'bo�K�}6��1�ED���^�Ukv\O_?�r�
b��C�O&�
�S�W�dC3�(�{{yMצs��y�0 ��-4����(g��E�D�*&6-1���d����H<�67 pfm�W�._��d?��h2�=1#m0]İ)��֦�tu�[:���� 7mr�w�9��﬈�����怆�).��OL|���y�j�|��?6b�.	�-s'�-Y<<��	�մ_�Ud^��mE����i�#�RWg1���y��l_�حlh?��F�$'cϊl�FC�Q��]�b���Ғ�L�(l2bW�&�Q���=lb�X�_��`o7&-*J���rPnٯ��s}R�hr{�'i�SUs�[5M�|����(��.��6kg��;P�gd^�`�Qat��c�H�Vxr����(��N�r�����)��3��-V����
;T)�{#追bf������n9�!+�jZ�\�B�y;���22A��'�{�|�*��������6QTr"��]H=@���(0�����6U3n����?ޗ#߁Iw4��V �#�P� ����O}y�ԍs
��w덄4�ձ�[�'���DJ��i*~}��{a�b�z��T�jq�0k����ݡ�QI�{��V���kf���R?���M�%���1�xx*�Qg?߂������܍��~hb��� �5R�c˪��VF*��|��#��Nf�@|FFFy��"]��~�({��sz]��>��?دbٟ{�<��"6���')�P����K�����EE$AQp��P�x�����\�d�&��v�!��g�m_=A��F/]�7�����W#e~�9�ҽ�����[�J1A[z�� �������T���f���I�ܗ��j��k�Z$`!K����]
7q�ۜ�?��Ԥ7��_Eyߠ�ߍ�/4��	i�4��"Nym��u��W�d7����$7��m�l@�B��~��?Q��ؼ�g�վ�e�V�׷o�"]�܆BJ�ǰ�W����4<���'��o	o����q#�8���55��������fϻ'���j@MSn|R���K�[���&��hh��f�f���զ���4��LՊh_
.����w?o�9�w �#�j��&�Sx�1�BKw;������f:�w2�=mi�Z�޷���q��B_uG�I�T���=� �Ζ�������Ξ��``���l�-ED-Q�~�%;H����
aJ��4d�	Rp��^,�un#e0�Ve�E��z�A�x�q�z**��߿����a߾�p�r`o�n~�U��<?�7�[,(x��_���Zq����F�I��Or?+t~�����u�|l��'��O#�F9~'kg��C,�ꋼ<��0��_/�g��T���rmE�]qKGdI}/E�ϧ���H��G������Pm�kk�"�����kO�ߔ��
c�`0�
ȟ"�0�ͨ�961���hV_}.�$������^�c����C,��� 2����[������5�M���6�%��%N��$%q%��$��� �qܛ~�%h�$��iq�TVV��Ɉp�$�����Jr%C[�*���Ύ����oe��{�ju#s�s�bSs��.�c��A�B�e��~��.�UCSs�l{<�l��:ӚR��X�ԩ� ��H�k^��c"�����[^��7�N��+=0�OÓ�I�f;qkn`�K_��,+���u��󊉅mo[�b�j �����f� ��B��N�}���� ��q�kc�bbcc3[Z�o����30sS����
��)��K��U��g�c~兓9��o25\:��������tp�2����**)��?~M�-q�9�b�:��5�hat��
�P����9�SSe<=��m-�?��)>��Ȉ���e�t����ذ�c�{��>;�g����.ѯQ�E����yZ�f��]g�
B|��9H��L��o�π�&C����bb��߃��������6�R6r>77Ǥ0s�F�&\J�R���$6���Z����\)���d�aC��ӑ�P҇(���7s����T
0!��4%s'`5<�~����/��/�v)�3/�����=?�ۛ�Q��dm�74�`���㹎_C�J�h_�WW\�������wdj�EAv7��!}Q{�����'Y�{Z�����{��_��JN^>�8=���:�8���/��vIdp`l�$>�!^z�ط���D�6��Lo��3?�@���������ׁ�����X�K'dI���!z@��vAF]w�#abk�\u'K	����^vkMX6{>Lȕ�x2;c�	F�Qō\��]�f4�*S���cjz��b��kɖ�C������ϼ�o����� 
 -1c����B�0� �yW;��wJIp�@@^��J&!3Ǟ�0{��������]}ơ���64���kD^�^/���d�fߟ�-T��x����Kw�1=�'b:�;��弼�i�.�>�l�/K+�����-md�2����ڱ��M�p�p��^d�!���T�SPP�2EmR�|6�,�p˳��Z��������d�E;�k�u��1b�!v{�ʷsJ2. �VvώR����V�>��5$�4��e�FY�׍o*�� ..0��>yw�f�dr6�DZH�DҬl ���re�7�*^�W�P��᱆Z6�� %�J��-� $���;�K���:�����������iy�\�V������{]����-$�֋U%�b�aU�q�B��UU�A$��]2T223Xg���8Zr8BhڮfI���HQAO�s�8�YS�^P���<��Ԑ��=���6´T>�X��w ��Yϭ|��:E����|��YV��3 � ��5l`O�`�k1�����@��g���h�~M"�� }_%�n<ܸ��C���+p ���+�S�{K%���*4�466V�{�}y�n��\I	��|����Q��(��X��+�����������A��D��n~^�����2��ǀ���O�W������^]��=���2�Hp!~�6Wm�p�I�}�<~���s�S/o�c�	�=��f�KS��Դ.�����%���5&���&�6�hѬY����?�+���#㚝+��qd�n�'��< �#���d�e{M�2/�Kj���ဦ�-�9�q����7���55᪝7�ebuq���{���P�ұ�{rrB[ 4�
���w5;��="���e��ݹ�ɰ�!��e����=7��� ;P��/dk �i[[c�6�Т�.��w�Dtz�A
������C�����)�B�,QNNOV�*k<�t���eQ��DO#���*���;�Z-f%e�i�%������9Q�g�ٞ ��6aߕ���Ybkt?���v�������Rw��>��jQ�%n9Y�{t����7���M�YM����6՞H!��`�^��n�/:�w��J=��kr�K���|�~aj*�(�ۃ�<�EE��*�!l�+]k��Y�Տ����C�K-�vZ���uu�Z�s>�����ۗ���K��lO8-���Մ��jX�4Q��c�hAw�:%�+dV5s��f
D�����F��fΎ=?W��sÍ�T�q����g�z_5ha;��K��>N�p+"xǄs�b�Ҿ[� #]Yxӭqtt�	(T����jj�ep��Y��JNiM�NoWm�6��n�i��XY���봭{=��8�w��s-D�O7����I�"x����^4�VM]��L`����R�444�o�R�; I��+;}S�JN�P��	��?���.(,�<�.x�'�S���N�A�0�S�+��T���A�`6�m奻��o��pՁ��&���ٿ�q<�7�O(�)���.Ѫ��JQ��B����S]�mlLC[�A��3$��(�6�Mx���ӛ�����O��A}��y��ރ��wP�,[ܯOb��j���h�E\6���Rp٦ �n�=��=_��6�tv柝�S32�x�F咊sV��S;u�.!�5��S* �A��v������Qԕ��mq�K���6y(�df��Top��-U���UI[�3�u�9jaaa�vv�����rÐ���\\��������CdI��N�7��k��on��3���;³�����7���]|C�����2��P�,U����_�����:���͵h�֖��G\� �ֻ��i�EEX9��3������TT�䮬���w𝔹++I��_dd�, ��Ȅ]��t�@�>b}��iVE���Ń�Σk�c����۷���W@�X98`�e�C�c��gH��P�����j�l��ν���'E�loo���'��D�J^^��_�2��TYii<=}���y;�+�B4�Wi7�k���@0U��b�Ҡ�ᯝ�g�������S�6N0�J��o �r�TE�m���=��殑�e���zݏ�wS�Pk�G�n)����D�a�����-��꾷a��A�E��SB�FR⡻;�K@@:�S�FZ��C��w���oƑqn<�9k�uŎu*�.��+�����I]�YXX���7�s���qt����$������E'd�ۯ6'�+d����u���E���?s3|�Nslg�Ư���,o����{dWk��k�Lu���7��555�Y��Q��(�P�xtB�Ռ�9�������
�(�S�{X��>O���?��(���86<�]��*`9���G��Y���1(�}k���=�;�ׯwo���`@��g��������QW1������ug?C	q��*A*�����Z�ۻ�mfo_���̀�R9�,���Zvi�W��H��;���zr�P����CG E��=����Ǫ���qlt�
%u��V���ޣ��̋X#vK�\e�s��Ж�fT�%����T!�m���\<��N^�;���0ҭS�R4����,,-��U�m�ڟ���ř�e�̷������属-��PR���c>]Y]��6T�lVM*����՜s�ʊP3�Hg (����8�b�ҥt��%u7,D�V{%#����sk���jP��ݫ�Z���ߜt%k�Y>ZukIqu�S�-.EiY��d333��<1�mlk#��V��P�s�PqFD4����`�A��t��9=`�^��SV�Z]m���d|������@�!���ڛ3�ۧ��؍�[[Tbbb��@��~A����3d���-6�[?N���gpX��L���MK#6��+�.���ɉ�9�+J��ۛC?8�_-�\�޴�%)-�S�����cc������j�m�,Z���C��`�7��Lv(.x��FpQ4L�(�n'gg��{���r���8
�`*>>�9C��/gj�:|fQQQ�7{3e���g#i8�e��|�����U�p��]�X��~A�Ni�a�%��#l����f��;>6�ɡG��7\�ʾ��p�8Tc�j����ݨ�����O|&��.:U�}��Hu���ܷ��lnY��Q3i��ɠ���!Q���Ekǐ�z�ذ`
K�W*�j׍}7�B�����{�/��r�`�W�3����,?yN��8^����'�]����=��ֆ֫�R�֮}V�""�>�������Ņy��lᒽ��k�/X@2Ì�Oh�MT�8Y��Ʊ`&��0��]���v�S�D�J7*ӿUZ�U������"k�Xސ�lSE��ܪ�/��R�y���RSX<n��05?k`��v�r�P_��F*�D^**,Ċ�J�Ɯ;��{�5����W�;��_#|+߁�K�~��l����+0&EMO�s	��U~�ӑ�g��T[��eϬ˗�^y{��^�k���S��n�@RM��UP��-3@��:�L�z���rtu�A�R$j�- &	�s*���Ɋ��&п��88@nǩ���8n���}B�n�9�?//�ܕ���h�����o��ϡ��!3��Î�]���艌�oܑbA���c����"�Z8
��+)aRŇ飯�>�q���o�C����k9�I/&m�/-��o��'���~m^�;��}󗂔�)�#S� g�+
�ȵ�="�*RzA���^����JF�i0�B�m�C���������8ϖ%Bs�dQ��ؔ��(u�|Iy��OO�,�s���|���E2$]]��ي�V� ���姞+!��r�ͽ��7J�'/�;`+�����2�EMH�uU+��o��T��<B��m:R-������*.���K>־4Q������N���	II�@vT-��Ny�#�m��O�g��558	�Y(�8��3権�8��u �ѧ�:�#]��v��AGgy�Y�500@������А<�A���i�̸�aǷ��9�U�CujYhU�sn��C-r}��תj �BBB���x�!`���B1|֌�W�_�ް�M���z�Z�f�&�z"��k�矼UU��!��`p72�w1e��+E<�j��# ��Ny�B���+�Y�Q�]~@�������� L	���y��2�;Ǧ�CD��g#��ӨV.�L ��*%5�C{Z1��CUE���� )���V�߆5gD��tTF�RMaiupO��L�8�*�Ə�(�Bݴ,Q&���(ny�1|ձ\N����.��Y��A),=-�z-�Į�E�pPl,���jY[[<}���¼ee#���
\�_�z���\:P���`
��r}jVV�J���{ը�]=��CA�I��M��ll���?��	�@�P[]����16~~شM�#I��А:��o��,)44�r�KWp��痵}� ���w>@w�U��d��_�}rr2J����;?�V�KQ�7�����h��kRz�	y�IҔ�)����0:rK�>�O��:�UQ�>pkɉ�]?^�%���%r�\ԋW�9���Z�w�0����*�@������8u��c"���H-�c�����I�)��bb����xl���\G�B�e��v:+�2�!B�''X(�Up_�nf���R|+��QP@��4������� ��vɼc��rkq�;��b}�b���?�~�{�Ԅ���R�!%I_3w����o�%ɶ��/45G�,�c�M��D&�,:&�s�읩)<P�&&&�h�/A����i8����g���������VH ��k��B:�1 �����������IN��k�E5���c�H��q۷����4�V��VU���ч�����q@H���T��y�������q�5��-��cN/`w�=��7!t�|s�4����=�L��t�o�����%{,����n����\`>@w9f:\Tȅ®��<�|>����O�rJ/��Wk�j�������s�7�JJJ_�^������yK���	�[�����w7$��1,-Բ]��j�ͤ�����rZZHD��\,-���:�����deb��\�?Ivh��� ʄ��hH�36��S]��$�e?ػ�i��|��7yY�Ka����t���;Z3�k�q݂��k���Ύ��WH@;^�1�{~�4��"�Y���Y.��@Bf��[��������O��� �F}:�F��W���$1��W/nօf��	a�L���8�,_�����Z��~]����Ibh�^��}q5�S�P|�{_�K����ll}d�K�P�~�[�XR� �"�T�)�#���IZ_�G��a))a�]��Z?JY�s�/1��S�D�����#���T /(��ZgY;�Z �w+����K���u[��_׼�5�ꩬ��tx�������o�l�/Wƿ%��Uʓ�Sh�
��OJJʓ���4��O:��0 ����	�GN� �EPl�ywV�ɳ$�u��k��M?r��Dd�+�����se�fQ�~��:#�[��M~<h���I���>����R5��~|a!����i�q��Kc�&Q ��#*\��:�(s�^��M�E�������}\�f�š��DR � -"��r��ޙ��6�9�'�Z���!��r��ɠJ�uޏ#�!n^޼ϟ��]���D!.E�����P���;���A���i�R�B[\Y�&+$lx��n�tS:���g��i39��V�;�����+X��۷���l��򟪻}�Ԥ��^S)}���6K��s%gZ"��\���� �ﴁ<�%�*�"�"E$��~e<��x&�o�����N`�CXj�߰��;>A�+�ҵ���+k�ɜ�>)���6�t�9Kf��Z���9vh�tP\ZZ8C����W���ϣ߮^N�ec^mz>�W�ۓ#t{֕w���^^�<<4͵��%�����)�G�=ɀ���g7j��K��Y	�~���չ����J�:�=`j0����a���۸�̈"�L
�3��
Nxx�@��Ij�=O�766�YG���	��(�"`��&|jJ���I�,	��,8DEc��*�23��Q
������p�������~��Z���r坴��:��s��N��KL�F�3m������]!��.���"��'��[%��*t����(.MSm����g�XC&��#�^�	DT��#��v�Cy��@� �n�Iސѯ,5�I�-���� L�KL\1�!���/�� �x��%}A	�	��������M]�|��Jz�,�=��ߵ�-˱����ZZ@���Κ��tQr�Qq�7��fWy%Q�+W�ik%����e���}qس_��0h�z�J)�Y�DcՎk��{���Yf��u���wՄKvV	��'C�DD���0�dGu��޾3����\��{~���o��D�4%��|�(���[��DP�|y���q|�g�UD�b淛�T��|�-	0�7i��9W �_:}:u~���g���Do��Ѽ/_��y"�I��E�(�`�~ m�����TTU����S�Y�\L�	���x�T��4�U�)!��B&�ֱ�WT�Y%A�#L������o�`�^�mf���f�9�y'�o�8�����!��������JEpC?}N����o6(���!����	3��vd��N�O�����EQ��4�[U<К���<4�7$��4Xj����֪��|2=-P�h̙(42��'J��q:;:v8���s��sW���&�ۙ|�!�;�����F�{Y��B\��K��}�'�2��5S�ߵ���&��ЩbyyT�
Pl����jSd�s����@�xq//]q����q��ɨsIձ�R�3�Ur4D�*���&��4�x�!~׽�;���KK������\ �񤢢���.t�r4�W��b�;r�w�CI))���ؠ��t8�+O>��f�T�F������䚫c�j�D���TM�q�A<�Z�w�>r�2NA����|�Q�3P �걆0�T!�`z��о�9`f:idU��9U�Kף�	�q3*|I���I���n�F����xC�/���7Y}C�/�R�j������v�5x6ǲ���s%���Q@<��I�J|Ս��#����'�g >��66�4������7i2O�Zae7.n�Sĵ�SR�[P�yc&Cɽ��[A��PJ%W ߽�0���bM�]C�CP0D$P捂��R�s�P�`ww7!9y�[{4�����g��GҕI�Ʒ}��UUW��Ҽ��A���|�Ǻ~Xh9ݩ�<��;&�	��/��z�/<�56�&��M�5����Z&^ӒٵW�]9���8���:���l"�e��F#�+'0�u$.�j�A��o.0��$>lQf8�����43~��g�� �sѣl�XsflX�챢�8����rl�we��c D{�������j����͗\3�Ӕ�(#����������VS�u*���8S �yq����hQ�r�
 b_��"�����8C�K�%{�J������X�����+nv��*�r"@Ct<\(H�h4�۪�3�f����Q�i>�݈����>��ʳ���逸��Oן�7w(;�?������10jV>�-���[�X"'%}?�R�Bۈ��~��H�/��{���Ó�!B5/"n[[P7���	� )��ޥ����qG��/<:�4ssJ\dx\�֌��ܝ[�ve��?���r+,Q8�O�L~�����-�Sg3礥���?&&�r'ڪH��,P�H_�����.^_Ù���R����Rz[�4������м�a�A�l��<�ܮ��^��ܕ���[��=0@�v$###rl�[�:z�<��%q�e�ܚ�*������QB�UCA��٤_ثl��]]XHk�Ҧ#��Cpv�le\�l�kׅ����䡼������z��OS_����_S�k�&`Thl5����+���m���Dsh�69o㲤�F�ӳN*�k��JCC3��"�Ðe�i�N�w��,�����4h��j�V6iқ����=���P�Y�R^>*o�C�A�+EE�i���]��qJ<12/�5�d^�2��E�/q��qzܗZZ�Bs=��g�r��a�S�%�$t&�dd�WVↇ� h�����2
>,��������k7̴����(~�
jOn˫�m:=�B��swu�H��Iނ�J��Gqd8^~@����,A�����ڍp�=Wx�С_5���	pB�Ȉ4p[���[�s�	���_��\Y����m�������(�v� &�[tKN�=���]C��U	r�UKl���o)�8z��������B4�eЩ��6��F3T����	 �n�~wN#�%w��}��g=W9���s)8C-�sM��t��n =L'��[`Ʊ�i�"�#onn6��&��G*�!~:�]`<99���]�m��}\4ĉ�Ũ�[��mEs��\Cdz-n�A���4
�DcNH�f̣;%��P�lT��c1����5��D�z�;��i��~�[�&222����ɾT��AcMAժԓpt<�ӊܞOM�1W�l'i3P�5�8�8
HZ6�¸��}+�FI�h��&J<N'�(|��u9F(��S";�r��!o8e*l���BzҪ������x�Z&�f'���2�-l�zk��+��25�t>��Szzz�����@�����Sd�����ܓ���I�����W�@��n˝
%Xl�.}�"s���p��'���e�����,�C����H*N.��Ag4|-: w"�Q̰��#�R �4�47�|Y
����E+3�����BЬ�637׽~L�۾`c��Q�Y��H4t���Bĺ�:B
�㤈��2��=��Xw��SSp��3�Ҷ�g�E5}�k�&:�����e%%�?[��t'Ё��nVۯ�^��.lHc��T13vrv~Vj���.p�&th3�aԱ��$�Edu"b������ޝ$	\�n_l4���V���v�z�|�8�X��=�4b�N��ZN�� �@=�P�콅���U ���krss��cqo66L������N��8MmiV���g+d��F>Գ��w����eJ]ޛ);����ck�|�f��������ff�C~��t��m�d��Z�^RES,M�}�GGq��N����/Q�?��x���*��Y1Ǩ|����b��Bn�fC}���X\�n����f����46�Bz���u���5��u�U������5�^k�� ��D�kvi��X����>#�\�x�T��a��IS�~D�V+�W����闢�"y����tt��;DT�x�ޞ7%��X9�+e[��%<�M<-ԏ����`FqY�߯��a+++܊u���їz�ys�/b4���T޾��"`c�e}�uǧV6S�'1.$i浴�T�:"��G���� ˁo��f��F���Z��F��>�&���E�n !�� $�p��p�5��*����7���s9R2��֗BP �ց!��a���j��YLi^/�.c�:>J�.Hل����W~~����	1�
�=I6�q�;|�+��ᯜ�c��>�>�{�RR�Q�gM�ީQ!�C���gTe%�������֎3�e���  u�]�0��얊�o^~�x���_�T�5�+�g
¾M�_�~��q��Od��UhF�Y��	�˔m�fJBI��}�ۈ��� XZar@�8�E�xR�SW���=����u&����ju�ww�rJ�N-D�[L�CJJطo�)y��#� ;^��W� eSM�oo?�V 9���,U�@@�N��-��^��g%I�?p{�� "���?�%7�-��6�b@�5 ��A �.sa��8Զ*�Ȅ������5�E����<�$|�x�P#]5b�����jM�/T8~�����9���}xx(C�+����)��6���XyE�ZadA	[9�e�'�7s�Ʉ�R�I_,�Cʇ��2jj�y�J3�}Ts'�,-w���4$�R����	�d�ۗ�W�����`?0�.X����J�{(��W�GZTdd���	�씐�R�'�A�r���{~.Ãega :G�����[EQf�V�|=���P���6��Bf||�����MSI�����e/_�������&m�di����7.��n��TԚ\D��i$@�D<2i����h,9r�"�ꦖ��t!��x�#��s33 Uh�`rj���T�i��}���Ԓ5.��6o�����H:�R���@�?�G>H�W��}q�|��w��w���t���y���|xV���9�I��,- �*'���ݎ',W*�?O� .�Di������@Mv9����7�%����laa�EA,UAZ���Hc�9"F#<8(��d�	mل�㻵pǈ�������T��Nm�����@$��j$@��!��>b����55�[%����Xq�bk)�Э�gԸ�#N�s��,���f$ԒS3Ԟ.}�7��k>__N$����U�貁�.�ׅ�b�Ap��.g�B�|w勋�?��ϾD
��HWz1��,�{vh(�l��ۦ\Y0f��ݐJe[�������� ����/!�V�Rg&������I� l��ի�߀�	�8a"�p�iJQ�3���&�f}�9V�)+G}!�����#����������:ؑ϶P�Qۍ)�F=H<iy���(�mF Dm�/�Ό��`
9wLf�+��c����Tjp�};��e�-P.-��[���)�r��T�͝�}�����I�j�-��u���k�����K���D����{�eUU�:���%@s�=[qH�����k�}}�T�m��iQWS�� =O����o55��E /���7uhR�
��� �,g�8����8�_������,�k	m2Ҵ�KY�Z8��	�2"��'�%fw�)x����_��V����W����^it\"�+���zB���������п���0r���J��C�*�Ғ�@3IQJ����@פ�_���O�j��b&D�)� �y�"�qŃ�jRb�י����RFBy�܄⃨b5I�p��������104�C�����������C��i�hUG����qP�5�"iq?
1o)��N�$�,�����ll��%�hfq��Ue �Cf��pFӒ#<<|�q�Ă<�����$Y�=�<-&�����5�Q������\�}O��e�7`n���#t�XR&#���T��Á���J�����C�ex5�����ZZd%�-��gZ�!'''4��#������95{�lN�9�a��٭f'�/L�-7~��[������FHV��|�������f2�܅m"�d�&=�MSV���`\����͗u%h��^q\�����دξ�װ�(y���[_�9����{��1�I���`�a;;�McsK''l��W�kX7 `�r�V➞>WA��)�If<��>�iii����2�4U�e��H��1��-צ��Wu^^�<�1<���1�	b��۬O��6�l�}�>OX��X�x���/�^>��<#�E����^�����꽻��{_�3�H^�Yn ,�6~�g^����sU)>�%�J

�3�GGG}3eZ*����`���(�o�U���������Ē{q���<���j�f��F�M����i�Ҳ2�eU����]\$S#�6�/�L�||HA�V�d�C�K��i�q��m�Ad��^ѹf�tEIsy��4I��	Í����+�_QCt�I�>:��!ꫛ�7�rs㵖��(3�sku�z�[ww�%;�7�� �O|_��9�թ8�×�����a�d�-ll�]Ї*2�U��>��HS��%I�UF.R����w�4u!.���!�?J�-~�C'��K�gaa�O�����߿���T@*ּ����0k����rRt8!�\v�x�3��<�_�]�@~��V_MMM�(+�����|���t65�.{��-#cԤ��ν+��(��|:�j3_+���@8$܊x��)n�:ʦ���2 ��233�}}}�e#׷�ԧO~���R3윔��#Fy�4�GU04`��NMo�� ��;��'�i6�|d:�����r���$�_X�A�)�4*��8Runl�܆e�����*&G鋣����C����0�S�ʪ�U�	�9���K����r��O}^M�j�U
*�RÍO[q�/H6��
]�
*e���iR�k���r+�:p�tL�j����}iI�gˠ�̬V��W+u2����f�m��{k��X<(ka�-&����-'V�������puU�J++5]�y�04�n�V9Z[3��n�$�=	F�B��z��S}�	�~2u����W7�h�H`�e: %ۯ�����3!�Q"��P��F�NS兾�,0~��=ɇ^��}�4�i����kt����`�*�� �B3m+��KAA!~1P&�"�v�Q�Eߧ��7��ܿX	*�E���F��|=a�gF�ګk��}K�Q���ԇX���y�+gzܮ\�0��6�<�f"�eV��m>�O�{�MN`��,�
rs%&p�i����#��A��������XD2����Tk4�gX�b�~LI*�e���5[�� �qu�G^Mu�50q^8Yg0"��5�[��
�����-<��v�Y'�:�����0O[k,�6��j�Nu)*�'���N*ޞ����8WUֽn�/�����(�r��mͼ��sh��i�4<�g�`�h�{r�?��Tز���؛�U�oUT�L�6��Ĉ3ss��E�U����������o�tX�q��n/{�����9j������
\$���S����/����9�}7��K��96vi�3��v���/�Lԇp{,[ˈ�ƌ#�á��h�ρ�˲��� MԭQ��(�V[QƮ��&߶?������A3Q�'^�+����1���7'��1N�o��ճ�+��2����4Y�AV0��m;� O[����SJL_�u�32HA���L�?�o=���D�^�&�F�Yo�����d�IYWO���/ ��y�󍎟�N��;a2�kX�� ϶t��������Z��x��X%4�7_s���%]c��/0]m#�kL1�%)^�����gez��b!&gH��nCK���!�ԏ��je��
#z 5���#G�&,� �׳��G/��/|y�Tp��n��k��s$#6���$���<�.�bl���,����k6M�S�/��-����^���eƜ�o���	�^�WI�w=1)q�a��XݕG��qS;ϕ\���Qebd��m]�aƗM� �-�iw��������<�B�@�S�P�-?;����T��U\^i�\�̸�G��++��+U�K����h�iL�r���p�-Z[[�;f�-���"�wL����(ur�4�Z?^�Y8�Z`�N�3�O�}�LϽZh��_���<.�M��Z�Q����D��ܭ"�)�z��(���t�3�+�XZZ&$'�V�֑-�|�;y�O|y�������U/`l[�Ưe9���%��c�܉*'� ����G�Q��t���XD�:�I���o�����v��R*���ؗ�X�i��%vvV]�z��R�s���U$��������i��-��W�����h�@� =���k�V#���
 j�┅RSeUm(����韈�tOA���������T��U�Dk����WRΪ�G��*6v�����lT� ɳ���y����M�e�D(��*T�hd���Ţ~/Y{���t�<zh/�H�`~�21	ɚSU�'��)�JP@(����3%JJI�s?�19*_ι�T�n/i��2�%Sނ63�@��(M�����S���3�tM[k�Y��D����q8A����I��P[`�`��H���XY5ˉ\���؁���)� ~���n���2Jt�˲���S�{�Ղ��D��b�|9�5�o�oZ8�p�����d��o`��ؑ��W���G��� ӗe4��Z�F�9X	ӈh)�ˑ��FB���лIQ*^{Bc�P�4��s?m��i��k4S�@����Z��T���b�:�.f�m�g�Oګ��]F����y���Kp3����P�|b�!BCP2��X���g+
~�ω��>5o&=���Y��I�+��zC[������p��O���oX������]PP�E>>9�zF���t����~��Z\>��5��cm��ZUH���?�4\&������v:*�Rn����k�Q���w΄�)���,�F���𐽚<b
���l���Q#�đ��U�ԃ��Ы���]Ϳ�7��ybU�|q���7��p*����e7����J��dx��D�4��חvA N����ݥ?��o�����e�K��w���t��pQyP
�璘7�	�,�R;�,���d(NZ���"О}�/T�P�?�3H���f�u9]9��X�Ntrv68��7k�X�m#�lY!\��\-#�F��O�J�W�U��=��v�A�B�;s�.̀�7ͩ��ޞ���t��<f3���z|�8:���B�����x� �_S2%F����Y/��r�C�����P�_��뫜5l&ggǕ�3��1�����obbbaa�t~s�qشmD?Ԥ�c�"
Wm�2p��L�^�×�l���7���*M^��(��s�-F	,��E3����g�V�NN8lm�T-���w��(�ӻ���/[(���)D�1�����T�1߭��D�f���yC���
܇`��d�Q[��5?~1���"ֹA�jm���T�YYB�-�l�/��-{m]�'�}�VV(����í�k�~�12'M�A��0
�h��Bk�}���~~8N�Z����⇋3[���X�n{�����b)C�K�1���j6��yS�Fu�4l30���*$<�f<n~7�_�#L��;u@���H�9��*�~:��Ň�����%b�������f�5,�5-OO�F�Hy���>�x�'��u�q��P�߉�MA5������H5���r��_�cޙ5�F 
1O�t��� ������j;wT!�v[n`{Z{ҵ�,}%%E�ݧO����m~-��۷1�.��w�9t�9��*YNurv�K����jV�k��X��T�U%c��j �p{�z�#ҩ����Ήm�r�)|Rx҃��p{��~���݊��ʒ����ů*��}�N/��׺�N(Ј��HHE����;[����i����Ɗ4Cc1��"�O2r�{䝐邑�F�D}܂ہ���#�,���n��BBn~4x���e��e\]]��=�h7z�����V;5D�4/�<yO�?��:�'��T6� �2�NNn<�W�&5Qu�5��D�Eg2�P�F+gfvV&�f�������x:��
�onf�"(��5&
l���ꖂ�׆���ߪ�)(���Kʩ�w��/���,��݉3�W��CT5W���gy��7�\�>��EFg
8#�eH�f/�L��}�Ŕ�?y�E���f/��ۧ���<锲�o|�ch��L� J�^�2rq��7.6:��OZ��T�������c���ۓ�����On�zƪ8-sG���_Q��x����Y�?c��K@����Ωoh	ѪGƺ$Jq�8�%�z��$��'��WP@GDD�j���u�������]�M?Qg����|�0(6���>��l�� zQ/�~TQ
X�5�~�=�����(�v�5�� Zm�L�In�3#���Ů_����8K�0F��5���Q�䬦7�Sރ��i����oŉ��F<��q�*�:�Ö�vkџ��jm)m2���hT�~����`�o�~��k�fRT���w��^�:�<��C�L�f��!��E�~>4OI�Ɩ⓵��d�x-c2���zrs��w�-���{<�ق���(,d� ׉������x1�o��q�$멈��?d�P�퇆�|~�.v�P�����Y���`~Qۍy���$�zF̈���Ϧ��
l��u*ZZ@��f���N*����a<���(�Z��o������4��,�X��c�����i���Ӧ���z��+Ր�Оw�o ����B�h��H���2}�g��W��4F2W��3<<��R	#����e����v�Ҹ|H#bǿ����&��BGrV*1)��[Q�)����k%��
4D�KQ(F~�b�n���߼W�7���t��?�0b_�	/gYiދ]th�z�L@���e�s�>�Qj�DI�¢p�l�I��CE`������2�T&� �������g������9�0ho+r�u�Y���l��.�ަ�>0�r܏�m��j����M��^2�LI�:��T��U6в1�5U2|0}�v�SA�s���vFT�Q@�ڇ�	`$�C�����'����w�Yf���A�ЪRZlF��J����ᚡx��d�E�Qns��D\�U}�Ѳ�<?[�i���@o^��g	�����8"������)�c��w<8��&��{F2O]_���4�x�G�̉�x��<�n��_C^��X�k��6��*�k���6]�����̞ɚ�u���?�U
+��2Z��L��_:���U�G�|���vr�)2�c�XC��Q���Ι��߳߿����|�K���_k��"K��l}�|����qn�s~$I��{�����Xr��G>�d�%n2���,����4�<|���)����J��c<�ZFn�Z*��p1S����Z��%�1�GtDɥ=x4��(ꠓ���'I�M��Mӭy׼~;M�d���>�_.eL�q�E��|q_��m=����!Kl�D�L_�1:0W#7�A����sz�x�L��������X �+�8�Ͱ��;�#Ńlgk�sw��@L8g:P�aJD����dΣ��*���dC��}��=lg1f	�׆�-��A�	�������b�ʸZ�W��#=i���N��V�g/)/GC@@��Iw��G�8�>� V�>>�w���%�U$V�ݬb���k{V�h2���%�码�y��F;q� ���X�[&b����}�F�}��m�"�T�E�-�'�qq�iԫ������jd%�m2�	+�1�g�@�5�:Hͯq�{�7Q��hh�n�����8e ��~�����"���ԞjvV���
�Pk��F�I 	���vI���9|��y~�!쉓�L��v0���nT��.�mn
Cv��*!"A��ك��Nt�cY"Q��a�ጭ�#�{��^�	1l*���1׳��v��Up��ܡ��]5-{�]4���1.zII��޼Y�-��<����I~'���J<C�p�Jhz�
��`.���ҳ�Vd�ӟZ)&�98kv�q~h�G�N1��157��E�X�K�P�N����N�j#�����#0_�g^4��P#��iqͲ�/�����"mr�01��s%����"`���_��V�Q�m��5G��K������F+ѝ�X���vv2JJ���狳у;j�-�o��[0Up�NG���(s�|���-�C+##�G�����4�������Y�f�`h�&�a�ͤtl������y##<�)�s�l[�#>25�s�ۼ��D2�����
(�#�6���b�՘a�
(*��jgv4d��8����A�q�ܲ���������?.���\e�I�:zVV__ߥ�J��#���\�r� |�H�k,x`k.W�1�x9~,.'f��o�=�?f�Lˇ��w�L6����2^�}������s~|< ���u�g12%��i�X�u�;.��w�J�l!���+U� e�����q�\�h��ŏ[[����>�t��"K��D�_*-eX+s���]�d��ϙ`�3�5�:՛����c�ǘ�����k�q��,�=֡�����!y����%&r��P`Da�'L�L��-�v	�TS������8����|�AB+�*)�lI��w=��'>���@�ro*:��~����)���);�8/��)�n�Z�iK`r8->ԋ`]Y9�:��+���=���r���-���*�ꥼ�ֲ�Ԕ'��sz���8����2"N	�`�n|VV���M��!%�7g*��{�5���� ���9,��R�P��z���7���Y8������> acӈeAǦuc������V�YPص��O��n_L�mBg9�����TW�5f'��,��ᡑ���-�d��������1C�����c��[��rƮZWhƮ�`�蒝����)���D�juT���"�ņ�SdXh�\�%[�vOm�c���d_�-6���,;��h.��H�i��Hۀ�KMM���Sh%6(��̬ӆ��Ɛ�B��"���ݼ�JV���9�>o��C���Zڷ�u\#�+Lӕ��׀-:~���eՄp�ֺ��w����	&HW�G�pc��ũT/*
ʟM6"h���HRE��ʹ"��\���T�����#����\;Dѫ�_�7G)u��P��0�"5n�4�� �`������@o؍�,R�s��u���f1���A�,l�袈W'��]��Y�?b���,��j��)��c��1#��҃�HN.|������oB\�~w��q��ᆮ���$��Ze��=�L�unYD�*���e +��]�O<�e֯�dBj����>}
�y�i�pf�m�۽}������><�\�MdMhQ�z� �@�b�,�(�� �ê�%��s999)��D@;U.��13�lr��jLU���IH�;��>+փ���H$ħU���B�V[S�*�0�Q�^�ĒvڜLF��I�O��X�C��gg�	Ѻv]����d>c3&Ev��K �$|��C+�2p����^�v��?�g�o�L���<)<a��S��x���9llU�I$w5
��Ɍ?��u��Q����*>��J�������Y�8��*d��Ԫ��7ݠ��5��L���
M��6��{-/l��W"@��00�aa&�����貿�N����ϳ�~��&��b�f�����:}/�	Ϊ�7��5IO�I���xrgh�kc�:�=���N�$�/eha�����-�`�!�!�f�kD�0f5��i��J�7y�!%S�[�����J<-�7�_��W��F���)���5�:�.�A����NX|t!C�f��<a��OU��p?m嚯�2I����N$
)�i�&=�����m"�{>��^֕��'�5��#h�nU ��'8�)J{���s5W�ø���c������*z��o�3L�8���_;�����1�0���#��(>��\!0^��*)�V}�z����<��8&����Dl�
�VU!�f�tܸj�r�Q��#}
�`0��joCg�>����?䞜�̙���B�U$p�f�'%'�MT���G1�X��p�9�+���81�k# ��;�J���������]( , xcs���{�7�҈G8O���t+�y�XJ�#JK!;::Z|m�g{�73��!uO#��9Ȳ�Y#G��q�cfJ_���S��Z9i����N<����6�V�y�z��R����tW�{xl,�7�����kﻃ�j�6PA%�  �H��T� A	2� ���� ��J	CP��� q�9H@��4����}U��ڿ��ݭ}�nz���O��<�i��n��EO��P�,��R�|.�3�S�b5�@3��� ��-BvD,�8XPQ�Q���i5��S+k6��/�BUBpa�Ao(h�?b��_4��z}���E�w))�{�����sa�m��(�շ׀��q7��2A$�#���-+�At�w���-n2�1;>:����:�a��фk)8����!?wߑ�Cِ�b0ȹ\q&��yp�����d<c)ߗ�-w�{�J��Y,��<�ڪ:"D�Jޣ�OCK�qs"�pfNK�pesݜ�{�O���]�)JO����������%���WW����:��r��`Ik�����D��`�y��Q4u�[6�b�o�͝��s�2B���@�Q�z� w��s:O��t*�ݣ�L���祥���%�¶w�o�*o�������)2|��2��NL�Q�Me-X<�w^�mXXzb&-�9�N�N�#�*���Zr2[�I�dM��/ݥ�*%�>'i����dg��OK��!>�غ\���Z��kr������/���Cm�ӈ�Ly�����,|�z��!J
���w?>�}�i��eh�*y`�		k�]!�����4N{5j?���䐿<@b*�:E���BZԏ�w�4�����E/o�E@��Q����K��Kg����u���d�[?�+a�A�U�O%/���ϫȃ�E���Z%9@��o�h�l]�WJ�-����ܳ��*�yF�73�t_8�)�I+I�%���P���#˞���m#����\��_�
C�Q4���X��Ո�6�6? �@`q2S�a0l/�����O�I������H99��r���R�/\����c��w)�\��()-�6+y���
��/5ן���h�X�ӻrN���}R��Vh��T o��b�gdsgx>=��YK���dhhx�`������x��ƫ�v�f����mji�]�iV��`��U��	�PǤ��X����-[����Yl�/$�I�f��O�z�0�j佐���;����fVm�����T��8��뺻���c�K����Y�?O�3S���Y=�ɸ@��o9Q�u��4�dY[^�	��
�u��g�6��l=��\���\{#&�u�N/�/d`�}[T����9�[�%}�O^p�U�f����/Fg���r?~�,�|�M�3�S�~��*X��y�`��P�O넾{t�/�&ԡ��zzz�V������ܒ�7�����Z�շ���������7�|�۲��}���BU����[�A���y����*wIM�nر�4�ꈼEZWݶ�n		q^������}�M,mr�M�},�v"�js�!{+g����M��g����IZ���ƍ��8��"4M1��{����a11�ܔ�ܧ��M�b94�D.4�T%���r�,%��;r���AJ����o�q����Zr��6��&��A�����'����Z7��Np��g/)vc�\��O�ϑklGM����\9wGUUu��H@h�?�)�/�����x��7��T�&64c�^�F�q��P#V-V���gm*Ն�A8��B�l�S���n��������M���]���A��i 0"
8�]PMif]�ҾBe�GGN�'՝v�r�*E���6t�ϯ�ύ���9b���O�)E1��X���zs�p?{��t�lD[^�E�$)7�\�q�3��Xt�c�s�߈!](lcZ�b(nIk3E�^^���XY���ά������m�x�\v����9 �nB�L�D�6�p}�����WX�k��e���Q�y.Z������M�m[K�!G�X2R�UHS�Poxi�~���k3�/���55T�q�;����R��]�9[�4�9����*u�aT}�C�f�ze��]���@pp�bK�/�M�N�
���A�p�	ǩQW���?���0����8j.3�v����%L�Н
�&l�}��0Té�0^�0��KnW�6'>����'b$<����I���v7��.^��g\4����=�4�v�r�/�h�����
U���p�Iֱ�EqA��������RR���x|d���<3MU����n��𫦼�w�JdI��*oU�ĳׯ贋9S|j�3x�e��/0�D��=���fBz��p������h9'?����!	�ڒ'��H�����l���p ��#S��Y�s0:+Yj`rVI�|sCC��w�9杴�!k!Kfh���|�W��Ӈ����YS�q8���'c�Ԯ��D���ҟ��-ќބ��O��;��=_�6���wu\?<��'=���rG��ؼ)��O����N�1�嵗�0�*�e�,�L�v��(��|iY���년��./����&�2 �������!�[��/ڙ����b��Ue���h��b��$Qj�7���w�;�0.��#�Z�����+�h��7���?�9R��^_�h�A^�����p�1?�ZUU�<�r�������(�s��Yg�#ŉdWV�j�p��8b����3LY+~���p��3%L'/P�!�Dݫg��Y�Q�Wu88j=��
�B/���H ��A�B��J�!UC��0��34�$����������o�|����xx9ꚜ�A���@�O?��b�J%���nJp��������>B��%@,��+�]}��b��Z� ��Kz�wXA�:@� �Y�T��Cg?�ߩ�8]�pbz�Ò�;�_<F}�S��Ǩ���d����N�J���Uv��LM�{�z��ēf��~9�j�R+��|M��߾��ֶ�%��2ņ�䯟Rd0�ki���v��di1sf��݂?�\Y�Ys$��L��3�,�2�ï�d����G_v\ϟ	����gG��e_��r@;Rg�-�O�i�8�C	���������N5�팭W�����h��3����^�e�
!t��KnOU�����ξ�k;鵵�qO���{��V-��烊t�F�hAYP���837dJ[��S����W�#�=79����=*�UK�V�'$�y��*'�f��>�o�����(�d�������e���N�v��i��1������A��j �m�����Z�MV�
���}N���}����m�S�F����|i{YYY|��[^�S?N.��ә�$�9�,�?��s�4�qȒzx���4ɚ���A�ӳ�x2<y��wБ���[s(j��5���s��L�	j3>
Z�00iܘn6ÿ[�z��-�w��Ƕ�W�����C�x��)����j_���?�Ójc��7�%�	_��cC�?W��t}(|C~��"%>*"<|������緖e�Mןy��-r�l��5����v�e�q/�t�z��y�B���Y�ǩǪ�����j�x[�|��>��ܘ������/K��x�W�[�����b�H��,��_�d�ۗ�e�iD� ��킩�"�4k�[JA�wgx�����'�����ꄩTmLMa��o��'֚�(7@|(>j�~�]�����	 )ݶ�+�TW�ƅr��z��`�|ɨ�~t�Tο	�����۳����ljjj�7i�L=V�m�nd�cbB�L�����U/����_��Js�1�g�0���[��1����u"?Ǘ.��7�&C^O5�b�.:o�d��$[���"��iLLB�	���z�	��7~�w�����8�$0	U�zg�@��X_�Ǭ��T�*~�/�![�-���uz���E��n6XMr��Ϭ,��)����zC�|�"�oXr*Ϡh��Ή�ͽp�8�F�{'zztj�3�]~��θԂ��+�#�ON�}��������F���N���s~�x�{	ZMC;�w�[x#4�tI��M5uuk���� Pk�DNg���Д��P|�.�mc����f5���S��O��i�l�X+}(�|�"9�詩6$���|u����W�Y_��ؗǫ���9��$��"�O������_�$���Ă��N��O(w�*�]2��>T�'g�z����©�̀�+�Κ�~$HN�XM��MwMr�y�f�]W_��KJ�;����;e�+���wutz�y~��כ��>;/�arr2���ҘWT�vd�V�n���J?��M�����eS��Z��v�Bϯ\
�z�|�wB��ڹ�+��ܱ��;� ʭiA�y��Y�|a\�P�qhh'��T�忬��ʹ:�`Ɯ���l�� �jL�M?� kP��g�?5<�@3��sc~��|�̫!��5O�Z�̀Ȃ
ϊ�}��
S�cs�����dZ�@����;6F]�m����u\Z8�&��P���(*����Oi3�~�
W������rSsT��th����Ubݕ__}����K���R_���� +k��@�6�O ���3N�{ܧ�C̰�̑ryWY�<�ϝ`6��������@�o��j5�9��ԊV�J��&u�Nhk�&�_�/^@�5pq�%��3* �}|H�Y��&G���0;���W�㇤,�6}���n���1{�$�,#��B��o��U��禃�`_��|R�ʥ_ ��b�z�(bbcc�
������$ ��r��#�|��QPi_�R;�`�X9�Wv&�8���Q�ߢT?�$�%�1��>)r��e�UzEI���O55�}����oL�\�HG�<@'S��q�k�8T�Z]��q�0�R��UQq�ߓ�A�E�̂9?y��o�_���&�ȸ{���>�y��LU�Ж�HH��+�~>��
4��z��4���7 e����ʅq|�ˠ&	*�5<���y;sZ��\f����:�ӗK)ھ����b|�?ύ�4� �ڦ��7u㿢>7�������
��x.hJ�L^�"/..���$Oi3~�ڪ
���zxxX�QY���eIg���q!I�	K��%�"�)�t�U�AjЫ����ݳ����Q��	��ł���\�/:�t�T�ղ����o�Q��;�'&"�ހ��=iii0��Q֫ka�����m�ݫJ�b�^��+�/�6����[�B���q^�(# 9����u����`h��m�-�[Ё�P�,BI��G�=EE�?��f�,��.������?�n		Y�����%�[��
�Zu���J�֌iZ=3���kkz�+�M�g��Z�+�V����t�����p=/��nK��&m8���j���Ů��"u�u9���3>��-(��Zg�ߚ,��֪�����'���d������D����;wdd9���^�}�+�h<��.��������K�J�j��:��Pkq&s 
�Z[[鎪�7$9��t�]G\�~ۆ�E����kb�w�I�n���@��1��U؇��i'v�8a�����~;�Y
O_���P��x�~:h����"j=q�������_T4"��uVm��Nܻ���g�'}�@�.�[�P���1?��ʁ���Vqe�cB���>�b����(1�*���[����t�"�¨����nk��AW��?Ǘ>�y�K��w'�j��F�DR"�
��3�8r[ZR����ow�L9�&����6G'�ă�:�>raǇ�����r�3v�z�]�INW+(��N���	����?��:>���@*��df=�u�pHf�x��'@
�� :w�'o#�J\���>}�kkkˠ^�z���h�ׯ��P�M␉���ZJ3�o��O8����Bzx�����Gyo��r}��2�|z#CL�����X,�SM�]�k׸���1��CKO��J�J�i壽�c�5�1��Ǐ�-#cJҘ��Qu�3ͩ Y�轻>ߡ�mO�N��l�BG%]om�F$g���Ԣ�,O�w�K���ߐ߆i�Dt���:ZH-�l�&�G���Z����z��>/ �@o� ��WMߘf��+��Ϸx������!����jo��.1<����|8���������������F����?�ܿ��rʷ��9>������.���`�c����K7U��Z�ݜ�_p7�:Y�x�XO�$\�-��M��jA<n`:��/ak��yΞ=��a�{!�Q\R����X��s���h1h4z/�x7ꀄ=��'-����:��Jv�C}�{�<B��G���
��!!�x՜�g�"�=S�'�L��/�d-����8d�fƽ&p��{�5�ۣ	h��bꀃx�ׯ�@���rq����I𬶖��N�[_���ǭ�:zzzWW�7���''��;Mt6s�')L�I�K����MTG��W�4�3-���pmm����cv�m׃�m�q�)����Ԩ❍T�u�OuH�M+��z �<'��%	�&�7<�̮�
��r�iE�����㠣f���'	Z4��b|$�Ǉk�@���1>�e";QC"�t��a�k}��^Q�Μ]b��|ŧ��Δ�>�;�ܴ���5W�fw��2���K�5︮�RJ�;p�l����V��ks��}U�'�z���8�x�Ǳ�\ve)�N�h[q���OV%���:����L�i0߅��]���544\fg?�r�U��G�t��M��Z�&NV�qK	�P�(� �BKS���Q ��o#?�\��U�m*+J�u���c��%p�K��K�92'�晰���(�
d@�
U��k�j��;��45��F4=����&���2�;8 ST?�:�<Wx�."" �+�����J����`���Byi8��Gy�}��}���*�*�7��*��̬*v�y��4jb�LZ�����ph��9���ŕK�� �����<.Зz_Q�rz���꽃�.7 �yLT�u�C���$�}l�Fᩢr4����r�P�d
���t�����ڳ���pv������Ǝ�CL�_�o��׊,(wo�?�J���#��G'n�l�v��_��t��Zk�JE%��#�P�Y��2�-��A�AN/���|Y�Y����12�F~1��ӫ]��ӫG�*�^��7�J=�ӵ$\��#�':֏P��܀n�p�\ZZ241��L��O�,��L ��C\�]���SVnni��/{�d	�^�[�a/.���2Ԗb+�Gd妎���5�؉r�"Xq�0���a�rs��WI}>�Щ�0�6c�;s}�!V	�@����Y`"�vV�ۓe�\�����~R��������/(��`�}̨���>��7�L������ĉ&����.-��Bd��w��n`����+	\��`���+���A�����VSs��Is��� <�spP������ƒl/��l�z�j�uFd�;dn��ɸL��&��g/��ɶ8i���<1�ٚ~X�P{Qb�KD{�m0IU���S�R�~�UU�D"�pW�ã�J%_''{}|dXYY_ .^�����Z���4��\�s)̐A��,a�d%o�n���Ӂ�kTP��
e!L����M1
+�_ëZ�H���z��j�|H���t����a�wَ鈣Z���4F?O�Y2`�'ة�2|��7m�#j����M��g �Ŷp�ט���!�b��/���\^��,*t��	\*b@���鈝H��=+n����s;1��<;;"5�,�*h�lV5���=���LLǿo(0(�_{B�555��r<d�<����Y�6���I��Y���4bn��-c'�ȳSr�[�U���l�&,�a�1�vz�E���=��KIIĘ4�:�s��PS{`��Vh�^�M/PT�i���4���!4("�c���9�K�ƖjRjJ�0�����S�MX��f��?Z�](�j��*���z�sI0VC�yBȐB��'���������V/���zP=��;�堯�V�:g��7[�v8� ��^���V�ě~(h8ԠD'�ʵͬ_/i�ٗ�#,��k*}pT�����W�^�H���;e�G@���3!��[׭�*Ѣ���zzz �o'���Q�Us_
����kC"�� fZc�0��Oh��&o/�[c>���V��o���qݝ�ie�\@%�ɪ��}��9W�.����w��)I$��x��1�I�+u��\�����n�� �-A��{ˇ�?�0a�f,�uR0ǃ���Ta���-I&x�������[�ܟY�X
� E=L ���*���}�.�]� ���R/����~�٦ �Xa\a������$�n"<��їf�(3V"Vz���GC�{��rMlE��+Pi{�G#����f�uia��rԩ������^㕌�}W�[�d������'n�qs�$x�v��hf
�z�<-@�/w\
�1v9��=h�eg�=�F��,#8��J��4�x��v��k����P?�i0�2����ና]�D���Y�"�/�C�H)g��j���+=9���x���,<��4����,�� ;oU��t�`���m���`��ziZS�= �?��U�s�A�=��������L~�O�n@�(���l����cd�\���5U�˂�d���S֏�/�L����.�@���K�o���L�#�5�/���4�p�t�3ܦEk�8V�g����VC���|`���y�J2�*YS��&R�Ԟ�D�S�`u3���"��Z��m0�W=��mbc�z�X`�&��shel2��ļß����s2�5}�36�1����.��e|����ϳ��x,�Nn�f[��f��u6a���յ��R����`��88@�� pK�݅+ ���;��4��Vp����'`�Q����$փ%a��:D�$/��.)�d���nEn0�[%<o�.ic�\Ztˢ�z�p�(���h&E==���'y����a�A�Vrɬ�c���I�t� j	ʄa�XN.n��ڻ�ᩃ�0k���tUet5��0s
�m��b��MG�[N"�As�ڳ.*�6���NDl�w:_�w�y�]p̄i�7��P׃�f�Z�ؒ��f�إ��]Oӕ����G�����f,���+��&��sEH���ZEmc��R-3���X�^n?����OZ��Hl��?�8����e���m�L����e,Y�������eX]��i�n�n�p�71�C�}8�>�|��N˯���\iL�i ��4�䟼��G�U%�t�"x�6��{st�G]'��'�������u�1�`��@�p-��U99�SxD��{I(=������S$���`^��	�W_�1ǀ��F��-���f&��$T������}��Y�TJ����m�9�T'Z��9B�0}8�����e�����-�����W�S�yHqT/O؎h,u�i���h<���1֣�rM-�M��x'�g䰮7Z��:7�#�\s1���vE�W�����ǈ��	��	��;g���p%Fg�dD��X�u�� <�����1¾���M��!ĕML)a�� ��� āh�H}h�@d�ȋ�s���o�]>=;̜퓵�$���P�aB�늌qs]�mx8Ǵ�Ͼ^�<�g�P��,��7}���x�CK��_������)�6����~��$t�MB�3}�m������;~�	��|\��Y��ȏ�9vO�p���+d����ui�;�`�mґ�tDu����[$#l>c��^ʫ%��t'������8w��i[�t�HT^N����\�28J�����\=?|��fM
���>�Im ?�'�g��ȧ���z_��֓���(�Ubw_�U�5�^n���ʡL+�N�]i",E��NrVP�������k~V�`�D'����l��=w��gݜM��.��vy�X݉��(-+r��>���l���->���g��W�:?�i��a�k!0�}��Ʉڙscd�v���o����&�H�0F,�ٗ,�ǁ�����K;�40cZi��}0C�550���2MT�5�L���������o��C����Z�Y2�h����~�ۿ����ټ��9n*�5'�@���׼W�d�? PK   z�X����U  8  /   images/68cd571a-d128-4aaf-a06e-233b43cf9b16.jpg�VgP\�NHB�!�л�4�R:�QQP:*H	AAAH�(H�A��&=4���/��;"\^��~�ϝ�}{f��9Ϟݝ3����׳ ��U��  �x� g� m �A�s�@(�tT�s���R��aLLp��ƍ`f�d����9yx�������ܼ|��?�RB��xY�,��o9k�� �iP@����.   @ϫ�o��k��Q��&�  ���������(@`��������7+B��e���a9ylvnea�MH]5"�������Kȩ�q��/���;�F��� ��Ϧ t��tp���hn�IXl ݽ��6N㇤�m��,��E�W�2!����{�%a4&�}Yj�t��*+�c#������UOI�`M��ο�١����(|V�rh���5*��A��u�3@#���f���r���Gyr��\�!� ��_m8e��(�˓�_��ϧ�����iRbȫ����py��Ո��Â���q3ubi���w�v��3}C��O�}�2b���L����'���y��D�U��&�	%��f�e�A��u���?��v�.�nZ���G)��x�c����#zɭ�y�'���r������G�u����`�B2��ֱ�_ɥ"�wKZܔY4n_��:��v���*���?���qu��-����^K=�U�3��z��,�A'F'����.�ߴK��=H��U�#х��e����Y�C�����t��j�����wOp�户d,(k,��cpsj�{�(Q�D����	N���8p\c����I������I���%�UU>�*��X9yO6|�ڏ7�ӧ��jd�	
R�4IN���rz�J�jo�ۓS��{ڏ��Ի��a�-��*y����\|��"���7��ث���!󡛪`����M7u�>�`Gq�qr{�� W�x���c��w����M_��8g���9�՝���X�?�č+OyG�0X�-�UX��I\z�A؄y��B�#_�ڱo���������}0:���� 5W�������=u��5OG�z�OU~ׂ���]�aBSSQ��6�_�Ѷ,(�ˢB��7�B8=X�bd�U�S�v�W���`�!C�VGQ:�+�U;j�ρ���D��^P�E�o���bk����4*t�&�b!�����M��I����iu���N1g��ށ�5$I�P����x*ǯ�qƕ���2![�P^�A����w��U�zN(1��W�^	FK�_�Q����Z�y	1�`km<�L�d���9V��=�Y��f00�I�<����e��.�����OC�r�7=�A=%i*�#6P�`ˢ�2\^	�n�@I��²X�ύ��߻�2"VJ8�[xL� �3D��<��.d�<�G_[�\���'�doPI6Cq�C��-�мb���F�|4��"�|�=�u`�}���b��Rq��#aw�V=F �/���`3gnh��xk=�~]��?�%2���ҫ�+��V���ͯ�Y���RL�����
�����[�+�I��7�ڡ=s��4.���"������}s����5�ē��,p�����������N��+U?�#]�7�;�ݷuU���V�	/{r�E��x��liQ�=Ȉ�ORhչ9{��_�W���e��x0�<�|~�b�o�Л�T�P��L��T�{���@�H�R�l�5]�@ee�)7�b7!3)0M�4���څy`9a�2^�pgZ��QG$,�5>yQ����?C� .z-���������&�ۈS��:i[��1P��<.����#�I��QQNa_���%�&��k8���P����X~O�L�6u.��P;�(~��͆L(^�"�&3�$����C�C�T�~�K�|��H]��sŏ�Q�CЋ&<��VP��	ϔQ;YtG�1Hy�	 �m���n{��De��"��J���D����*����;ֽ!��M�c���+d�ұ���&$�,��J=D��ʌ�a����U��Sr�w�vNK��(�4ͅ�\.l����y!1���>��m�<��7�nL%��J�fY���@���@�bB���U�;��}Eș��A�L�W�(�0����<je�+�=���x�Ǵ��]י�r���"�"�_��	�u���(3�(��k[����#|�����_�P3�񛱘�û�m]���U��4�Ot�7���Xcf~r����|����I^��mѵ*����@l�5"�6|)�hH���ه̴�(;dJ�њBN�0�ͨ׌�*c�H	����_�9���!$K�!K�A�ž��=�����?�����`�סϚ���-sJa���R��!�&D{�S�Ǆ��
��o�:��n����F���ؿ+V��e٩��\�����G�l3�����_��Zt�"Q��(�',�y!�Z���[�n�n��,��-�����@����(�>�QZ�Su��Z��K�[��>�\�ʊR���ѲQ�Z��A8C���0�'�Y'��#��xC0�Le�(��>ˉǊer/�P���<"�2�Q�1<͚�"�Qt��ͽ�ōw#�����y�SfY��nu��_������.�Ʌ^b�(ź,��k�6y>������W����ǌiM.K/;��[���%�d���$�8��/��W����^Ej��3���Z�+)�"�2QtvLۻe/�;`�(���Y����8�X�f��&Д��]�M����ɾ�m?S��K�J������eu���c�+��-�G��X~Q����]�p��>u]x�(HZ��o:��L�D��;>�����Y�JP�ʄ"�"�7�}VJ��l��iNN;��*��?h�X�w�0@��+Hn�Ĕ?fn���-�ٜ)��o!aF��i>gf:��ghN���\�YBݸ$�.C��e�U�e�M�� �ԯP��n@>k�+a��c�t]$.��[��^DS7���b>}N��Ɲ'�)2 a��%'�X��Nń��D��3 ��U�P*rH1������@i;�@��ְ���|���`B&����c ��o}*�9-:�$���xo�MM�]����䖪��"Kd߽�6�� �[�U����B_�
����h�����q.�����
�2fz5:��GA��8��p����}��Ȥ�Z�Y�\[�w��O�S��7�_W.�_y}��\L��Qs\�zן�e^>��9��_�N��2��t��q=m�-�˹#�>�	:�s˸�Sd�ŋ8@��q�.=��������0�WD������ x���Qm�����E攝�^тq��qi��!���ӹ5M�.q?����RY���e�f����JKf��#.�#����r儭�C��k����p�`X���%�K�����/�k�klHs��=��u��V�$��bb�����i�Q*p��7�֫G�'\�'��I?^�dPr�H��R�g F����:<�p��ka�oeo�_��P,%��w�7>\4��h��7�%<���u��[��i"pVyItp3�%]��o�W�y0B��F��΄�j򶄚���w^#�k�Ic�}H�MX��_�b{Q�{Rw�I������a.�c�O���������4ui�;�1���U.R�9��l���0�wr�.Z�l� PK   ���X�\�#W 2Y /   images/72f7f29c-ad5c-43c9-9f1f-56c5e6d4e935.png��S�/���@� A�[���]�����/�www�w�� @p��|�{~������f��9ݧ�tz�'\Q^  �HI�* �a  D� ��M�h$���;{IM' �}߿8dWj  R�B*�^�ej��J����i>�6��t�D
@t�ԭ����W�A����-i�BC(���@Q41�e��[sssϊ���ϴ��wM�|�^;�]S
���<v�£�è��6�|�ڴ�E����F407Ĝ΁:�Rл����������=99������P)���d�U۶�����i4�V������X��E�^�@+�e;����X��j3�H�{N���aⱋ�6�P^��6���@���M��g"gF�S-��om1���IfC��cw�S~KEF������mԛ��5��Q}���������1{n��p���FU'D����%n��aΛJ�L�r�uYsu�M�v��T��<�T��#�AL: ��,�5��EEE]302")�q��p'��E�� Y�Y�������6x����XȱZ�i���0p�FLo�O�կ0��ooG� m��~��,TFh���x�ۜX�+8�!w4̝w<0���z{c�N���N%�r

�{�(�@� X�j��;;��GG:���H�T{-	%
�^����H�o���S�-"��b�{o�ᑗ���Ò�M�>'�85�!�?댆�����5}#�VE~��!B�06Ȧ|
ف�~��-��gĸdaI�vwq:sQ ع�cT�lA�)ƿ���>�G_�����el�B���'j�]�ؓ)޳a����?��5l��Q|5MFsź�J����@T_� �Hƒ���X�z#�R�Fc���� ��U��Xv��T�\����^��	�#��H���xqĽ
>�X�Nv���������.ڦ����r����D���=R$lq���@���w�5�n,}�l�7���� �7J��!F;��<�P�z`39�;�+���1����?�v�b�����ϗ>�{��i���]Rn_L��ݼ�Iw:�P�끢ڨ%?�M�|��с����vDDDm>��OB�fC�c���.�(��>��}&�$-�3�}��ߚ�2��5�s�M�:9I4�Ԇ�#��P�z/�d8{���X�%�]�O?�{wf��D)K�#�b_��#�tz�7�U��QZ6�a6P�t.���`�k��/7��g-�����{�x�^��b9o���F�ڕ��M	D xښغf��HlF��C	�����d���נ�K^�)*X6�m-}Y�����4VX΁!�BA�a�C��5�\����5�.Q�St�5ږ/t5}^��?O�ʤ0DH�T�3�VW�M�&ߊ�C��\D��i�@�Q�[��[��Հ��4�/jq43_���I%�4 ��x�>�^C�qN�۩�up�n&�~�R]6O��4Π ��d(&kszn�in~�B�U5[d��f�f���*g��@1R\K��,CΓ�4]���4�V����ɩm,eh�����\��0g��]u0� }��mj����Tz1��X��hu:��恅͡�u��IR	=�'hWP�o����V��X�$�j�H�*8l��|_AO�PѦ�sv喼8DS�����!s>��������v�?��Mo���2F��No����Y��1?i3��=5-�u�GM���Ho�A���'��~`�	B���	M�t��d�5��'�K�?Y3����hrI��������SY���L&X�]��v)�^`�{0z��u�N��>���'fcc���	5�Y1�%>}�&��R�J�` � i�t:+��1��.G���Kǡ����w��iTW7�M�\���}a%�=�1	�I ]p��+�%�����P'������X�E�W]�%�B���~1�P�}�(,�V�/�SVnP6����:��N�W:;����]g��^�Qj�V�b�)�7�3�x�U~����K�ۿ��i��䰚��lk��c4^��t.MXI8��b��SFiZ3����'6���5gS�4KaB;���T�4%R�t)�����{8�QP�Zc��T�����:�k�K�v>�g؉��K�ϯtJ$J�0ʽl�痗{Rꩁ��rc�׆T0q���D,���n��_���Dz�gy��`���H	���VV����</C2�CF��xv"쿛����U+ik{~,*�U/�<���7 ��yϼII�\���M�.�k��*��mk�q8r��nUJ> U��5U'���U���~%!�4�̇��?~.���
�m�Y��`��~vo�˞���� ������nnn��e��޿���k��_�͘-����^)��fK��y(�F�/AEU��h d����*������=~X���e4�MY��k *���5_L��M�k�P�P�᯴h4Ӹ�A�3��~�� ���s%
oѩ��ҽ)b����V�EK������A����=6��6�����Rc���.�c�d`20/8���*�*fll(�KdM�� ?2x90�� �Ĝï)x.׭�[�,Q����w�"	��W�@eD�v����_:]\]o��]����3t��,m�G^��}8R�KBVa_<��Y"U|I���@iKn$E�V�۶��e�9ъ�ڢ��O����#(��@��\�SX�Ľ��p͝�\:�e�{�k�?��J,lxi:�z���/A<��p��A��Z����o��_���n%..�_�3HC���=�e����D`�j�J�03_�v뀼yr�U"A׺���X<j���d ��~~~�h�ly�W7�v��,�Z��<_n?h��b�b������5��k�N~PI�,����B����(6���2K��|I� �R1����v"�+��K�ŠPӷj�)�l(��-��5=U��H�h\���-�^���2�渌�D
w+�L��z�N�]R�k�#		)4�/�D;�0�I\�#�Z8�d"��� ��f#�2E�H��آ�r �7Icg�B\�n��4J�)�D�r���O72��V(|�	�"ﲂ�&:Kz���j~)��!��߹~Ж4����O���Ws��Φ��ڔ������{���C_��N�+�Z��x��Z(�kC�k?��q�s�5u�%8�kka����јZ?�+
3VM�`���p��IX"�N��W���|�;Ú�!��6'����T���6����nM�ѲTg�t}T��c��+!�� B�\'��Di��غ"�o&X�}G�������J��-2R���^4@ve"�U�������:��X�m�����`X �O1;�`��߳A���(����'V�e��]�C�^��|uٷ�G)%+�Q��.ХL[Z:b1�Fue���b�uCY&��So��%
̓�V���~����8v��y�xB�84��k���H݄��|���>C�I�ŖMp��a��k	 ���(ʏ����h�ŅmS*	sKqqUJ�y ��,��BSl�/>D�,2�-O��A�
���Y��"������`����G�Ò���� gm��<�SO{�
0�,�j�@�K�2/ۋ�[�O,jAw���y���k�ġMhnŴ��x��dS�<�g0�,,h��X�z|2���G4�����j���#,r�^J�r�%��y���t��+"���Z��C�6W4��}��mm�[�P�����TVN��j���x��=�l��q4mͶ�m�U�����������()�B�/_k�[��~khr媓���{�hj�yQ8��/e!t�����v���,}}䠈uy+�Q�PDo��%��A+6�� �26ƶ��V��el[^�q�,z��t�m�r�$.L>����6�]��C�Λ��b6	s!"8�]�_
���6-Z�Ry�C ���^�ռ�Һ�$)�X��3��v8�jT��l�N�<lAz����+|��P����H_�Ύ�c�͒X�K�I���gdѓ � (�o�x��A?T���,Yd����ۊN�[�7Z���
l��W`��nݧ#�T}au��@L]�dJDs�����+�� ?ݝ����5��0�]d��m�)
,�3?���#�p�O�D�:��[P!�ܺF���inܵo�P8��}�[����7VX���Ih�p�ؔu��^P����CCU��`���!�2	狠|ј~��{fۂ���"�r��AzU,Yű^K���r�`&M�`���E�j���ɕ�{9:��JTýS���2#7+F2��W;ɮk���S�Ӻr/nn�b��,ܰE$�2�5����jƥ9?YV}�i8�]m�6���HH��%�'55�h�h���G�~�ue�c���G(|��� ���i3N4�.� 8	�猠��e�l������Z�X�W�t��"�+��(�n�O!"st�B8�ÕVoi���Q� �7�+L�y�����_�����3�����[8��b���E��#<*��F�a��)��ǚyL���r�]������2�
5����Z��k�g�
}�� �I���M��C�$�Udd�`�SP�����m�qF�#��?�R#�;���8� �e}z1�c�;��=�8�C��F�� ��ȣ!��q��<��;�ݑ*�rbg_2"ъj�_�ƈXp���a���ć{�n[!��g�����U����W�5t�'���ҘЯqӌ:�NK�^UW�a��O�Л�e_��YO��-p�y�&v�s�b�S�X8���AEt����.��Q�g�lC��;�Ǡ���op<�&]�!Z�(�׼��-(Y�����)s�\i�H����eT=I�_�,YQ�����z���哕�GQ�~�_���6=8$����]�;z.Via K}�\:"�'/�`�z����,�F�$�-7��V�� �b�7\�S�����]@$��X�L���6��p�@����ճ���6�F��]���'h��RA��%n���ϯ	��C%>�B���-��\pw޸��K!9.nV/��ީ7����K;�-���)�N{������N mߨ�"|j���M��*co4��	5_�pZ?r��.�3�UH��
�7�/����
h���5(��i�H3�]�#ĳ`&��DD�� �0�ߜ�)TS�si*�����Е�l��i;E&�!�Tt[���%�E��B�*��5&�cS;O�YĒ���kf{OKV֐'uUkK��Ewd}�7cr����h"u�l;�n߇"׭�$���o���|c)<��.

�ZY��[wV� �T
�R��Y�t{�J�L��I�J���~�%Y'�iR�n��e����Z!�
��&ɲ�����R�����~/�kr)ۢ���]�/Wa��j����yP��ד�a���-���
@�����=~�3�7ʨ'D;3٥Y���)�o�仮�Bl����R[E�y�mK�K�
'*�y]>�Cc�l��k>��A�ޙ�����u3D? �N.p�Ө:@���xn>D�Z����#'E}��+<�'�/�e�ݞ��U�����9Օn����$�JIj~L��7-�F�����4�:k[�������i�\)7�oi��^;�����c|C�J:N˔���~�Z -���r7�+�"�!x.���w⬇&2��{Z���{��Qj�O��}���b��p�L,�Wi�I�廦8Z�|��n_ğ�GggS�k��{WS{�Y܇�#yy�3tM2�Q���	hKf/�v��җu"��ǋ��4��l'��w���a'���j����{�ބ<	�OԔ��W�Ūڣnb���$�$�0�\Z�9�.����ĝ])P����c5Ә���W]w�E�Ͻ�H	]^��hR��|K�}�;s-(��23��8�m�M0i{�\p�z�S3S~��=-[6��I:���pw�~�k	�x7j�"Q4�����a"�1r i��#��x�M��5>��B7�l��q�yo2�gJ8�����4h_������3	���>�ۂ�Vp�nT��K�3&ߒ%gU���9���`,�7'�>1����r�MR��b�8���L.�A���<�Pm&y�c)sű�nKQsvh%'����~�aVf&�ܱ�P�9�͵����uW�e$���&��ٱ�c����F�rbY��ʭ���̳w���q���uk�jtt�<�*�G?ߗ��)����iP�%`�m�1�	�l��)�J�h�OO�;CQ����Iz����
ʘ�~��qp�8��}�$>��Vg�����7E��N���b��BΛ
�w&@f�$#�.�G�W,|��L��5�������8l������*@� <�bo�Pt	_��O#�K:�MO		�*���\ '`'�"r*$$D��O���ʤ=GEK�I���"��n��L���sjGD��+
����V�_�e:�X�pټك-��>O�_P͊\Oɭq���Ȕ=~�u?�W�_k�D(�s��d4�?����-��Pv��3Pdʢ�l�j�6�z-�E,l
�m��v�pk�?-*�2�n y&��Q����/��2'��	��p'IgO�Yw���?�����F�U��xFJ	s��a�_��HJ!��YYY���1	V���Л���;�5��F��F^����Ц�_+(����C:�����N�TkS�Wi��3���&hc�د>�Ե��O1m��00���X�_jU�XĿ/F.B+��݇#ɣ÷���,Y>�y��"*SjH J625�XƟ��M�"�al�$?�����F�%�^FM�,3�v��3�����7Z��V��j�!~U�r98P5R�hH��_x����B��bh8�3oc��9�R���������d/U{V��)^�Q����0_�D	vx;h�0�ϋ� �h��a�=bNﲨXѻyuׁ)D��z��+���~��Ն����4&^���S��0�=�v�3)�w�R���[L�_;	�I��o'o/z�+J�)���*z�+QJ��|��t�)pr��D$r�(=Nt��)������3!F���-����u�c��ccﯽ�4aqO7�[�Аk^?��!��R>x��g���� E�z��Z��4.�"(�%WQ��ol�#����Q𑛦xhRS��qm�*�	���Ed�M���o��,�]{���j�z��f��� ��H]MM�^ǋM7���_6#g�^�T��؆��'�^�u��N�%�}AH��|�XY�"1��`ϭJ=t��w���?__�3��A���<5�^sd�Y/G~=�l�JƦ_k{<����/��:3y�n;:����§_�>9�j}c�ѧ��rbh�=�`���W��l�S�\u�8����f(�����څ���`�B���}b%�(�&��vjO#�Av�Hf=�ڡ�'��x���o��,�4Ϡ|z�+3���zE����*����mQ �HyW�鼋��K���[�4Ipo6,��(�.��z���p�"a�����q�����z_q�U�˶?#�z���j�'�y\��R8�]+F���F�?���k<㙧�=�r\.�G
w��W?�@G��A,�K3+4��c�{C8=DE�s��B���V�q��6��l�����Zw�4&@7J�D�v"w�P�^<�R�B3�4�SB�q��@F�9.�	����1"��>f��<��4ؖ?�Y<J7$ШmZ�]��4�4��+����f�j\Z��@�P���g9�Bԗ(q�kV�([r'R�>��q��~��A�o���QbCs�I�թr�ڶ�EB�]��k��M[�\b�#�.0������N`��\�,.bS}�U��@ˁ2��)&P��lo�R]�Y���.�Y��Q CbAE�6(h�aɥq��iJk�K�?k�T�s6d�s}�']=�����+��U�u�0�翅�շ����JW�h\���|�ؾ�.�(��6�d�ȡ����^�3M�S ��!��ҟ��#�N\b���\��R�L�^R�k�R��^���Cd����hN۴���s�U�o����6dM�eRJq��k��8_'��E1�̬�p���<Ǫc^�P3X����v�J��n!D�5&�b8�=��Y"�f�c� �6�T�)��nŇ"܁[�?�`B�E����n�7�#IN�qnS#�s�OSQnq$���8�Q��9��r4�Ȋ1����s5C�c�R�X������ ���4ɹ�`a�Xg��r�
lu�Ґ�nqD�y�tUb��A4��I�Ϗ�Ǟ�(e�x������6���d�T`�Xd�Z!��L�b'�)��B�J$20�ߧ�ڗ�����\f`%��C}6�A�Ru�=��ʋC�b��i�V�\,��(_jP߽=f��n ��ԡ��F��QU��>?�teoY�&�B��~�X�jdS�	�{�L%'���	~ ����z�(�F�\�w?"�eO{e�w��	�����W��2c��=wM���R�Ql&�1�^dp;@LG&]@&i	�¨�#=խ�;"��p`��-8����F�Z۾�Ta���<̴��JE�9��P]�y���\>҆cD'�c�r���E��[S5��l}������q��v�E�#���
��
WoO�H�q�ZK�ך���^|2���K�5F�����B��#0ی(NF��e�
U�Q.V��p�r ��d�U9^��Lp�*��~}^���N���mξ�U����b�Kź��j�ɸz�,�W�B~��])�y�l����3�����6q���J5-V6��t��/f�*�L�C�4��
7~�n�ng�j�"l}[HvSAJ�+�DL�F_ۋ��>HFӄ4`o�Y�Gp�6��r5G��B��k������j��������D��6+�f��z�(A6�{���U�I�e���E���}���%�S�D J���9�8e��!���fS�?�=�&��8�0��3��gNQx�b�d��e�?��K�Ȼ�n[�OG��D�-z��w�WQ��Wf����a�1u�	Bd �rU詗M�mzHG��xd
�=K�7w���^6���������"q�ɏ�$NK؞2@c��%���
�|��o|\EQ��#�UI_�wB�%}*6���2ԥr��rO���#|�/G�H��{j�?ﷸ�SZ��� ��zI����7�Jj�q���l��lA��6�4|k�t��G�����2�)A�f(1����7�����2&����Y�/�sq��7�%�v$��o�>I����.�'�f6��$K ��U$v�j�ǫ��ߥ";��L5�fY��L�"ƚ��,���M�Ċ�.�Yn���~�����?b	�o���"fu^,TX�͖�\��Uz�� ����<���+���;AwKp��p�p�i���t��f0 s���Y��q<�����C�eJ�*�h����)�i�7R���c�t�r;V�ҭ,T�y�0B��!���(,]�UW�����&S���mQ��=��S�[4�^� �Np�ِ7W���+�V����u8	/�]� Xg���r�P9���Z��S����4�]�̌HqSդ��0Rm�+ꛖ�k*܃�
{?�v���������C2@��o� �1��4_	�Cz���ݵ���֖�����B�(Mx����O6~Q�P�V,3M�� h����[Z9���E�A�uA�hm� �
�4G��|'Y&Y������l��'�+S(H�8�	��&,]��6��a�����FS���(�i	�%;�P�v��_��6��o{!��'U��Q��wn�����V��r��k���BƳ�Q�d�8�Ԓ�WbA;֑ԋ��a��e��v�0�g�V��Xr0x
:�N�G�%��2�e_��;CXJ�?��b�JJ�,�/��YŞ���~��Tێ��a;)�x����<[l~������m�/W�m�M�2����_R��_�Q�xf�iҏ�߁�&��o����W�t�q�#�	^��{0�j~��%e�JwdE����?�S(X�,X�񉊪1(�|R8��'��G�I �w�֡V�����u�$��
�`�������i����5!:���\݉��Za��7��JS>`��`2�����H��؜��p�mjEn�C�K�D�? bw���]��e����ּ��5=Ku�p�>�_�*�CeeeC�<<��u��ׯ���؂��'��dlӕ��9߿��0v	�������bg@ �=���/���{��yA;�3T�m(v�e3��4YcD�ʢ. h�x�����d��s����|뮰��j� ]z�0:����v��M���#�Җ���bYj3����ɰü�����o]�a�b���ܿ�;�����aj|��.	G�qP�+;�0���x�svqy�ِ`sQcι��'���Z�% &!!��S��Y8�д���&��>�n����60�'���0����A�Qp1f��\�o����uκ��JB��gwww�n���ђ��H1<���>J��?�~����17�YXK:�]Vt� c�ϗ��O�ښ��A*k#R��f�1����U� �^��?���c(���7���\"�$ֵ��h��Et^���0����0:z	d���_���AŹ���K�������eR^�V�s�[�B�>H�v���U��`c�9�M�3dw4��7E"��CZ��d�(q>Z}�8�C�#�q��Ή�H�B���[�N�+a�_kc㳣wB�ہ]��v3��n�i8p����=���֖n��?�K2AGzBp#�)��Z����O���j����.O���O�ffvg�홵���)�J�Z ��O��SPx�-~M��it9�k��r��y�u��֦�\rj�kqu-G��P���eK��,�8D=Q^��p*��\_�g��N��Yr�W�w�h(օ����.��2k��d����ӣщ��ܗ�ك�mϨ�G��������W�����o��)��f͓��ꏼ�W��td-���jgg�_����z����ؐ:Vn��2d�d}����2X1{l���#Jx�����_�vu�Ԗ��<C���5$;;{]`W��i!���(����&���\^& ��ڭ4./O&}Ă��I����~�A+ŧ5hMq�,ZLW�j�]j�a�nB�l��Ǐ��qv��=m�����q_��&�UOѴ%��R�t�m���.To���2ҿd�g��_I�(%Z�%�}���՗�)�w����֦��T	�N�9]ﰋ�]a����t3��iwz|�:����:��̔�Q��(z��~���L&���#�7�el�e�)֨�R��%-����B����o�S�V=�<���b�`H%zm���B����ݞ#�m[v�k�G��Z ��84
�f�:�$*��������8иڞ�@7����>a׹�W�הF�g�z�Ko
��j��$J-2}�/���S7��
g&���dg�g�(��R�S��%����4��s4���!����88��݆�c���p��o�Ћ�����Z6$�x$i�q�؟vTG�l]�%�(�{�徏����|t�ѹ���s��&;Ǣe�u�_�"�R���	M[[��Yf�(&�d��si}�d�)��+bOG�Ws�3[w(��aZ}m5�܌w\*V�-!:�Z" �c���éF��vȬf���'էW����\0����^�y��y
�M�<��G��I�b��v�D�%��m�
��?
j쇶�*CK�6b��oZ��D���v�H{)�Z1u:�8NBu��ߛbuK�����z��?����0�"<�֟_�>���c��e��FG8���B���DeN����w�� N2�|���2�|ENh�����K�C;� ��?;��$O~4��e�S��Og��j�B��56��.Xv���GLU+�5x����*O��m{h�F��e��D�v�d�G��n�"rps�N�v��o�ة�-f杦a5��(h��T�H>P�v���R$-�Ρ�Dn�8ԢA�;�Ϟ����	�j��j��{�֌����Txy�1bC+Z�|�B������aư@���I���k�bE��z�8��3�?�ĶaR�#�Qѐ(�X�
��1�C�@p�g�dO�qj�մ���b�N��:*��n�]�0�O��!U�]^�h4���w_Qǚ��lt	��A�,�u���c#/.dޯD�ol�|�|�	�H�=��ɤ��$-<`os�%�/]
w^W2���I��U���XI_�*�ޞr���g���[����4z�{�'���B7b1�:�4v�5���䚒�
M�ɆdG�Kf)	p��r	a�r����3|
n?��
Z)���q��a|m�j/�a�t�Z�GǽwBg�� ��_V��Ύ�}nKr(K��ݽUq��tc�~���~�����w�����1��_b�ܹz}�Y��?���Kbe�?a�\�6v9`M���<��.�r͆�\l�j�k�����.,"*� ��f�s�(�=!������;�/��B%\��
M��M��
M7*Ŧ�-�M�v������jXj�- J�S��-Ҟ��]��lX�;���"��%!I$9u(�IXv>"0���uFC�q��}��ͥ��}�L-��O���^�GFh�V���&��8���@�U�sH��d.�Ė����|2�=�m�twe���$��_{a�a����m����y�nԳ�_�9<t]!I'ݟ�Ym~W��ޅ�'X�<�g~���J2�%��ZԲ��_?�o�,�	��6Ucms$�a��k�U���(D��7�~��;ڠ��h���Qy�o�MW���A��zR������it�,YN_n��#��1n@��Ls��S��k���q[`��[�Y�	%,$&C"m��ǲ[��b"x��.�S#$���*�९��n��3��+'�-j���e*�-!��)bWn�/�rl63s󕂩�R���8y�Qf�"O9�=��Ak��c���*�H��~n����OS����Th�����\�n	k��ғ�V�h$3�i}��x2M��%�f&��u<z�7��L��?oDl8��B��c:��Q�df<�ާ��'+yZ���'*+r���,�zD����[D�����C=�+�o2��8����H/�y�e7��a�K|���
���K���J�3G~����Rh�~/+"Bn�W��i�_p0��mv{m����OM�^��{|��u����Ȩ�/��ғ�I�͂�b��>��_�c5?�{�ꌆ|��Nu�]սNbYJ��_��t-��"���Ѻ2��صGf�o�r�Y��

#!E[�F��C-v�������UG� 
�D��py�9&Clv����o�c��𥒓Q	g|��L�p�00*p�4Y�34(	�0��J����Y9�^2;��+��sѳ 1�ܷ�MPr�;]Hs�ܸ=;���}�4}��P�	Z�_�-��2.�Uԡ�#�K>'���x��}��>O�n�L&0�i�|�c��x��q)u��_Lt����;����t|�5�ϋB�x�md�~��Y�cQCw����Ҹ<݉��i�;��a��aw�]gHc�9tI@)�'S�d�.�+��燋XLIqZ8�Z���<x2N�jG��k��jV?-s68ei
����ca9<�	��Y@�w�rR��tt�7�+ُ �0���f�������|l�@P���7�:)N���!O�;�Z��7�J�AZ���[R#�L��Q ��R_s���Y�{�F���>ݦ�d��jۿ�n�묋�����#�N�9��Ts���f�򱀡F��>�e��̷�w����7���V���������%�؄�9�LC!Ś~Ut��e����������L��0l��_2:N�;��&���d&x�A���a�똢di	������yk�J1�P�e�v�p�R��U
�����4�T����^�yoUC�Q�(o��h�;�@y/.�����Ɔ����\
"��ͼV}9�7�nE��J*���Eq��g����v����!�������lE!����X/i;E���V&H ���F_�6J�VÞ�������_��%o��+�&w��<�X�(�J�<��'�"(�a�����j/d�ƞ�3Կѿ�r
D	W\*B�g�b��H�sf�="_��`�ݻy;1G2�Hp.ע+6j�[a��[SSV�Ii�ȼr2{X���Ka��|�l�õ��_�H�Ri|U�`�g��$�ŏzz�eJ�_�zn�`��
3P9.�3ƫ���G��o���(G�P�fR	ȯ���1�1��3�2��_B��4���lO;U)&�"��8�lL=d׽:��k�T[��RP�~�8��	���쑝��}���|��0�f�*]O�᷼Gt��c�cN}5� ��?B����;��D��z�]���f�.�$�7�a'�
lؓ���'Cz4�&�}' ��?��<H����K��t���(���^�F�`����(�Xƶ���I��jy�e5H��<���E�©m����-$lC�n�k;��g0��м����n�.a�f�PqABϷi89|�O`�/G^��'��%���c�-D9&�Y����	횈�)8�Ǚs��H*������Me�a�
��x�zz˽���k�2�m;�1���<��l���[��?�*���9hЫ��?��bЁES~��`��}�|�gC�l��2<��r�����#��Vr��P����kk���r2�|`/.i:�hn�C�e�yp~�.��Y�V#��4����ِ~���c9�j};.w�)o/��ʔ�U������������/&�6���x����Xw���Ib�'����m�v�C�?���������_d�]�Y��PM��~�f��������J������Q�vT�����G�Ȏ4fqH��$�}J�O("b|?Cȳfv��t�3��  i�|�Ʃ���5���n'�o�$�+��Ӡ	m6��FTT+Z� �_�1=��d�P��o��i6b��O��Pf�n���UD���lY�m_5`�>�üCm$l%�V8�٠�Iό�]	�K��^1E8��;�09b��~��I @@�ڹ2��Eo��������If���K��s�j̄	�������T�N4B�9��!5A���{��ų�I�Q��ɀs(�h�k$��_B��y0��W�q�����e�Ln�˒��.�lJʜ���OJ+�e)��R�5)���qq�F�cs�W�'|�:���S��6N���5P�[W���"�aCd������a&�
�k��� �i�.��N�� ��j
��[�,J�~J/�,�M4VJj~�-Za���E��ÍHQi�4L��Ty}sݽ��,�y��%�N~>��sw�	�exi���޲c�����&�]����W#`^C�"���ro�"�4���MxG6)�9l�er�@ ���OR���y���$Nv��0niMzƩ��wa���qE�D+�
1@ȅ"4��1��5(�s����v��IA|�����Xx��a���J�1������/�K|��ˍe��β�b���,O҃m%Cg�$}K�D��^S��(~�1�i��p�,���2���T[�Ƈ��l�M�yˈӄX2Vq��֏>�/ߠD6m���s�U4)�)�q{33�(��#�#�Gc��Z3U�W$�ʪ�s�4�2=��1�չ��ɕ�9�aF����'Z0,��޾�A'4��A�wڻ�`n�Ix_*�r��3!��ݙ��߇�>�8�X�^�^�غz)�<.~�.X5^�\�O�sAN��C��岂.YN���� �|��g�뛛��11�)�	�Jd�H���%�de�L�C�{�="q�5<��^�3R����s�# ծ"���E��K��W��Ȕв��u"~5Wj`�(���H�E�A�[�k�}]�������&�zVD�%�B���=!3�,YKÍd{G���$/);n��3�F���*�%���98w�p��&����a�(T��Ų�a`|�S3���ݕ��jaVkW	� �U�й�'+�~aX�f�"�O߮gm�>�:�����{V���P3��E�Z���=�H�d�x߫�[�<1��%�u��z�c)�N�[Z��8�ef�=`aG���9`v�&���S��K-K�b/�ԡ}����ph�a��!� 5~��Px��d!h5�M�Ma,E\_ ����s��9�Pm��SS �i�"	{|e��-�}Ze�o�W�����^m�us�kG��BV��P��f����P�]S��0�m>�o��������Y����uS�>F(J�L�=���6�:D�	��E���[��[��-.̙Jc�b��-�6Ħǣ:��}z\ yo��1�9/7 ji�+��t�"SX�]nh�t�4g���2K1����� 1@οɩ-�����\:	B��P��cܡ��H�0�Wb&޻V�a=^'d�Y	�e���F�v��k���M���54HּI�|yRL��.��R�_i�8ݤdZ��,zT�)T�Ѯ�.Ń���O}iT�Ѻ� !%��s�1�$x["�x�z���TmNc�Q��o�%��Va��$��T�����=#3�c��NL\r��a�l�P2NP����k�o��z��R14�&��'�T6xH6w�$m��jB�-�Z�4Z�� (hg�M��$�T"j�]X����@���o�_����}����t�RM�h�҈#@f^$/�N��-�PB3�1M̂X�4����;fPl\���n�_���S���N�g_��v0��kk�ڍ������
�T"�"Ⴣ�$,�B�>���2��G�^���b�5-�[I�>�����[52�?$Qz���L���v�P-�w� ���%�=t13d�#���i��K͝ZT im�pA$XQ�D���Ju�b���}$�|��_�e�5��A���]�@��}c�I���4�ڲ���gyY#ow����р1��sr芙վ��^��|}���W��I�D|�D��L��n�~I��G���j]hp��̨�&��ԫ�Y��\0Q��|ll�=�e������]8�Q��Rh+br9�i�b_�%��d֎J�Hev��Z�
��`��c�=�L:g�3�M�բ`'���CPSf0�sO��>(���<H���v�9o�ֱ�O����P�<�x��
�զ�iݪ�諹�u�~��Q���EBǕ4{��n]m�����|]������W��@L� �����F�8���$B0�E���Ç�/F`s�b��&+BH��\C��%��Rz�h[b��$d0��/���.��A��4��t5��f����Կ�$d�(�f��h�O4EZ�`bQ3+��`�-[���6:ڡ����D@l�.F3����˴��5-@Г�G�Q�DMa��yӷYQI~��f�=U��9uI���X@˯4Y��M�S��]] ����\��5��+0�a)�R���O#g"}�� ��A�����fȜRt �"���6֐s�V����j�΄^>�0u\���F��v�H�� 8���rK��\�2t�ܹs�, yO3gh=�;d~6%��岈�*~ �1PZag_�x�2%{d�x2/,��Og���ɥ��	pR�fǎ��w988�s���zZ��r/I?0~����u�`I�Hww����M����c� UX-eo�dx"��ַ�Ӗ�0R�5f�� Y C�Zh��Yg���zz�	�Y�\\��騀���ڢu��;J���Hr"�����Ӗ����)޻�x≇[c.[{��־��G'���
��#�����|P��Ԥk����	|SJ���x2���R;QhsW�ȑ�Q&�����w�Wl߾ǵ��ͩ5O{�?0ӡ�ۍ:MavvJ^�`5��� ����aL���Z �E�Z�]3a���j@���T}���s�h�j�$��$����F�/����?ӟL�)͋]�Ѷm[�Yt` �lWA�<G�u�!��Hƃ�x��&|��b�?$��T�$UZ����� )Ѫ���/�g���Tp_���7�Ԩۈ��N
�I@L�̈́6T%��*u ��$i���ua��V����� �۶�r�����;��h�$�&09yY���<��a���1��T_}0a�r�r���^���-�Ns05��pjjR����tD�j�c���h����E�b�'�����nW�j�6"w�d�'U��$=11���c g�GI4ͤ�>m���y2V)l�ۢ��BswJ��}��Hh�A�H�`Q�I�7�z1�a!w�rs�do/]u �6�q]�J4E����)௤����V����}�'�v�3dh��Νp� g��٣_"��:����bU�j�jM�Y��s(M���ȴ?�̛Zp`��	b.�'��:��B�s��zkـ�0�%��y�&�mф_ۧ>�ʮё;v�[/�d���1�ɒc
B��X
H���/i%�M���>��O�	��à�<k*Ʉ�Ivis+̏�K Z=� ԈTh%}�D7I�if�gl�wu��(B|�[��t`�G�fY��T�M��h���u��rQ��h�d�	���� �vx5�f=����F<�K#�]��� ���Q�z� H���M�	L�&`h{Q�>�9�����J\"Q��M��P���5���7���t:�k������Vk��W�]/�|g�稝�ߘ�Ӧ��G��*����3��Y��DM^�8'&�\�ZLYL*K�7S�������95u�m`�jC`��嫿KM�lN�_^^p��[��"����54ǒ��3,͚�<(�3�L�f��#��RM��֋����>�f�e�D"��<��q��LZ���o��5�����5aâ��k�oU�X�%���x7���G1�|S��&P�	�i����4�l��%-�#)TG��,e�o��g>��k�#��jZ��EwD@e�n�2K����:�i�@R��.���J��d��C��- ����MB_G6<�Q�զ��Z%G7X������b�;�L|���$g�4M7��'V���F��(3�ul�8���3�;y�	�FLo�#�"�o�z���:��ľ
5! ��U���	־�F���H�{�J�%�s�;;	��}��V��e]�K��[ܔ��rY��"fTw�|JOIZ�LB�>���}��爆~g �����r��Wϸ6�o64@�"�/����d.c(��(B�bR�ԍ�"$7m׮ݮ�"9P�4n���_Z Z?�� 5�"A��e���٣�G{:�\XXrfر1̰l�AW~���s��9v�s�>C�����x��233)`y&w��.��СC�4gE�W�l}7�����}�$� ? N�N;W ��W�����o�[��5j��4 ThK��+KimPD`���(�a���Z&�T5���E ꧼ	���iI� �_ʏ|�r��4h��'�):>�P`C�`�F�j��b �m,=`�wy����ۤyQ3����/%W���M�/�$>O5��c��~`>�iyl���$lLP�l��0�"h�H��/�D[�1�K�V��h����=�-͋p5���W�*C^��3��C�&�'�^K3�⺿Y~O�h�z0g�SS?O�ź�:S�/��G��1�O�t'sX�Kg�F�����bA����f����PpaeE����0�Ǽ�u}w����[�^>��`DP����S�k�Y�YN��yQ�4>JR`C�l�q��Pk���Xs,v�f1��n��ɬ�9�tV
�����94|��i��O�f��Q��::tSwtlv�SߥK睦k-� M4~(i���Q�j$�,�m���D��5�p��	)#6�j��ر]4��	3�"K�Ȁ�45�*�)�9����x�@��v��O��b��
��e���E�5a>���s|����N��4��U��d��Iu<]�ɔuD�D�EC�U��?RQ��=��;`�BsL��U�Q�'^[��4�Wi0��>����L%
n��74@�"9*r\�Ƈq�T�p&��*�{�7��d�f��a��ɩ"x �
&���=�<��ƊM����ی� ��˽N#�э���� �
����]*	�u��4�I4��v6�D����ȑ[�<Q�`b�����U�{Պ�b�^�N��~G�`�?Aa�B�?���P��`�f�9Pk�f��_'���6�����u�=���1K�7�ۻ͹h����o�X-�)�&S��9k�\5��GG/���h�TƱ~��?����}���i�Ke�����(' �S*��<yr�9w��g�e���ݦ�@���'��׉t�Ν����6Bi1�$��4��W2��%L���t���T);���b�0��?���x�{H�u���C�c���,�/h֍U5N-�G���Ϣ��&�G}���
� l���''Y+�崞��o��zJ��l�u���������c�Y��������,k�Ssd��Y�V �a��3IbAC�-(�5j�5�״v��?��7@�>H;�wT�}�`ji' #�=p���w�@-]�ZI������lr,zgi_�ݯ]W@Z����$*��Rz�l�g��ϸ� R4�qz��S��������*��O�H�(mj5��i/�I-2�c�U�H�$�����+��fi��fd0�� ���iI�0aԘ�z�@�S�6k�o���A�����4%�J�T���疨n���GV���8�����?T��]���P�� t�t�����$�V,Bx(�󇑥�J�0C�S��_��� -��"hp���}��9g؉#'놦� )�(;�ܽ�A���ڭw�uWN�3����_����(|R��}H
�k�h�3o��l��X��?�3s��ёK�.ly�ӟ!�k%��/}ə1�@e���J�Q��X�֘���+�x�ԅK]O�ۢ�L�����QZ��d�R~���C`.NUId:ԴXЎ#����7�2!,e3 �_���J+-�:�s�W��$��� ��ɱ�2��6�Z+p,g~�5O��J��p Xr D}�Ac "�/�`�Fh��L��y�iz��a3R�N�D�����0��O�)#�Q�8|��N�S����i��Њ=�hi�E��u�]�4V��\W4�|���[E(>-5[�/�|�k����Y���t�-?'�K�$�B���v����׾��|��@�9�y���S���3%�9C綮��Z��_C@,��@04��$
��?�"h��/-�i'6�r&��d6@�&^�I r�h��)��`�gћ��L���X�I�i����9]kyjR�/nn[�Ы��,p��IF�f����2B���a2 �y��	 vw�Sxj7k٥`���Dz���$M� Mxd�������@@�{������,�߰� IhC�3���ɕߠ��>}:���<ER�nt`y�}�����t{��׻TJ�i�����?�����G�$�#'O�А��Xw )=��	�b���I��� �� hÂ`�n��vg��d�g��o<���^r�N9	O���e2�<��4P&��k,|�J$G,|	���h���k�k�0��/�n���u�A*�W�M��h�\�Ԥ�
���`]W,��x��ƈB�s_��bp�2������o���T�9�����7B�F�jp�5�VϞh�j�'�H� t���T.�bm �@��(L�$yW��+1�M�~+k�nW�Q�1��#i���)@�^8���*r�w(��[*#�塇��"�ܚ��m��V(��>г��_�_?~�m'N?Q�n�߬�3��o����֙3'o�LO�9`NnB���8���Ǥ�#��姒�d��v��/�_�n̲��4�i�{�]b��$j����=D��>\-���Ԅ��9iZ5�	����|ںHhw��i�'ʃ{ռRMg��4���W�Wl-��߆��:�$����]/!��ߛ�f](ԯgi&��O���WI-��OӀu-ysg����*�	��O� }@���Lⴼ:w�l^h��/RE F̧���u�k�� ��6�@�C;��\����(g��g?ۙRY�Y���Q��F̪nM�䉩��hϞ=� ֒��s�����+>�ຍ�m[���l�[�^)���I����%�Di�R���;��-V/����g-6=�c��ǜO��H�Ql���&C*~��=B-!뽁�ΐ{f�Z5�c1o�B�ռ:$zШX�Ӏi����H��ѣH�'<T;GsGs2�4U�\tZ����C���Y�|C�Ԩf+%�oQ�Zn� ��z�@�͘v���k�s��YT�1%���_�\YN��F��H���w-����3n�q{��]t��<`CjB7�*NKܔ�W- i�u@㺒���E�`���άH+YscA�h�<��~����q~@_{���KN�k��+�����?g�w�~�V �f(`�W���+9A?&��#�Ƥ�(~�a�@��Ĝ ��#�֍̂C��4�FI��S�_�B�X+��q6 V���{�V(Yώ�fL  ���$H�j�~H��4��~!`�
�ˮ��z�A�$�{@LW׋T�ρ\�a^����gI��U��ſIQ�<������+͠�{¯�f2��H/(hcd"ډI ��}��9 �hdaʈ��|PN%���v����Z��L�X�'���g>�ldl�1��<�Gɉ���N�*y*�Q{F�5�!����6ձ�m�"�"��_�I{�<��0k�*�"��7�講n��i�H9��b֜��l,5ils>e(�(y�6��o���)���<ITv��pa��R����,�?KKtP��J9VZΛf�Y��
�#gј��z�MO�J2m���0��_�ԍby�S �[җV �F!xd�ac2=/� ��'i��AX_���.�/��	��(�Тx�>)�=��;����M?�8x
��w��xn�r@��G��������>�w�^'$p-^�S��s�/������Z�ъǷ,@
~��F_)R�uHDh�&�1a�� I�Dg9r�Iu�\6i,F$G$4��>��ϸk�u�r�W)�T��r�U�~�%M�!��A5�!��	-��W��1��j�:@�,��6��|��H�w�c��I rwȆs��i��O�/\.4@f��X� D�������	�0�9+�f�d��N*�S�;+IHa�$��A$>3�|5z�̴�~ȳ��~��NS�R�F�4x�{^����>�g��Z��� R@ί���oI��D`��k�`��RqPcJ��Z�F=Df�a�����/�u�@3#�A����~�R@Y8���K�Ij	Z����W��58����֏�dm-ϵY6�eW
��F=4�Z�Q�~a:7;�4'i2�dbM��%f�X�Y1e�@ڏn�3j���%���6Z����gJ��O�y�G@Uz�Y�9��13��DRr�����ڴb�D�1h�o����p~4�x�0�{�]��½���s�{����Y�X��@
a�0�W����	�
���L:y���̔�ԗ��(♏ƿ��:��P��i3E7r���O����q� �_��5�m�A��	V9�+E�-�<[��|5���M��y'�΁��CMۚ^�o�a�qlk��Q�Ո�D�l˝���.���(�w��Rih�i��M���,�1�xe��*�B�Њ�`��:�u%@�h�������s�!>F����E��6�8���OR:�J�5zfC�+E�����[��$�֟��?���Z��dޔ�	Q�!0@�KI�;��5�_����H�q�L�Fx0%�\�O-8���"�|:c�ّ��%4��nh��!(�(R��em���2���_��I�_��>��=ZMMԣ�(6�E��u�V6"BKO>"֪�T�T�jA7�:�M���g��x�͟��\S->��$}IO�?���,���}8��I]`M��_p��&���@4܃Ig�k�Y iڙ5�ϝ;�bh|���b0Zx&<�����V�N���V���Q\>���?��p��e�E��O��O����ZKky���B���� >Ɵ��N3�Z���e)8R�*"��c�� _-͆��Q$ ���i��ssZ Yja�{J;��kEnv��I$[��S�H�N��*���G�"�h0�h��O�<l2���2�̄��8����Ӱ&m)z��$V;/k���S=��k�8�S-h-_� 399��1n5�j��F]/'�p�y~��uʸ�R�h��C���R����Vmu����d.;�tR�4іg4n�aB��� �&���n�]I�@����h�����8�P��3	���������vѭk�b�%��e�\L
VkQͩ�|�3'4��|�LۺI�H@8�i3c%���_둪��a u!i�(���9����tŁ%�28�ŁS�T��.J��%s���Q��a�����E�Ĥ��l`�h�t�ot��ݛ�j���n�v9Χy� �z2�C�qK�P��>H�x�gE�z>o��ə��>̿g�Ҭ����[� �{R��������
��y�|�%)��R��� ˭��`ҡڵ���b�� 3�/��Ѡ�'���,��!�ˍ�h�3��
��4��Iw���O����T{��|§�o�؈v>��7���/��|W�7k�e5"�⿉��g幙�9ϭ:�i��8���I��������?��95tJ��Ģ���w&�t����g�F�Ѡ�b�ia:�g	3ț/�k�F��umC��,!ɒ1���9fh���Z��ϴ������qۨ��l�s[����"y�(����o�2��a�@&�L73�#=�j��4����S7f�kJ&�S[n��X"�������ί���i5�qfZm�����"�r-d������ꕸ���V��j]B�]p)��S�6�$Z�v��"Z�����jNůg�Mk�s��H����Ѷ\���� IJȥ��flVs'a���雾	!��o|���k�9� �,�3�1��D�n��F��H-G�8|�Y�hU����L���yp��g>�;~��st�# ���H���R��@�ާn|%��0�޵������o��܌�XW��\<�b��L�i��Zl�f-ʫ}^h96v^����.���	�PK�a�F�O�)�q�8���s�D�~��L6#����o<�B�'B�}�9#3�+��U�>W��cx�)&���z����i}�����jSD�FVHV>֮��_��*���������X·&m��{]����̣i��	�A���U�	� �3���9<u5�o�snkME�/x����?���=��>�� )*�"Q�y۶�� ��h�E����#1��*��#��9ʴ�&N�
�wz�4*�y�S���!�a�,�p~3W�t�x��{�E�n�2��
}�Oh�ڋi=]�����T%�Ae
6��k&@��4!�p�k�yy*ei?!���C�f��dlzVx݀�4a���>���H��}o�]�HFR��1�����K� �8�!�Dޣb������5H����Yc����g
B@�<)��g�-
�K.�Q�:�����D=lx���.����������MyH��w����Q�d�I7_�E���hZc���@ u�4G̪h��Ǳ��o1?Wf���3j釂'@��ϑ����IE;�X; ��]�5˞?Og�Agr���/��?�)��NʺcMb������䴘�.�4�<����N��߫E�uݔ��HR
 +�Ϯ�/:[˭�$Z�c�4��_�es�՛ZKk�66>lh*�h[:�T��7�v��Ҕ'����f�[Ws��1u����Z�D��Ə�э���8��7�W�)�.��G���ՎY��d��\EĐ`)r���C��l�5yަh�;v����ξ7uu����ق����l�=�T�K"�-��ਦ�1�sĬja��B�1Yz�LPL>�ng��g��$M�b2�	���\O��٩ \���,2���h�D���o��JR�Xc��ѬUg�	�N�tq �gxx�=an,� ����g�P��*��r5�dy-2)k:��6h�%��X�¯���� =�Qߢ�H�� �[��ct� F���,�k��Cx#�C#{-p,�!�������
�H��[����?�8s���KE�l���� %'iOGG�mڄ�CE�^�O�t�>�@�@��L?�����?߁@�����5Q�	�	}��I҉�!h�:]���$�gj���Z��}j�$ꦪf�	֮og���>�����'�Ngd�C"y^�@SKʩԻ>���}QLO��ÇotsH��G����!g Go��=��`�*���V��	q�5��4I�����O��( ��*&'ɽ�t]<4@��X �;����SkN�C�!O�-"�o۶ՙR�8�WU���U[��l�+�.;���6�M������B��Dֽf����#� |��/~��Zk]%G�p�����e1��k-/wHY��N�>|�P8@���.("b�l�dA���Be�
M�I�cR�}���dl�y_�RU��6�h	��HX^9���."ڴ���E�w��M���FR�EN2����B�=&�?j���nc3Ÿ1�QU�rN����Y�|�i�᳾��	�fe�X�tiM@��.Vw|�G�/F����w����#2]�4����ʣ��^M��(hS(��d�.F\s� Y�MoY(=��(�K���0~�J���,si����,.%,gk�Ø�ܗ�WJ��o@���f���n(@�T���k�tA&'^C�W�m�1���30B����Ӟ�4� �B��ڶ4���h&��+�!�th�C�vL��ư��j'��*�����NL�����TjU&��<h����I�D�D���S��@Y�l�s\h�К���w�'��̙�n�v�={���\��o|��j�ݚ����F]�M�F��Zz��9A3�kj�M�0A���|�R�R'��<���&�#��9ߴ�ڭ>�j��M����G3�K�&j|4�-��:pW��_)�@�9�=k��NU�{ߛ��������Re�ku�Z��P���}ƦM[K9͙���+��|�s"� UmO���Rj��j�g,Z�x�����^��b�+���O��]U�T�v<��4�������9��EÄaipOa�[t,��˱1���d?��h��w2j�]��v8��ر�1e���)a�;x�@���11e����<��A��k���v�g��I! h��F�IS�,�5��5E�'�3,���Ra�oO	��\v�H*�B��b��`% \UMqm�Wx#B>G��VKE�c���a�j��p-�\�`&������C�aY�l���#E�?+ɣ�u��G��ǥ�� �L��1�A1��������N�@i&��­vA*�n7�&�@�ل����~K-U���̃.�%ǐ	&@�m�!R��a�o�[z_I�c���F�0���]T4��E�3�/~�>'��۷��Qa��$�pn�6�59:4y��}a&G5}ZK6M����Ġ��K��1l�Z���S\G����h��T(��z�j:% ˂���}ocZ-a-ה����K��i!N#-D��"c����q�?y5��4�[_��W�����1�J�l�)���,;xz0���9��H>�I`k�`�X����X�q^czÛY�!*<�4D�uv�o�	2M�PJ4�po�lT-H@0�j��c��ǣ�aϜ�;�LH�	�jԥ�>>�C=e�==��~�{NMM�sZ|��e�(N0�v�c��젵z�ǹ<���>���%D[�Ym`^��B>mB���!A1
z�m/�q*T\~�a��{*�����iڡGk�j
O�6�ɶv�th>���ſ���T򊅊T����ګ���^]�k=�����q	�y݇>��k=O��o(@�"�W݀�ov��I���'?�M�Z�X 1�X�=���<dŒpZ�T�=��g�H~��M8�W��f��J�e��ЁI�s�wI�r-R���y|ʘ܆#V[�|@_�AlB�����$���z>&�)>ch�|��_t��G����G�f؃���#41}����M�M�b ��#i�T����S펵e�����xokP�5>"@5��
����A������HO[���T�>���;�Ѳ78/�d�"0"@��c*E��CM�z�i��4u��/�T�	+��ͪ���5��sS��Hk���`� �P�D��� �wU3��<�� )W{i������{��b��N�^
��C{Nv;I�6`�)(̈́��E�!y��dH��]c���N%oiu��]U����}%�vUW�\p�h��\^�:\���sN���XmM�j��Qz�!�k5o��:X �o��nQ���v��O�u1�j~�N,�[��#cU[}g^�13`X�5i�T0;��v���e�4�ˢ?���G��ɒ��`��PjL�@��b+jj9�y�ޕja�*�*���OC���sW��G�c�l��Z<�/�y��A $��UӼ(�PxA/��s�vN�Z>�-9�V[�k3n
�H��C�$��Z��ҵ
�r���W�b-.v�>����_�{�;���rP�j>�΢����$��R{�t:Gza&7�m�t@�j��,������LI�h��"բ�h��Gz�������W�	��5 e�Z���	HR� �فB�y[W�F�|���������z$�g�������*�誮h�T�eI���Z
0�,�A_<5*�����"hz���±��)��n�]͜�Z�ş���.�4�մ{͒5���P�>�>g¶��ɽ����Ռ��c�r����x��c%-�B�X�<�T�Z,��.� v��?�я���g',t�/}�K�R ���Ҳ�k��/'ZǮ/��=�f�d��8-���s(�D0f�f?X@l���nqZSc�A�x�
c�f�b`�`�IlR"��"�Z�����H��5p���w6��^3뽍-�t�_5d����y��<���YjI-"��9N[h��0s�c��w��}�_l�4�Z�̐�N�R}t.�����q@� ���G)�*��#d����
v~��櫟�긵S	O�#$h+7{j�g�	���|bcҦ]ߣ]�F����'[�}r�
ꪹ��L�cc]5/Ɓ��g:h@;y򤳰Yǎ�ZO����~���խE9O'��կ~5w�ĉ�_�B7/& X9�O~��|�����V��ȑ�����__��
I�!f��9��%/yIYI���cb +�x�>}�i{0v�l�S*D��#ͤ�5]m���d���u]1���~�J�����:����װ�`(�*�RS����1�TX�I���j��m�)��3;;�L�&�0�!�T�`֖M�$���Ɗj҃�����j�j
� b%)-�L��j���]��@��:�	{ƋJ�� U�%Mc�E�#S��	mSjo�Zxdd�����`���&6}o�8rͧ>��kV���1{<��ˁ�ޕa5�|��Ͻ�]�z�T8k��T�4 w���9?�r��d�Q�L>]��v�k�"�l]�2Z���o�Gٹ3g�&����D�vPȒ��i�H����-q���I�Go��7)s�ܦFi�� ji�n�&~ˉ�qi�s{KFXV��zH)k{��� ��)[Fz��]�vm��J��z�d� ���8����C�k!�&y��T����J�����)I��P�A��ὤM������<M��i�&h2�.�
�٢����Z
�����e���ʑ�Y����g��Q��vE��-ci*��CC&M%]f�4I�Z�����˿������_ճ3G ����+g�n� m�����]����׉Ic-A���>���4��&�c�`W��b,gC��ƪZ�J��w��8zM���#t�e=�� +$�i��_�(�'�[�陇�����E���E���&i�Dpjp~`5���N�,�\^?�j,@fi�Ob���{޴?�O{��8Y˦��S����7K���n=�ͭ)�i���"��(R���\=T�BSԠ7J�8�f�d�b�y/�tAD�ď��:��Fb����5i>o�f- �?��CN ��zhV5�?A��E�"�����]�gk$@�	@��� :RQg�|�۾����^��9��JB�~���B��s4�|衇���uCM�֨ YH�ߧA� �Fj>G[��D�x2ZG_߰�T���c��d�Jid=�2j��|�� դ�͝�TP�hD�"��e ���]��i���	�����^�K欪0��Uvzu]�{ֵbB���"V4��L�l�ip��x���1�:dQ�v��u?x3hv�J�%wsqt���� 
����"��O��w ������iyinU
$��6��� $�6;����0������X����>n메�=�;�"�������ws�l @��27w���ඁz�M�4�{�Vq�>�M.`�B���;���G����w�}n��\7\�y5�o���V��6���#e�M9�"d�V+��0.[�,����� FL!�[nyںH�vMU(w�-M�C������h�K�K3y+��i'����� w��2$ Pik�%}���;�?ٯ�74Ǫ����܎��girY��$4�-@�R!����%�!��=�I^X �]��S�s��K�@�W�k����.E�w���__��L
� F4]��\'[S!x��~�U�z��c��m@���unn���-�{�H�h/_>�{��-=$os@H���j[�(uR0Z�=�ܓ�6�- ����=�f��U-@Y��% :X��W��aFG���cs{F����ph��~�{̄���d��@G�~U��O��6ɉB����4UB߇e��4�1n�
障 L��k'��@��)>+���(HjpH���l�Z�������~�ou���]{�4-Z���\S�gY�!"NGݜ@����{�o����]ZjC�J�+L�D�8p�)L�9�U,cc� ,Pg�2v�3��| N���[(��5����|��[-/_���;��yJ �g5 ��h���܋^�gcg1�$�Q�����o/,���|��2Q0Bצ�=A�9h�5��_��:�L�c:tߛ��Yt)������@�^V���m���o����L`ѵ��ֻ֝	}�#��VW��L�� W����虚Y��{ �s��P
Y%�j����Q-�%���vH�߷��I-���W���PSk�S�=�]��Z����S�Ui>J}��9�M�Dk��0�� �ޙ��w�w&��<G��Y�zV���8�ڲi�Ѭ�9t~������xn�ch�q�ȝ�'��(�}{�K��h�ё��wL>j�%C7�8vN�4���(��W��3A=:�4�%���Zd%p�WX�A�>``�AZS�i�3�<�s�,ӷʱk�)��^��i� $�"x���� C-����<����VU�j�Z���]��>V��f��|� �`aJ���V+"!4�� U���4�(�����p4F��k\��F�̀3�0R9����W�O�[5�f~����<;�����n�<��տ�V��FV�i�rK,΋'$��	aT׺Ōd�TB�0�o��op�Y��U���!����W��|��I�C����Ν�R>�,*�;�0�$��	̀7$o:<�ߢZ}Eh�eːt���<��?������s��Ƃ��9��բ�b�*8�������F�|O�yl�oԛ���V��w�1����	���~�H�8�C�"���²z����厯tLҪ��#,hP��c%���sc���͜o��hۤ�a��ω�zTj�A��.�5�A�vn�Iy���z H���Q �D�: ڷ�Gh+������9-6jg�E��8�ߌ��h9p�ԏ�' >*��^� 5I^��Y�9�)��B
�a���$���ҎG#ǯj�k��5sժ-Z�`< p��9�,i(Y	�͠{<g���SM�	s��"{�OkǒE�z'���$�8��iXj&�<LcޡOy-4�J3k��%��P��x�S*�-u�Y���i�Z+�p4�GcEQ!���)�-��YZcx���������ۿ}m%:5���i}��)�v\�X�V냴��X�ӗ�N�7I����Q{�����ѣ.�������kn�&�tH�%�i�+�)*,^�v��]�Y�̪�J�'�%��Q�dT��p�t �!�wjj��QR�u׮k��o5k7��;�>z�$4�&�#�XM��|���-H{�Vy gb� ��/��m�D E�	�i&D� ���$�ROju���RUwZ�i'����c�/|N�"��+ ����P��X��E3�2L�ԓ&���"g�E㡡 |�������}��_~���i�A3��M]����16m�u��g}#5h�����A�z��]�L�L�֭[��� K;'�N=���z��&�)�o�,57,��hҖ�Y�tZ=�y0%0c@@
 >e0L�;�,��5UDxԴj�p�9�ͷ�b�*�Z��V�v
�u�Uo։d��-�y�f����8[�4����F��*���F5�Τ��;�0�v�i�g�_W2��{
���C z@��[���/��=��!��X�*��r��
@36�
�ȐGUH�q��w�R �U��܌���X#�A>!��4J�4 a�:��1Ǆ�%m�e�]�3����˄"�X�W5]=�6 D�eAQ2����N���4��W�}�J�f�MHTKo�Ѐ�Mh��enM$+]�u!j�?Z�8U��:��h-��8\"aJC=j�� � ��\g.,.ΥW��O���6\�Cpڞ��R�t�����6|�� ����B��-Y:�
�<��ŏ��V�X;�|$}���3���+hu݈� �Fk��#�\U
�jw�U3b,&�3�r�m�9-ր�|�i��2�?O�bZ��罬�����p�`h���	�Cy�n$@2v��-����&��,�cg,�{9��F��ت�U�w��'FP����!D�&�.â�l�t$a�IZ^�����c8�
[�"˃��>�jE�L�R�w��h�ߥ�<�[�1��y��gf��U#?d_]��Z!����'����5������\���Tb%�,W�4 ���z�2��
�����@��|J[�u:�0)L���'��}�5��s��9��W�-�a�V����P�Bx�!D���t��RU�)��|��4�:w�M�bo��k�I$ZB�fAȵ-L3��� ��O��}����y���|��*y"�����F��T���Ǉ��;L"~�f`<�+�ӧO��[�:^M*30��~�t��,��!���~�h�Z�rs�_��tC�Z����Y-�Z���#�j�|W��y�a;����$���!L��<�I�H��r�أ���p��N�ul�C��� m����2<���iC�n5ƻ�����|i���9�լ�҂a�;���4d��[�D�x֐�$zb&�� on!mV�<������ ��$1e:��1|C*]l��1Kk����aR��G��~��RntYn��*������j]nS����׀��ǔ�Tf=Ԑ��������N�ÎX"ɲH�a�e<]�D��ç@�LLT�,�������Xn�4NƋp߾띉Tè����5����aI�zt۷�ZI�y������Zo39kO}c����N��ӿ	[�%��.2�3h�u��l�6R('�#��[t�����BFcWO��<�_��U=�&�ýϱ��;��4xO��!{-!�LƖNҬ^������x j@� G��
��n�Ly+��:{_���t�u��������F�q��h��U4��+�K��}��*����|��ɇf�PZK��i�����3.L`⽙a�����ی�IKN���a�E�%��0���i�XH��%�r���>C�7�Y�4'��{@��A�bŬ87G��ט��R�K��  �6���,���*/���Rv-���(}�Z�LZK�巵���c����4�lW�L���p�4�d֙K��l
� �#|<X�,%#mi�8�:�1l(�;x 	036��\o�K�j���Ja��`���e�c�z�ė��h�H���c��[7gᬝ�oX@���T:���R�zx�D����I@��V�����f̒-L�mN{3�{��G��
�0{{�Zd��aY�O3F��Ω��`255!@I��|��'L�p���(䣧u�Uc�ߖ��+Q���t���Z�\�y�?v�@R��G͇�R�0�����0ܻw�{�2���	�q��ҿd�a4���,��L��6㡫�]����PS�gi��1Kk4�j�����-oy�b��J3hW�H.�}��������T ��ͽ��/r�|C����覨����&���PXTh��kfp?�D� ������"ArlF
�-0[�,b6����?�/Gi��Bd*�p��i�/巖K���2 ��\D@Å�ܵk�3�R���n�aYش
@�
�k3ë��ߦ��Y�%{ Ԩp���E�%`�f���h�Y�i��,�hfOhθ�o�g��N�.�$��zL�O�G��8C3j�����tУ���Y�jY��x�;~�mo{�[�f}�U
����_�4�;���� ����n/p��Uz��P��R���l��9��D� ��,$1&�%�"�k�L��t�F�P� ��1NL 읅ڪ��֭;��9�G��5k���y�M�/_��X�g�$�����( �ҩŤ���$ׯ�׸�]��ݤ��i��� 0 !��W,8���c��* $�Z[�� ��Q!tؘMʹ�= ��X�Xw�=�o����0�O��<�k��}���6�4F�D6��=y�x���4�4����PɄ��}�s�������j~Өc��dD����I���*V4j��y3߼y)���}��ҽ�� d��K(��$�J?���)��,L�D}��;6��[�m�d�ib�T+��4��2x�^SS��D{��g��*��-�Xu��y��S4�V;oat ���'\7Zf�G޿��]�,�"7���5^����z ����*����x�@��7�4-޳_ 
�0�
<fE��[�{�����fK�gcg�f25��+@��H�����1��똭;K�!-�/x�[�I��r�um�q)�f�|���������(k�1�*�s'���<�\[fv�Zy!m�z8��k_��'�=�Y�WCR���l�)�n������}�]����(�l�I�,��d3����ą �4i�HSz��h�t�6��%,��e3h�6��f8a��6)�Ԏ:����k�P4���1q4��hY�L��Y
V��`^�B������kj<<<��AW0d�m%�U\��Z�k�҃n�#h�qɽ��=m�x������Y��I�&Z �̃%��p3�@�fV{���k�X�x�oyEg�2�n���=�m�����0<6v)ZvO��Y���A�{�{X+j#��(״f�����Ѕ8	d-Y9��ʧf��?� ��/G�\�	� u��"�F�[ꔿ�}&�{�5�y�S�����һ��7 ���w��IAh�7	��7_'�1�.h����7PR����$�,�94���X_���x"�"���1}�J�>M�HC)�Yt3څR�-3� �'O�pLS�yffN6݌l�΅���z���u��Z��f�O���5�� $��8�d�-[T���S�S���� ��[����ڤW��yT���6�&�rU��g�R�nhh؁ah5�լu���|3~� D� ƞD����%C����O8��C3�b]���M7���{�S��Q=������~��z｟w��tV!�d߾=����i��Ga~�����o�������z�X�o
�2!���5�v�w�d�����f�C>�U�1����4��d(�d�L(-���cf�E*B�#2�M�{6�i-u K"����Y�k�l	6�:��jR,151M˜�#�k���O�*��9t9uu�i��q����wa�n���ϣ��ܛf��z6K#c~z�,��.��3� ����{�up��<�\��d�֛@�y�2�=��	�͹�<���3 d�`�iZ�����;��� Q]�96ˢ^�J@�\��!T����<�	�OU���^i[g��=DN����AGxd��Z�ǘEEǣ���?"��X�(�~�B~���h�;�;(��'��}��ѿ���xc�׮����ؾ��w���LM�6-�S�Sl�r/}鋅�4����ʀ�Q�M�i�_���i��Nz��f>� ��'��?��Nl�@as��-*��߀Ӻ4DL��25a6$ H��E	 }�>�.�Q�4dm��%���6C<����@���>�>ro��ɫ��_�FD����']q*#i�t!M����b���F��炽��3�SKM��}�Q��.��X��I�M�c�F4�4�t��	^f�I��e��~gk����y���0�u �IyH��0���Sp���~�h���Z
�p^��V�R�1�6�T�A�ߛ"�+|cjjR�Q��}��� ���B��b����'4e����߽�կ��z�Y��
�ٵ��[o;w���@�0������ot��<@��	A4K���J�X��d�+XL��6c���,D�E5�����X��e�V���3&�I��&mA֩����z����>�#� dE��C����*0�f�:4@/�6�&Ț�zuOh����$`��������I���װ{WB�?7ƫB�f��W�[�ks
z̯���<��E��t�N��ZU`�����	�9�0ͨx�-kY��u� y��m"_t|L��k�E����;�����A�;���?�G�n*�q��>�f�իy^[����y���+җ����܋^�b'Ak�:��������X
�Z�����q��R��17Fр9����}�7>Wـc��4�d��2q�4(f�Ts��jdN.v�Wa%��k ��'ѐ�`��c��T�I��$N��d�-���\��j�i���L�T
8S�ƨLY;«�m&�3g����5zѴ�ޚ�k��[@e�=�������U��˭�4F%��x��B�)E81q�'���ȈZ,_M��Iǯ5d�mj�p@��y�O�Ί��,�ߨ`���j�Ċ ��y�ݽ� x���Zh�Y��R��B��Z _������"0X.�5�m���T��*~3j#�:39M���?�P CL�� ��	X��m�cU�� �AhB����?#f�%���E)8������ܴV�j8@������=�q-n`yy&����=��iI�L��S\�^�N�e�ӗ����a�Ju��0��m�"2����&Z37X+!k���J7�ʘ��o����4�F5��1+ck���<�k�F������iaXL;��)O��4�����~}?�PRO�7M%l�dm�L��W�eQ�#y���Mj�t{�I���ӛ�YO�홙)�O}�ai��^��ۡPFf��͜�5�����«�.��d]Ͼ3�Iak)�y�&��Z?մ_���i����V�O8nTL�$
�8p�/!���p�x�88B�p-�c�_Ä��?���z�D��L�ȅ׿������ٵ����T��������iD^3���r����LiP4�~b���X�,��ڳx ���22�G`y��N�s�L2soBIks�L�:~ՄL[2�+߱��C�7s-�B�lv��L�fֲRX0A|_f�5_O(����͜�R��J�>&����Y����T�W����ӂ}��,������c�I�XkW���M��WkeڢV<������@�5L�V���,���&W��j���c��n�m��|�f}aO��?�F@?��?��8����}�3��E�vL�;w�v�3�v�vZ!���;���
tY-][����C��������w?���ʯ�Ҩ鏆�=�w��]~x��kF�=zj�>�)w�d�$'�ÛB	64�����$����i���;�[t�As	��8.��0�p>w�O�:���mWG�b�"<	�����ECӯ��p��/�kLD��+���5k����/|�\T0u1���-���-H"L��O�����څ��YK�r�g�WN�1Yֆ��H���4�4��gtz`%��kx�����׻������9�8e�H5ر���}����o��R'���t`�и���J�1�)"�~�;w~�+������z۶���ܹ�.L�H���({�l�=�9/t��\0��OR�v��CmҤt@��c����&:+�H��R;aʚ|{�Oir�H�î�)��D���'�����I@�{Q� f8�#e�Lm�dQ��G6'vOhRNo��@Z?D�2�)�/�W�+/09��p�	���ZU�t����ck mJU�b�|������$�=e{-��l^��?j�Pf��t#�����M��@y%���&+yv��ygQak��K��8�뮻1�ԧ>�Y�X�����m�`x�W8k
��g�G7~���{d-F԰���`�mzǖ-�w����
f���L��e����94�Ò�/\8'Z��r�	
�Rs����_��g���i�m���/��j�W��X�?�yjIm4����X%��yj6N�*<�9��uttJ��N�������Ǣ4z��	�h`ʫ>�{u'�<�y�Y���R�_��i�k�3�{��[/B��+M밧U������ B�m��}Ze�y��|�3� fiZ�����_M+ϤK-"P-�[����d����8���e�6�8m�ĒE���<���@����o�hjt3	>��Is��A2��|xhz���?z��e}e�CRG�"��v�BI�)�!��̕jnm�Ge�O$Ty� �1Z�7S���`Q�����j��	��.J�l�	!SS�+~�+����iz���4T}s�ZMG�g�[Бi�Z�'LIj�c�(�)ӾG0�̳i c^5�ÿ��ĉE	�!ः���%��`dsc%�H�2�Oւiu�5/����}��U�;����;�SL��:��u�]�\���]�L�w7��e=���7 E+�����/?��[��Bj�rZ����j�+�`�.�r�9�Q.\tg{���}˷��l���!:�jAl��ּ	�-�?��œ�35S�ƭ��Pa��B�&O��.��4+�,��������������\?Rh<o�;�5S��74S��$�(l�K	�����S�7�X]J��7�3�M�"8`�}�9�C�$he�x&��������]:f ��i���q��i����}́!�|�wI,�m���:ZQ�Ʋℴ�h
��Z��h
@J)�e���� ��4�.+���̌F*㵴�])PRK���K�/}�W[th�z��H�b>����D��/�X���)P-��͇�oB�>F0ٺ����b9��˛yϝ{�1J�w|���)�[���]5+�8a� �u�]_hdT�о�R��1a[Oinl��9�'.��j Ҏ	�bIg�I[��s��BQ�P˶��F��+)��u�iu��f�sl�!MB��|�a� �^# ��C|�Ø�뻾_�=7����j ���z��3��7@2%"-��,��I&B7~���ӤK���* ��KkY�4�����@�;���ܳ�u�h4\V�Z�1&�6~vʝ1��[��KZ
�^�P���̕Xh��r	�B���洌`���ͯ4^M���y�-���O}��Rw��ai!�	���i=�+�-fdh��A-kL��5�K��������g9�`-�'0�t��|�tuJ���z���5j)�A"��+�D �g��oX�b1 �pMM� �H�ww�~m۶}��b2���1�aZӊ����Y�y1�uy�w�q��;�^�����FK�W��:7����{�v�b̤�����H�;�����%�3�����#�E�q�\����I��Z��zL��f �`B-��ef���K)�K&�'5�b��ꚓLS�î��'�o"K{�����\0�����g���_Q������{���mc�+d{�9DB�l�_o,y�g�w!A6H�D��qa�_��G];�={�^�s���k�x⹯�D�L�u�@�X::n��ǜ��D��˗/J���y�Hd��L�͛W4���)0M>6�<M*,�@�]�����sw�(�Y��J���䆑�^���y_��Zi�M�t�T ��/�&x�%��~������4C-�r��ʊWn%
�p��$?�ON��jhhǐ��j$�aB==���3��]�xA�_�6��?�1@$θ�I�v=Wڄ��}��&I�|^iL{��Y6�[���ٓ.%u�_|��w���޽K��rUYH#�@!MA0����J4����Y�����i`A�2�#��V�}�9��2y�։�p�������%�w��t1m?Y@Q���dZiM���[�C��>���	�;%��>O�������q�8_�����-�PJj���g\��h[�Q5�� D#}���������DV>������n�F|h��4�ݻ���� ���FX�"g)���l��3�5�4��������D�8�@�c��ָ%��?����v{���zS5��֍��two�����/-r[3�H����C�/���b����?��&��h�K<���9�u>|����E��{䑯H龣��	Hnw KJ�YG*��X�/�a\���#���W�Y�1��-h���+�֊��_��C���A�T�?�*W���"�����
 %y��x���J�j�g���I�MJ�iK���X+
$�=4��&�&�s�D��ӧ��� ��_�z��,��~wG$x���H�u�
z8.�R�FX˱�s��0����jL�oW������>���|��4�/����#׻��Uaj��B�N�)��<և����;�~svv���C���t�ؾ}g,���_5�L{�Z2о8"�)׹ٹ�ot~̯|���^�G.��&=N�e�B�~O+n��xy��k����s�[4sm�&U�1:�MP�����Dk���B}�+��T���.�{�����N<����kE���y�7 5Y/�?������֬Sgs��Yc���8 0C&��<�����w�	�F�4ܤh_�Vڙ��oz���~h��|��^�_Ӭ�G�1�̿$���+��:M�H��n��P�.�dl�5�Vw*�L۪��cM ���.�=1q���yM�}�0��,k�s/��(`�s��{�i���	�ĉc�q&����{�ys�/�V��mu����w#��3��0�ҏ����L�ޓ_��}�7��/$y�`��}Aާ�99��7�R^�[��KD���֚]H�c��F^ߌ�V�:�)Ю;HP��;�r����gI�gr�y�kŔ�-�/r�{��ͷ$��٬@�$H��Ad*E�?��O��{_��� "s���]W`��ە+�Jk�X3��^zz�� 棟�v��Z�53]��KD
4�a�<.���o��$��e��ܧ>���n���/w�X����̃^y���E�i�W�����k���W��P�uO��$��
�[��6XK��I:��5�Ӎ�Qk|D
�/
��Rͩ�_���z��N|4�����~�_%��_�{��^�RM���@�����g�������,�6E���v�Q_���7��Ԩ1����w#��k����BFx��{Kw��OK��g42�&j���WC�|�ʃ��Y���O}P�Ӽ?����,�����L�Vo��`Z�V�Q���w���m�J��rZ�/>"�֭iļre���̬���?��QZ$ Y�|�՘�x�H��R��&�|�m��âݝ�}�C�J5�2ww��;�K��&�N>�q�d z���[�����/���ϥ��j���R8���)��R�o����u�ٰ�����K:���j4R�n��^_�:��w߽���ܿ���� ���Yj� h��4@�������s��=������z�͘�x�Z(��_,k������cp����?�!6���a��(���؈� �C���O�$�rs�~�gr����7�'�~W���[�==�]L}v'�� �oy�[�t�͒���B���H�xϭFźf��5�P���ua˖���󍘂5*1�x�H��S�4��?�9R��������⿑�o���ł·��J:(�9�����-��o�9���x��R��k�X�+e�����=sso-��ZB�^��J�H�֦ �<D��]�z�s����s��$��e�)��
�Ԃ�����\�%�M��=�qt�vWku�W �����?r�����u"Z���������[$�8��7�ɥlk�gj�nٲ�J��'>���?x]�%/y����[mB�x���y�koX+rTlۺ�����ݽ�=��Qsn$��ŋ�r?�C?�z@Ƽ����x�v� 6 �g?�a��%�+���|���5������ܛ������C�Gpl��� cEk�y��G��������]_\�۾�$7z���{����N�q}�Ҏ���j��� Gɻ��&�t���ɟ�����眹��o}�����8~����6���=`� Kȱc�~��o�?O[Kp��-�A2��۷�r��������2t�A��}�w�R�<5j��{�Ļ[T�쐖T�(����g?���w��B�6�ҳ/��*h�x
���q｟�����M�w���5���$��xq�+3�nz�r]Z�veo�$�3F
�
hQ�����2�����O�L�5�8��z��utĤLMM�������}��� G��2 ��։w-.ξ��y�w�P-�f�Q �ܴ��Y[�o�%;C�?��@|��_�p������o{�[��j���A��遁�WNM�}~``ۡZj�⿌�H�H����P�P./Gp�L�x�ZP�<ܙ��9����ǿ���~p��9J�_��y�?���F?88���ډ�����Q �N}q՝?)P-,JUru�����>��O<Z�o�}\�$7,��OH��k����5?��s��5�F'd�L<�S _��d���?U��5TH��q��}�}���7����z��ג ɠ%���'&F�"Z�k�����T���}��Q��ǨA��pu(�����G�O?��/��{�'����H*_�e�̙3Wv������g���?���K��h2�<��H(��b���%������4NNN<��w��}���'�3ή���J�$�3:zqt����#?�#�w7��E��פ�ք��q����R�G���H�����X;;���=g��FM�4<ZL�G�����~�_��ǎ��d�� �2�p߇w����.�֛��+KΎ=;��{�;�(ϟ'An�"�}�����^[)�vm(M�kC�{ ��TgΜ��W�r�����o��S[1�H�$/|b�Ύ��������O6s+�0==!y3t&�<ʩ�?���r�����ϒ~v�����BXٸ�)���S� 	��ƚ�~_������X�.K?��?~��7��?��v�� H�$�|��]?"��_����"q�,,�/^��234��K�y���I3؁ܩSgT�%�3��>�Y�Yo,A׮+4��)��,}�M!�9)J��-,,����|��_~�{����C_kwB�@�A�K҅�G��^.����+##{ϋ��f�9�*�\+�����n$�~􃹯~�>����op~���ݗl�j)`�t҉�j��1o����DK������������z�H[$��x�┼�uzz���[y��wS�H3����$���g���an�ʎw���Q����r۶�B���_�i�{��08�a1��f�m�X� 놠��G�������ϟ�����޶5�V�̶�R7t��C������\sӈh�Oڴ��勋]������_�B�;�.f�oȉY���h9֢��L��������۬6�~1�S�enn�2p�~�k_��ȇ~�����]��u��:u�q��c<�����vu~�h�O������zғ����r�v�s`�"����_���h&V�/��0_"���s�.��N�|����ԣ>���E[|������6�c�d8��N=xA�#O˭�z��?���X>i��=��[��{ғ������s(c����V��� 7����Tk�b2����L����{�]�)~I���bu[W��zfzC d
,/������'}avv��K��~�y�}�}:���|C�[�$@9(]�7��E&Rϲ��iu
�)Q�>�8�UP�
�[Z���쬳�MMM�~����>�����������{Ξ=�n����q����G����������ѩgNO��>��}�#��9rK��n�����;����z���,���֣ &V�AF�l���D "�î.��t:�5==�{��'%�T�S����PG(�������mccc������� �RYH�R��e�9�i�##ù��15<$�����vi*�C>ߞ�������=���*u�O/2���5���J$��d\��6�a���L�|Ls��eIo�
�������;wQ�]�2�T��{�ǝ�>,|��v#Ú�wC����vx����.pabb�I]����?rnnZL��t�A����l8w�MO�]{�MR�uH*����g�S��F��&+7^dU�>�U�oM~lڠ�'%gŹ|�;�gggD�$y���>��O�p� �/��8%e�6;-��Ѿ}�\B?�c^r��$�����膈H�g�64@
�����C+�8�2O��͑�����i� �����?�,�םb��V����Z�W(��kS�|�b�Y��7ͧ��b��t�O�j��F�C� � �>}����I�v.w��Iy976vQ̧S�>$��f�ܲ��� r}ΧMV_���C�rǎ����m�c6<@ʂ�eAbjR��]h���?��JAS��w�3�vy_���?+��Hn``D�씴���={�v��#f���"�˨en������bm�1m�Q�6���M��9�3���g� �xA��/8��9����ҙ���]z�4�+	yN�j�߻,J��6�����P��~d�<j�]Jp�e�+X*8�chh8܊�5.��wV�����^m�K�6�o�!�h��`2ѧ]GM���	�����}�������c*S���4����ю7��$����g>�ɂitrrJ4?�ɉ���X�����s�֭����L�0l�~o��4��]�'�L�;ڸGlh��EsF|�	(>ue�k�y�1 I�P
�u7�ϱ����0o�?�{챇����988,|���n1���j�%H����O|��Հ �ی���ݨ��sֳ�{�u6C5iz����8���4J���sڡ�Q8MP��N�}@���߽��5��
�_�<!~�1��v�8p��H�ű������M��o�٪�n74@Jt��Ν;�J�Sa�Z�	`�f6X�@��uЅW��q�/..���E����]�����@��-��	��?�Z�[�
�1@��-��~S�y��	1�]r�*��j�k(�B���.�^;X��Ѩ��T���r����	jF}��g��w��%-��s�3:[�u�^F8~���%�a�ԑ�3Sc�j��� 9#c|��Z��߭����u񋁁��-[��������{�������3TWL�:�A:j���,V;*������h�yL8ܩ����.�m��<w�'%��8�S��m�t�7�iF�M������ut�y�?:����[k۷�@��b��.�Ɵ-�2��֙�,��w�i_��(�C�=%� ��~��QL��N �\B���� �t*\ T0�"
���.��R�;v�p�4�9rD�-E�ء@�n�}'������톚�:nv�$4۽{���g�Ȃ�6P�G�9� h�12Ѥ_S�'��Y�� H���S-�[�qn-�I6ꔓ�^�3-���y�X�ݗ{���= �������׽�?�3���d�ou쥖����N�?.@xA���$a��D<��Ҙ�4 ��'��-������'?�N��9����j)Z� � 7K`866*Q�GE�;��ZzZ��#��L5Ws.�V��Q���#;F�7O��e����8�1�j���0�s�5�\#q�eAR��|3���'n~�'�%R|��@�<i����k��Y[i_c:�L�5D�ҟ���{6)aܘaff�]-�M�6; ��T��hڠ^S?�ڪ�Osr�IW9�o�N�h��h�<+�~�c�|�PUpr�P��O6( �s���=H���� A�Ć��;���gN�z��}�'\#UmI�ss35yZ�Bv�������gC	��8ZTk�F��M�|���u��Y�H���,:4�E�qMPPA�'?�'���h��!�czz��&��q����"L�j�R,^���X��x�X�~�����]���n׌ ��޽{�.��w�"�� �X{��������ذ����Ȇ��������ߍNM�����5�!��qj.�U�&W3����g�h�\��]�ҥn��^��<�V�%������i�k��&ǂ�M��D�m�m��5^��i(&<��)�t<��O���2���G\�o��5�P����Me�`b������["'�8s>�K@�����H��8����V�������FzJ:֗��������������ݶm�[ӺG�s���)���[�����y8/�!��%�}��Q����%�[�bz=q,@���{�L�!��I~'ǿ���ď^���n׍ ̘,�a6����+Q������dxl1 f����m��ivaaI6B�3�X�j!u�&-w�4�@}������XÇ���q{�E�s�|�6���v�4M4S^������BO��x d4S�7�ߧ����Ly�&_�'<4�����EC<�4��ѳ�{��������]��a:�OJs�Mqn\ol��8p(w�78��Ν�\"�E���K1�yӯ��%��y���w�	 �'A0�ϟs�@��h�ҒI"Ǐ�Fx9��_r`�k��μoU�p?����{Mb� i+�f,��snl�Uʻ9������F�����B�E��ށk5 	�
����O~�{����x#@��/���|@�w�m�ZZ�1	��̯��~���鰪>�YN�<���� %�0����Y��iVǙ��b �67k!d~�F��㓞���2O�<lZ$h�Ja��ozLyh5<K�����w���-�����y�)6&�g�|�߫��j�v�l��ڐs����c�2�E׍���K�U������.Go����_
8U8R0�|���;v	��q��h?�by?2B6e����%B#�}cm �,�z��|��/�i|������G������1�p:tح!?Z�=+����N�d(X�RΟ��O��A����U��K�]Ǒ��A�ճgϺ@ �i��>����ѣP�B��T�HG�={�<]��O$�mh?�"��˃H6hfi�
f�o ���gi�̛F�
S�Q�'��%`&"K��:��/՛e�ׯ ����Ο?#=�^$���/d�Čю9�e�5#�]�c����AF��ͽj�Xէ:����ͨ�44��I.T8(XB��� f\��%�N�6t���&M��>�� 1����/|�KN a���2Y��qG���
+I&_jc��9��y���� X���7Z&�ef��&��΅�jZ��'ǢE�pĳ�iD�Ν�?�@4��~9S���4���ZKOi ���n��}�S�X4[h�|�ڵ�i�D�Z�k���z@�@"L��S��ru��^�����'{챿��v
D�����������'&�k��lh�T�A.��R���<�<�'�(K$j�sP3&I�>�G�f�B�d5 Y�2�uo�kz���  =�*�z䑯��O3��� /�'�F�ը���WK���iRͅ��}�0s�A(JJ�Y�����O���	�����|��
ѓsN�@�!��ر���@�]7��(��W���ڲ���l���������{�.�7�^L�0`� ӨP���+��S4J|�Z�Ů�_�����b�M)�_imV�R�-����j4H޸s������0�i
(Z-�Z�E7CU���;fm �('����kY����G���R-,>�@�2T?�5b��l�o&�M�{����e��;�$��+�I$i�4m�u�*&Ym�J�X՚�X�DiZ�j:��h�.���v�ӊ4�zb���NI2�:.�v���<F��,�fl윘w8��|��NK%�IC��ħO�_P+��q���@�͛{]�����K-/�fhh��!�a}`�C"��j��cr>}�D�����[G�I{�v���]7��g�O��l��TY+��Y��*��RAM飁O�.�3��w����nU�IעO�I��Uc�;,er�]m����z��ɯ}�k�3���W�wJ��U����4�_����Y0��Λ���rIMNCx�R�h�g m�;��t�FeS�@�T�>@̐jƴ�0��<s�_��,�M�.��,6�VA�5=Di��*����r=t���$���BǥB���,�ѴE5ڢ�`�X�)UF�=t�T)]G�Gq}T/�k�z�R��U�s?���SBɩ����ԍHn
��HS��3�\
 :@ſbE��|�ŋ���L�(���d��@��a~\L��$�}� ��&$Z���\��Bj!�s������q~O�����	O7�g(!�+�^��-�����u��0_���Ν��I��.��4�DsQ�i4<a�!���Γf��j��2?����aA�H�(4�j~T�e:��B3g����,m mzt3��Nz���K��_��4E.��(��G���Z�ֺ(ԡ���3s58������\j�� 5�ͬZ�&����{�Ѵ�WH@�$�V���m7�c�d�*	)U'��{Dr�)���K��]��h���U䤥L���8�wJe��B�-pN3�mrc<t���)���kI�ƕ�v�&Z|t����Τ���$e��I����UE	��2@�UK�b����ٱm������[  ����ӓys��5��[&"��HS�D3��5�j̧�^.�	�`[
h�{Y� c��I� ^�]"Y�4�|%ʹ�D_�'� Y�ˢ�M@Ej�v8�Q������	x\r塴����O_ � W��MJ��`i�Q��IϦ-2n��h��g��ɚhY�ɓ�
��Z�n���^	����h�	K��-�H�A�:���j40
!�ۯ[�R0�|\-G��u�0���%0��գ��h�hA_ "���6���I��m���o�����@�*�'	�{düD �?�F{:��@�0u�.��A� �o ��'�Ɂ%��4Ŗ�G&5ɴ�6�\��(5����,ɚ�-|���1�$[��U��j�֌����y���5�>TA�;d=�[��n8! �Oք9��HԶ�6��?`�y�ԓ��T�t� E��d�p;ҥi���5�U2}��[����l�z�3�Zu��9�0�c�1��q`o���a9����x���z��>���|�Ә��\f�d������}� �n[�,P ��}37"�iq�N*Z���s]80�}v�4�j5Τ97�N��H�T�0	9L; �Ls	ܱ~t-�)R��|`����멹i����ã��/A:7��
�mZ�H����gb��k96{�.��#tM�5c�U��XH�����K���Z��
���ض��I��v��a�P59�_�ޏ[�Z�՜Y��Հ@���$��	��;R�FF��oZ�fɽ#�}����?"B}�d]"G��Dk�UJC�o�p�d���"$��\C[� {�V�v�nSOLLK���n�b��H93l(���W�~�de=Js���itN�=�"�������=��P���X�Ո5�߂P���dT��(��F��P��.)������_�"��=F����''a�t�)1�
毕�X�t��5�Յ]��°���M�IPN�+hU��U�٢������&(bF�jA���=�3��9��˵��4%0�����?)��?)��?i��7ҹ"@f̶�l�!�7�&������� �Q%TeV'uqqN5\���h��0O��1�h~�V�B�J����*XD*����0è��zCvJ��AWuƊ��T���Ү��%Q~id߫�~�f��ѫZ��u{&Z�iFy��p�����/�*���5�ӂ�L��f��<P<@h�Ϻg�ޤ+.����CNĪ�-�|�J(��g�����SN�*��d��S��7�r��dJ#B���a~����zC�o������i����Z\=,�o��o�]];��5E3Y��(�z)U+��f�ū��sA��t91�WJ�v������8̰H��9��8��.�V�ђ\V2
-��L�z^���6�X�����#�k3վ���/��c_s���c�06��;]�;������X+�"X+UmڿE6��ͭ
'Y�B-��A�j8�jex5�',kh�4�m���l��5��k[=�k�z���in���F�������=�Z���A�m�@ �D�;z[������h�, DüL~%��uT��GG/l�Hm+���YDs�%Yl�F�zSHXi�3��gK�J�
��g���5)��T0)=?ץ��1b̆
.�ߤ~��^�|��
k�6`ml�S0ohO/��9�*� VS��9��@�Z�!/��V��?��7�yk�����da�����A�
�A�z�V�ϴ;�Z�h�y0�C�.�?7�M���[p����b= �g_��,;�c��� 9?p !{��%h~&{����i��6�ҵ#4#� 	�Y�-�t�MA>D��*���_/�ڬ��:2�dA��,�?H�RC_A���G��2}�|���]I<�rfH�f��>���,,�:�u�5��tS�C[^����2n< ���jo^�p�	3CC�¸�{�䪫 ��iR@I�^�[n���d��K���U�!�J��֢7?V���c��5 �PSLC>`�R+���']}VM��]��-hO�����c��LK.�F��G}��]���i���r��^������9���&�ɋ�����eH�k�g���HٛC��J��h��%�r.��	��;X,P3 �"�0�j�+>CmК���L
PZ���AZm=���7��8ۡ�����"��]�_���|i�� S�l2�%i\Mk��|��a5W�>f�ѭ�_;�����@o�1�o��Xr�������U�IR���'��@v� ��"�Q3�r-iO�>G�,�|Nz �>��a0�ڟ���Yv�ѳ��η�R$�>1��O�7fi�j�&(M"E��8�~�� i@j�W�k����*#U��>T�SI���sLh[��p���>���ޠ̅���J�W�%�f�1=B�)S�u;��ɜ��j���fs5 ����7P��	�6e��h��f��ҙw��2Ѻ�a�����F8F �h��Le�������� ��w�S@rEȹ�z���݃]?H�$�'���Ǐ�b��K����,��&&��T�[��U�S�/�le`EP9��Ij�c��?-�[ ���t�������X����<�J���ر�i�
�)�jn�����^�`�Dà����V�e��߫�g��F�������!M� ��3�25xfzZ��h�J޽a ����Cͧ�X7�N�-������I��]��[-�����%Ì�u���.en͛p�&~�{+Qy#��RV�l�{E���M%I6�U�I��Iv�W!Nr4I3�V�~�%}��|��H��!
slqD��lyqIZ���61�����,���M�{7�f9>>�J�a&�I��E�E+��W�Yӥ����5�f�m}��sƵc�jΡ��
h��X���x> E��F�������	�ޘa��E�z��gIg�=��ɽX�r�/����� �F-<�}?��K�_U���b�F�������!�A��д�r I���_J�L����]�>1��h���0�Y�5�Յk`jAh�T���lv�RQ���B����3�ϣ�෺,�؋�rh�٬Zy��� i���S:���SL�C�ʓt
�I�*�w�-��q��b��螝�G�/�&0�/;���๕�cn�4i�o��V`� RL��\��Yv�8�C���w��M�������C=t��a>��տ>θ���:���XS�2���VQ�C�C��q��U�L͝�<l�l�Dg�=���q�iH��}��߃�<
(p�ƽtiT�}']�$y{�bK�G����g��7�(��U�9M����僎q�>�x���N�ؽ��J��57���?mm�@g�Ԭ�4Z�v��$�2D�CS�j���uU�.�XJ����X~oe���/������4T'5Y�J��V����r�����|Gz|�fV5:M����z���~6	��]\� �,]���e�Ldq�}ֆ��8Ց'''��B�M�g)��k���{v��J����I0�s�a&پ�A�?9s����^�T�pfXL��K	s��i�Mi
��!�~�o|�c�cc�s'N�qш��o���5��n�-�?M]�Q1�g5Yy�D�P��J�79��^#AUPԊ<Z�f�f��C�[��jiXq4�}��^1kT���0�J�`m�ʚ_+��w��с����0N!�ƥ�ChO�C|����HY�'���d2o͛V�)�����ai=����ؼ�m5�� ��-��6�h8e �a���g�i{ffV~;�I4��2V����eX9h�i2k�)L�dM�ܹ�E$�k9;;����r��8RG���{}#�X.(����L������e���0�,��@PK�-�͐hK���@3Kr��m����p���*���[��O�r "��8�-�T+k��F��0Ȧ13����W)C��D�u��|�~WJ���?.�ǫ��Y6�R*T�	`<*�>�%�\�0b��Yl�5���V���V=n��ͼk��^uA[�coΝ� �Y2����U�P���d���n�xt��"^�^a0�-N�Ԣ�
�JO��ηiT���̄k�s����A ���Gd޲�W��B?Whf�7-H�V���55	�N[Q) j��jw��3�P�¢��5j�w�}���V��2���\� �n�<)�Hՠ>D[�����C��ǜԭaw��������'�=M�>H��g���J:�#���7�$�y�{ 	��]I��f��v>��H&N�"��H��H���If�����;i��ϔ��dV���|� ���I(<�J����Ώ�ƏY��f�d3榁���qލ�-s,�XL~ (	�!T���yk\ݱ�ֆ˗�$��KE����R�R(��t>U������͊�{��єY H����r��ym��L�~r������u�_-0�Z�&hch���Џ��GS�m.`�i=��w �� ������e���Y��'�(�d5FW�>��}�+qE��n >vuWzk_}��4�!��>�}����@eS��4`f�d� �߫���&�z?��\Cԫ�u�׭]�4������a����ԅ��+��lP����I��	��}4mk/�v](ܨ���E��9�z0:z�&�b��,�I27^31�Ŀ3��L���-,��k���B`�YRkj����4^���i�9C|��c%
����i�p���L�ӡL;,��{�h�4Z��R�Gz7:A��G�Iάkǐ����;0G���wܻ\�y䑟n�\��3mx�dZ��s�H�'��Z6LC�O�9+������l3[  �c|��c�]]h��h]C�sT2�V���k��d�I�浃;>$�'�I:�_/y[��>�J��*���}����B0�I���4�z�V�ǂ@B���U�R�V��k���X͡���_N�� <��4-34�B���,H���Q� ��������� >*� 8p��tX����;㳒r�E4K�7}L)�j���h�_�J:w]�p�VC�Q� ��ٵk�sD
�k�X���8#UmZc,C�4��~J�R�wL;�����G� �k�I3��<�or��M~�ȭE5�R`�s��tn $-��D#����
���3�+YH�8zM6�.�?�c��[�`��<��4�� ��h�Ⴤ�]����3m�4:�5�z5H� ����p����w�$�Q����ǥg"̓�'���S(`�o���p<�ie
D�h$��+ �۷�FJ�G�Zc��>!��{�䚮1�|�D��@@�2SSc"e�.�-��4��5�� �]�|)w��wl �̊`�U�z��u-c��M��j�<Ck���!3�V�*���b�u�BSd�7�YJ��h���|�Fhj�pR� ?������̟��O6���۲�ե}sn��k4@z�X-/�_ɳg�9P$W�
	�������[�E�$x�:��+�[�X��8!��g	��_���GZ( �3��$i�&-6`V�MeͰ ��Ϧ\Џ�T�܄FAAl*�P��z��N{��e�.j�vK� �u�����@��cc�҃�)� ��N��,"�"4��&�|�d��i��OhL:9׫ۂz����䙽���"�]�Y�AŊi�~�f�$ ��h='����^U��ڛ/��{Qڸ�j�A���Y���Q����$fS�sM\�Bث�g<�4>�5F��K}�8�ɓ'��݊di���|בɥ|���GW��6֯��1��$�/���3���>J5����i�C��j��) K�ø�~�_�MG���țf�L�,.^<��喧�K��9��_tA1z�IHD���1s��+UX��M)�`�7�3ױ�(�PP��m
t��u�P��` <R �g�jq�g�{��Y�߅�UA8��U�ZI3^{�L,��Hi�N��V(�tuQA[����w���K·��������ծ��7zEJ:�qÿ��V� K�Pl�C���T�X�6o�J�8�tg��Y�����T�0-�G�-�h�T��`�c�/W8�z5H����[o}Zō��e��g N�:&�0-*���4�d41���aʄ�W+���w�(D���6�
V>���9�j�9�:��҂��$i]�x�i=����^/����>�?�K%P�ǆ����J�j.@*mt�X�4�J�����}#$HC��*�Sm?�y��G9գMΘ\1���q.��*k��?-����v���E��0�"��Ha�$ ���>i>;�1�j�����e�4K�\s�ȵ�t�`y�F�}Z�S�/��o>	��M�� anG�> H�I���Sjs>I?�xT@��=`��`�x:-"���b��ªȟ?{�f�X�ҋ<��&5�j�Vfؚ�	l��ب��)iOں�hR͟LV���)�u�M�z@Ж�wBe�R}BRE~G��!͑gk��x�R`C���f�����N�&_%���4JM�WFW��X Ki���d���f����`2E��x��$@@�EE���r>]�3_SR7�Cu2�^��c��sk���	��Mc~�%`��(������XZ��Y���h1��`,�v���D�4h�c��~�6/gѢ�16��|f}�����L�h�K[�ly������U�]����	��*����H��?{�̵���kgFF�@SA/`�e0&���9n��S�^S�����k�K-F���t�n?�4�Зd���s:��
2��!ՙ
��6�`CӱFk䫥��/$J|l좳�X���Ȱ�ַ9"��=�� �_����V�,7Y�o�������U�yQ��52��H��7Ԅ7�f#@�@X����o�y��$�؄M�v#�LD)j��4 ��1��T88z�В��ja��� ���M��k�@���%�Ǥ����D!���-�5�W!����B���W�P3�^�K�KVM�3a�}��Y@��HY�33S�d|~C#��;@M���VM~b� XI�5}�rxbR��c��+�<.���x����@�*�,��DZ�f�l/��a��k�˱�K����Nc���9� W9'mF-�+%1�3J1PI֏@�>�05�X*� ��fyh��%'��$Bri��$��I�+�\%��a�5Q ۟�ʴ'$��dm�:��	|���@���|�j��@{2I�\�E-օ�j��-rML�b�A~s�������G?UL��#��qI+��TMD�Q d�E!��C�Y����v3�ht��أ9���ԜHvD��wMpY�hlj��H	z�͟�,pL�~q�1�8=S a*�DL.�uc��D�>4��ߛF�u�n' h��nZ�:>"��@����ou�ڱDh[}֬���Gx!����|�^�[�9������um���6r$�JQ���Q��4�G- iZ"�7W����/o�ry�D ���ro�|h3Uy�_���R���r��O�:A��řq\�2����Ĕ�ZY�7��8|h �G��&�C�N����w"�B���2�}�&����r���6Kh�IM����[�LE��A�;)f�S������9�/L��U���8�E����*�`��4��bK+]����iw�.������Ӛ"���}����D�^Ta�aJ����]N��f���)� \��F+�Q�S�����>�5�ұ=nB7��w'�E��)�}��~���i�h潭�s��0�Uϙ��{�l�f#�R��e���U]���[�_��;\;+@�Z��n�u%���&�ŃMk�� ���|����q�[w�����;����~��x��o_�'y�>��%����-y��c��>|�b��eK�m$i��]Z>�	^�P#�y�Y�}���L�t�F�����0D�b����1�O: ��O�#��C�&0�kg���UH?��iRl������$���e���v�c*�f�����X҂1�� ˾G}�*A_��ء�  �����
̃T�9/|�G�_�ޚN�AL�H�1K엍�&Y��D�S��M�ѡ�)�&I�����:mL�>j�ť�Y�re�� 	bJ2����ƪ������x��x����>��̻\��X#X�Ğ�^�����I��������y�j��^-�,� ˺	Ǖx4=k�������e��:�`�>n��-CY�X#�PBB���LFJ�I�r���	��ׁQU,��̭՘N���[�x�i�Vr,']��~&@p�֮K�}� ػw��֗�0���U@���r)C�K���#��'��������d@1�^/��oeAމ�?m�	ͫ��ff�)@*)��r�Vݠ�1��j���C ̂3���F��N�!.ѲZ�>���f�9wN���34��1"�����̠�������'\�h�	�֮5Y��^
 ����{�����4������ӡ���:�����m�z3��c_qGה�ZOJ+?�%H��YJc]��d�E��X^3L�muZ����jv�ր@KDj�2��^�ڵ��dr*�K0���_&��p���5�L`���%��c�����*�j?/��߭������5 �]��eQ�eR��N���Wh]� �ۄ��)��@��:-?��D�&A� b��̛�69�$-U�V-PN�U�I�_T�^=枸��S�S��T��ŀ�[����>��rO�`���L4b�7��Ӧ����,P�`z=�����|]U+<��`,͡x�I���گ�� ����˾VS�i���"���!Q�����B����K�Y.�}M~5V%�(Sc+�*�����l���7�����H_-@�;�p�A:�� f'���y��U{����yHˋ�1e��C�x]���A�� ��um�kuG;]г��I¿���;���eG~sq���yؽ��;��0o�.�w�5�I��Դ�15̈&He��`Yz�I��M~5��r��ފ^�,i������Ju�h_�BE W�����ԟ/yl�%�X�*���墡9ׇ��՗�Q5�����������yM>���Y�(D^� �fj�|L�R�xx����ߖ�f���_��k�kֶ����Hi���#Yf"�f�S&,r�#o:a3���b 6$�p�[J#U�F�nZ'��������[$�a�3��ڰU�p<�f
�PK��GGψv��C��aarZ�� 3�����d8�r�4�n 4��|�?h-�tl?��GV�"u�j�5k���d��R[[q:�� z�6F����D�)`�Akxx�p-n�}��G]+�r$�MSl:B��5����;�|�I~��c=�c������n��b�xY�3�����Ԋd�r�:�VC�&V�i�R0֠L+r�45U�x�_��b>��O6ϰ��v:��X��Y5`=/���[(La~�|y���Y]]rmv���{�9͡V������g�ү��ӵ�+��ܪ�MӘ��C^3&R��<�d�5]� <j.-Uޏ�z��Zyk�[U�6�]%�@R!������k�D���l)@�2��-�kq�6�o��7��U�?099�2�|�{;Z(�� �_8���������+4@L�D����,I�4�����&�OMM�|��gO8�ܱc�K�W��[�����ƣB
��ݲE�zs7??�����H��:�<x�K�!���f�ЛAU�6���vά@!�;���qV9
�%�"�Q�Um ��4a1�z��e�_��m۶:#� s��Ooa(�l)��;���8o��������w�	��y���mN�r��r�Ӛ^k�֭�oV���"�Y5	��Ѫ.�H�� ��A�m��,�_5EM#QP�J�������RD}۶���	�X3��NV\�֍Ώ��|��I�h���A�.�GV�@[S��r�%�޳���ThWwѲ��Z����4���7�&':�=E��A�X H�@�Cw%�v� ��$g����Q�q�V̧�f����j�6���i�~��Q�q�Ih������Ds$j5�Y|!K��vF�q�(��V�u��5H�H�Il�O��`C-�a���i�?A;lo:��:.�C���ȟ�w�����]����0+�]5����]N�|̥�PU�� ��`���VY�l�s�E�oa�##0ɝ�I����X�:�a���5��)!�����M9-*,`�A^>|��/�I�zϠj��F��Й��J���M6"`�q��н6"O*f�;3*�TN5�S#Ϋy��ӧ���I�M��ޮ�4�W�q���+Ռi#��R�fy��I"�aL�,�_Å�T�iS��uZYQS��(���lC��ff���t�P���D,TK6�;�Fq���{�4�%�}��m>�����j��>���r����������W���k�ui$V|��J1�#Ϝf�i��̟jz ,��+J��1�@U�г�<�״죭i��6	�q�أ�=�Z�8M	FF��9CXՂ͙�@S�j}��4?�/�7f`)D�Gj�U�T�}�n�ǆ��y�� Yz�64@����d��S����J��^[K�t4LPVЛZ�*����Z7�o�k(��Z�G���0�!5�h�|~��ia�ǝ6�y����?�x�Ej���������̩����(��+2㹇~T>�v>%����ּ�r�.F����/z��`�����P��tV�N˦i����+���	d�5�Ny��%�Q-�*I�r�:��x#�Z�8̦V�7!�����<�V�@�]t |�M7�����G�������3�?�)�š��.e��	��� ��f�%/����y'Śv�i����Zs��L5��,]�G������M��4��G�6��%�=#M*]�f_��(�5+�ŋ�e`nnF��͋t�q溴Ϲm�֗_���Z�����A`�i���8O?���P붪���s!�>�WM�ZلD ��S�r�XFS��z
�=NC�,��������A*4��{c8V5�zs��-=�Ͼ�o<������b��ꊔ_��E8�Y~G��2�h�����/��g�]��A�����-�����C)�j1H���Ǳ੽�iM�_�>�=6f�����4Bc,�TE�GeT�%�{H�4��	g��]�ʡ�g����a_�z������=f<;v얿{���$����sk��]
U�Bƌ=�6���g��+ӂ����X��G��g�ڟjN4�0&3M����M-娭�����<H TZ�Y�З��{���?5c��+{`����<�d��JW��{�C��yll�	��p����dkfX�N��J�gI��Gp,O��AJ��aY�_�rě Ze�ci3k:�U������(*��f�5ZɓSo�d�M����2"�Gπ`^����oQ~p����yg�ݺu��.1�9V�b%�Jl����+�ovv*w���"�\v�W�mZ�����=T!����<�\Q�E�3�SS�~慵������Ԍ�B�����>�e��*C�����5��h�ӊ���{L.�C�������ڪO�4H�I |p�ψ ����%�ߙu�h�t/�PZX-�ڧ)�������ИyZ�g�� ɴ�F���[��U9?J1f�[�M�I�5I�mR���VY\�zk9�L����2Lm��LT���	�ץj�<I!پ}O��� 5x}�
wUl�)�	D�vO�Ƥ����6��p	��Gֶ��
��q�����X���P�Ѩ�z�"���#:`4���,��fb��P/@B�-{�f�t�1kڢ�a�J[V-��;@��H��`4�q^��I3�ِ[�����+j8U{J�Ba��2�GX&%����}���C.��h�i1�M��,���O�3�ϒ���tl���6N�g���9���Յ�z��,̴���_"�d߾�҃�3��G%
$�P5���9=���	@$7o�1}�?s����Q����F��u��]<ޤ֧������쩥� w���g}�*���^�q� P[��=�%}�e3�f��bwAs ��+��.������O;<L��^��r��HoGgz��Ux�����I�ˏ?��;��-�^뙼J}]}2��]�v��8�<��fT�0��}��I.<��X �3H�0|%Y���� dx��
�ʝ"�ʸz���u ,�X��q�IS5AMO��k�F���ٛ�PL�.��Om|�q Y|�p��hN��쫌݂E 4s3�1����^
�+�6�[0%�9��y��nRhK����L��{���t� M-��ףYqJ��X��ݤ+b��i�f�}�J1�������&��A9�s_W��؛� ������H�8J0�� WISTpQ��F3����	��X�Yh�chVM�Ok�����CM�T��ȩ����i d��O��Y,I]K��ע6��'A"a�ڀ.`�5q�F d���IB��$��i}P��jv "��)�˔� D}��^;����L�O�؏���6 -J������j�]�����nd�b����Ϲ����4j�a!@�3��_Z4�?��OմX6�� 3�8�_)��ʉ�u�f�C+k�! �Ze�@�����@N�%�4�F�֌9[{���h�$h��z�ȭE�s=�)�?�.p�HL-]�	�d�Am��9����͙Ex�Z�k�Qe�����ko����K��\����0��lM�;�gW�<ȩ�C�OK�Y�I�i�O�i�|[����7��[MW m��Z�Ws6ϝ;�m����ݻw����=˄ZH*OZ��yWU�̳-RL��-͉��U����Z�C����u���J��Y�0W�M%�j1z'��
��@3J{XNLБ�V5�F�#L=���X�,a��[Y�ć������Xw �<a���J��k�2�����e37oj�vC��M��a&P%׌���:���S?����Ư�E|j�5��U�����y����"�[[�i/.��-(TJ�� -��g(@Q�=�Lmr��Y��Jk�R@h���VJ��q���M�5�<���IG���P����T��q� ˬ	��$�׿"���.�VF�v��`�f$���t��q� ,�gh$��W�>�f��3R;X�d�ՙX;`��_��|�� a.ǎ}��촠���xp�&:sYL>�Y���e�B�E� -Z�+ �T��Z)"ʼ-�U�Ӵ�4���s��T�i�j �}����\1��E�*�|$ E|�T:p��,� ��k�)��IQ͇�4��H��?�mn��Y"^�J
Ha�kd����;��Ò��k�1�!���c�īQ~
n�Jظ�&�XL~���L_f��M��s��Y̌X}�,���/�n���u
�Hb�M.��8��L,�5 C�@�4����5i����ZUd�q��Q�� ����,�� R���i�(y��'4ËG�5�!9���U_�}U%�bH�F����هz�>�������9��ܱ�N3-R�)9�[��B1���t�~:u������@����R����U�O�>���߁�"�4׍���K6��"�˕�B��D��b�4�����;���-{����`|	4r���� iĪdv,&�ڀ^�Nfb`�[�U}�K�U��B}����V� �qT���#���I=Gym�U�Y���K鄟ko�+h����;���%�/�h��i�QF��aRD*���Aў��_����JG�0r��,@Ki�ip,��������H�@t/'X@���}�&]`����t��<��Z�D}UUS
Ms5��-ՖHV��-�Y$Pz��v�&��
o��?�4B����*� �VX ���0�|�q��$Ym��I~��ô*��v���s�'�"h,"@�AOIֽW~����'�����B:�(V����9J��b�1fR#H� �oQvz�N�עG�$�δ�t~M���kǍ��(��s|9?Kdm��$���ކ��Y�_j� �^`�z�rZ �þ��62�V��
��
�*���i��ڒ�4MF.�=$@gZ����>_����8W� ����̧����"���cgΜ�]1YR�C��1���e*�X����9&ϡ�&�����h�A,cE������	�K��Rktt�1$m%"8WA���Owh�m�ax3����{ �������4�f���Z}Z@:|���A��.�H}b������)զ��1�%(��)��ٛ˲O����_n�����r��>{���?߶m��33�?36vY$�iי�RXD��)��#9�:�c5fU?���|~����I뤋L8���Q|s6$�����^���r/;��V��r�VI��9�c5-�o_�ڐ�M�L�VX� ��k��Sq�~��� %熇��4:�OI1m��Cs�_.���>�̢Y��7i�?�D�J����+�/�����|ͣ@��V$�I6-������|��)$�N��~o�	7m�aIMQ�XC)[[�;3%�.]" A�A����O��m2&��L�V#A;�|9��4�|-u�/���R�J��b�Y����YCd�n���Ȁ ��5 
��/f�y�f �����Qٚ�iĦ&���M���MV&p5�a��� ��Y�!�� ��n����$}}��3g.<v���K�\#S?"@�O��/eøچB��I�<�y�����;��)�˻,?�^��.���g],<��w֖jxx�hC�do��UE��(N������a4E5�MS]{?,-��E���U}{i���i��刂��]$Ǉ�l]���I2��7p�kij��;��U�I�e����a�	��0M�_3�ۛ�}j�~4d��K���t<�Dm����H���~�]�_hk�J��G�)�A����f���Rvvb��\�����%L�n���Jz�:&a���#Ta>��&&�] �1-^{z���#��d�x$;�7���4+N���ڪy'}���{�o�|un߀/����3��D�fX�T��ɓ�]�
^����e͐��5l�7��huߓ�5��j�J�aA!�*�T���͍*A�P�\�Zd�u��]���A���(�8;;�i��V*R:/	����xי%Z @"g�sN� �bP�2%K�li,ٲ�'y�=��yG�k�w����z�c�9��Z�V�D��c  X�IDAT�V�(���ĜI ��sN��{����ntuWuW7���5�n8Uu��3�-*~���1�&3��k�!�i'#g������*K6��#V����j�nR�ԈE��0���{E
UHU-Z��ɂ���IĈ<�ѐ�Y�g��ݵ����s�%'�i.����PO,\p^��5U�I���d�2���j��$ӺE�D�&jj��_�v./�wb�Cm(�&�2���� ���c���F �a�p8�G�t	N��̺��L�]\����)��-�ױ:���2M�y��K����R�:K���t(�q�-��(s�JOY\|��P�ܢ�̌�p���W��i�qC��-/�aG�p,$��)����(2�����癊��#	vv�dm��Ue�T|�s*\CT��4؜L�6W�b����X�x���,�60Ȩg�iǝ�N�.e���Jj}U�����L�0����R�$$,�P�9�8�$,�Ūf��_ڣ]��^��ա�(�����Y�/P���_H����Z�<��ɤ(j�&>��M´�����%w���Y�$7Bx���'�
����ӽ��d�?܆\E/
�B����xz�P��^�6!bqU�F�CGP��R��/]:#�SR�	���ɦdѴFu3X�RR�i�!)���t���p�Q��LR�su����U;yr.�
�2_�LX�� �@8�����ӽ��5zݵ���F��yC��7��;�s��yP�"�S����с�(*�)� �\���Nr���ʪ/�3%������<���uπ�Znڔ*:�DUl!�+:�E]w���ޥ ���Za{,-�B��$�#411IH�2ݔT��a-�����T�z�� ) A<H���3B��-.'g�HĀ����7r��Җ�!,�n�Kk���5�$龳�*R��wd8�@*D�ci;�]�K�fB�Le��Mrۙ�A����.<�A� \�7�����#�i*�'py�/�k y�t�nP��Őz�/�t��On���u$JH��p�ӳhQ��O���\L���'8���{-����&�MLkk#�ߗ;l����%E��"kKl,�<H�>��qIҵ���!*�!�@����b���	��9x�t2EY)e.n^��A�8�� n��e���û�Ɣ�<F.�2AZ�?;l�zM��N�m�n��3ۥ{��z1��⨫C�T�#)A2-ƙ%�$��Ti�-viF9���KQ�Y���^"�l����%��`F�xr��tJ���/m��/ëJ��S彂M��� ��$(�:��a�C�3�*�m�4�w������Y��� ��8�)IRa���4,B���㫍 �i%C縆y��A`P��œFzT��U�9)��1y����U�!�(Hee� ����B�T	���a���Γ��rc�t���S�,Ɛ.�^�*Ҟ�΄�W5���լjs��˿y��U�աJ
Ta( 7��_!$�6zOP�F��������;�
Hˤ��޸������(�2LO���HʁvU����z"v���8�C񾌴11AZvG��zQn[�#J���B�I�v���2�|yU���!���[II�e�W�m;�T�( a��%K�7ǯ��1��`Â�����*��E255Y�a�� K{B ��b�/rvTr&`�l�2%�b�jJ�Q�Q!샐��Y���j� �"�n�i)T����y��	g���T�^��c�� ���kv��h�-�7�;И -z��܄y�o�����Av���x���;��z�^u�����T[%jH�Ιb�0��+O-8c�33'��T�@�隚��MOOs���up,a�F�g����_�vM�B�C�(�-�+BF�g�F�)����q�1��J��Q�Si�)&q��ȿi��
��;f\��d�[j�	�:�=�y��B�T}�����Ď�b�P�Jwr���+�3ƥ*�8^T][,·7,B ]*oX��]��o�]+ӵaQ�%Uk���@[[[�9rD,�EMNll`��}�����񻋇t�v��*&Ry��o��N&�P H�'=����K���12��S��9�E�ȓϿs���;T
���*�0c����?99G���i���R��l��Az�����M��\&H?�ssٰaf�Q�O�,���0�����E�p�JV���u�]V�@|%�}�*�$��^�*�����{�wV�B���:(+�H���񘔔 ���!��G��$8�uD���Z�E��t*�Ef�g�R�/?P���(P�N��%��6�Τ&�N!��r�ϲ�,>�8ܦ��O��彑ie��i� %�	�Dn|�-ӿgFI��I�<�;,E�	�"x�(A��uw�E���"MUG�,�#_r,V��/�J`�ړ��#Yr��;�?�����S���GaD]d���}4F�ZB������VJJP-�,��3H;I,ƞ��?UVʐ*z)�)i�W�&%;Hi�A����|E������Z%�))R������1��O�O����If0*މQn#q�=��d�(��qq F��XO�|��o%��{�}�"}K�4*�"�'�i��b)w��� �Z�&�[jQbw/3��9J\I�:�Ʈ����zZ�kE11q$a���?��p&���3i��$�2�.6+�ٹb�F�%�O[���N�U�_Ex�uI�p��W_���ر�ս��W�H�LO�뱔>ǌ��7�Ր�e�S�&)�%�4K��:)�ɍ�^��!		�d��UY:��M⢪瘿˞[P�I�%qׁ��h��E}�A�<+l��Z����!G�����2�@�PA�� jX��.���겪*�_s$�Fe|�E�죰���y2�����GH@�ԔR�Fi���?<1ᙉ�=�
V��.�Ͷ�'[Qv;��,�9��}�`�pug�3�����#m�z5H�(+'3� u�W�@��8�D�چ�=z�85;���;{�zk{o����#�iCĴE��>dr�T���$MIjr�����MK�SJ�X�e�[YMBƖI�l__�pV ��I�(ݕ(d�C5A�
��C�	��X�����,��Ȱ�(7/z����˙�������s��g˚v�[J��U���ԣ��&��q;�8�)����OY�MtG"�����߸�:�z��؂hұn~���w�V���KW��Ls���9����e!�D:X���٢��n��bO���SI������Np�A���w'��
gp^���,�s��7 z)(��*��.�x�!"`��oH�R�=Ʊ	��;PY�1D'Dkmk}��Ro8�Н�t�����ف�6�!�I͈^�\��s�O�HO=Sʎ�mT��w��X�p��lQ"~tA�aIV!,A��3)I�$������z�f�"�2uu�t
����HҬ���R԰�c�KV.fp��u-UH��C(�T����{_��K�F��\+q(�H��R�r���RU*c�ƀ<����y;e$��`S"ۏ��5�������Y��j�Y��	B�Dl�d�!<�%y@d�V^�� x\\��U�J}Ԯc�m�����8׈���3�*�@܀Am2AZ �TAv�*2��ɐib8IN�t�xR�r|�jX�2�)K�HI%�v���D'5�w�CJ�N/�k��g��MHS�C�@�����滑��8�߃G�jMJx��(z���~���{�(	Q�B�*m��Rn*@�ҡI��h�*Rׇ#4Oω��k��
<T����8q��}�'��H1Z�w|\mۺ�k������ר愞o�����"�i�T��j5^�`�	Fp��&Ԝ���\�")T���������s��d���`��*�"��@8z�LId8�l��+T-��A�$�:;�(�G�+Dx���$9K��$wdq���[��<#����{���N)�������C�?�&�Jm����A��Q�e��U�gy��M}t�\�k
�P����Z���Q��E7�j ���ڱ�F�$u�ͨE�7��T�+�Rġ$C�3�1E��tǐm��4e�\!}B})CVT̞t0R1|z��t.i�qzҶ��XuIQ�.�^�2�B��cz�[�]յ���U?��(b�R�sh�PU�.�;ہ���H#U��{�@~� }���G�9�ҝt �R�r�q�`�'g%��$����/��o��R�o|�q� �c5���y�jbQ��;R����t���b��5��+����@�Q1�20^�yUvgB�A��"I��y�dU�3I�R��ٵ=I������y��պ�\}s 7�%5��ܩ��Ԧ��'ƨ�J��.�)�����@����"F%�gGԽ>�K�����;���3���}����6&WF7��=�E8�'ݎ���2jn�EMr3N(�~��U���FD(BU6J�:�3얺]R�,���J����4��T+U���X��3�K���Ĺj��9��=9�z�]��sԌ"-]��HV'V5WOZg)S�M�X%�j�ch ��A^oll�bvo�E`���wP:�Q���{.�cQg��#�5����&	�"]M�L���UUh��aꠐ"q��`�J�_'BW	�9m�'�Z�����j����nBV�\B����\ހ4O�L#��!�G�P� -����-���/A�na��� *�$��8K�����x�Zq���jeW���j:ӑK ����ڗ''?l�`o��<?hjj*��qq,��w4!!�art8.�Q|0� #`H�������TWW�o�Z�}A�	���K*����ص}};�U�j+��)���*��yF�&K��?��i�/_>M�2ߴiX��[&� �����&*��B~����FM�F�ތ@x�� ZK(�i
�?K�RYY�<�|&� �M6����D���j/ԃ�}q6	��¬iݳ3���e"��b$B�6lؠ�y�T4���f�4`'�t��\����inn�.�&�6yTf"�H��0��<#0"����	���F�>}�v�7�D�P��#r�!>)� �p�����)v���ɉ3��#���V)�u�4i~=ř�k�LF tp��$#�q���ڊ+�u�։T}*A�[�3�#c	2���T&�����������tGG��2M�VC���ej�P�ǐ[�E��iC!�T!)nڴI�Q�F�uJ� K��T� �
�쬢����~�Ot��մK�YOO�JJ�M�s�x�]r~��1<,�ȴ}�	��*٠�x������]�V�={�H(�v�)��lP���0�֝�i�~�D�Ƚt��RK'5�STt��q�⦩D�~5�1����M��rCc���Q?>S�;w�6o�<A�*_��w&H�(���뒜yj��?Ç��Ť~�9��Sy���T��Ռ!r�x��T}�n��{�̙3�����B	���tiq8�X���ac���a{%��*�h�'&&����XI墾��/T��di!(�1ڲ��������C�H��C[[+9�T��Ϩk�����s�=��*Tu�"���$�;ccpYz��pZ��fz��%''O���z�������LOHHN����n	�[p8��ϣ�ײ_r�F�Q���E�SSS���<�B���S�j			��F�"�s�l��9��1A�0��S�����C���������]���MT#1�l1�]��-�P��3��HE@�;��Dإ���	�;6�*k4r�<y�v뭷 �_����S�VA��Ƣ��'�K3L���B�t�J������xt*����$�Ѹ���I;�
���ώ|���`M����3d|��HR��P���UWWP}�q��hKKirRE��y�f�L7 Bg�8�X�b�7�>�B�.`��J{�*��4���tt�� ���󆖖�'()�
������'&$�9�y�zq]O�v읙�;�WC�N��8�s�L�Raq�UR��hIIi�.��edd���I�٤FM����AN8��˪Hv�p���n�L�#�� �DR�Oz�ӣ{z:g�׷����oJrr�r�����;`8@5��=��ub�>�����AM���I?��s.%�
��ԣ����o~��1�����#&��H�&����L6HV� ��S� �F4D۫��Ŋp������Linn�A/�2R�.��M�H���*���X��$�s%q�4��QxX#��m���8����J�Bl�bc��Ӵ���{�����HJL�zh-I����x�u)SJ�d� N�]G�n�3&H���n�b@���	ry~������N��hn�������#vג,���Ҧ��ZXc7�b
������Rg /l�`�T�pb�����Zll<�Jc) "}2�S��45u� Cd��!s��	2�����T��hxg܇N��i��%I�gV��Y�k!�v͈�J�����*i��ܑ���z�}�8/=}<-4ѴHu�eA��@)сpnPE�񍜳z�*f�P}����τ��i:z�fM�JPU�'}ډ[��g��=Y[�h9Ҥ�t�H$9N|�*�8ю"Cg�З�f�qL����e���po���Z+D�,6pR �aם�5�2�,X��HQ�K!i�4����(> N�$l�==�`�aH캱 Bm���<��(�j+Z��,=��&U���-IP��������A�	*7j�Dr1�<Ɖ����8"�,�zq���LID{�ҝ�:�S����9�*V�N�Н��$&Hk���(�r�ٳ�ݤ`�qb���7�!%F�E����J.��D��b��o�gkk�v��%q$K��RU3�h�'2��l";��꧝�\#��I~�����~�"0&1I2ҝ�\U⑑c(Q}�f�L� ���)�
M$�/I�@##����ĉS�ĆM�\��.Iϸj�:0��aY,AZ�o1A���h8���$%q��B�zTZ�LI�p���ѣ&lE K��Th]]�L[Z���2r���+�.I�ħ��6a�T�B����P��	���`I���Rg����r& �W]�9ՙ�{�^*�J�Wآ��?�*Q@*�]��L��  �U&7we��Iv�zR��@{��$�~�X5���$"������!T�GKK���8@��q*�|DՋA�T�Ey_�����b	���d�yL��92��0��8��!U������,uH��Ͷ��ZXxJ�l�@WW��4�D�G΀�mww��_xe��rH�m�1Au�C�pG�v|#	��n���#��Z٫efN���I���)�t��Z���L������'j�s���nM�m�D7�BF���������yN�B?R�<�'��g,i �.^,D��X���'M�>��r*�XAV��-_~;�<3H��(B&bcc�=�P�	H�J�Ǹv��T8��$A��棏�k�����Q���oݛr����SC�Z���ƦS��$�;�b|�)��8"�("g7"�#")T#���4"��0%�Z��.���k�ج��T�d/V�W&H���ni�0�E��IV�yo �%�N1��ۂ��"��w߾OH�<��}�=b���Q���_���Ң���މ�3H�7�:��\O�ˋ�e�~�'��{��y�d|#@O��*h���Y-X0��h�w)����
���9l�T�-�*͈M%�s&�J3��hmP��f$���mi"�q�����6#}T	����I��Is��	c3����A��~���o+���G�o��Ñ�~�r��gR��0v̘1/����м�w��*��h�K��x>/o�-��d0m�����[m�YL���9�-~�J�R�*���޿?J���n�� MR�bQ�fvD�X�������	I,Y�f���D�{��YwQ��o������ê9��N(�|��[�C{���j�h�+��ٳ�iQLUb���'Sz5�)t�M��UW5��IH�f�q��Y<4D�.I���w��j�-��{�c/u��i���JPGA[L���&�2E�����;x��A��ݖ�"##'z���~�₏0���%P�7&F�aU%ND��#��?	2�%T�exa|"d߼�]Pd`���U)�:/ �DL��G;�D��yG�^��2 ���@�Ր�=����ch(���̜�6H3虸V����8@E8��awm9A��*��E�E����^��U{��Fx����A;_p_�܄ˎ5�w)��3A��Q�/��!�!]�"�z
$}3�Yݱ�a9U��kT����N&H���k䷄	ҏ���K� �@qD��W�"�I���r��6�H�P��f�fޣ�>r�q$����,�<��n8r��0A���	����x��x����51��(�I��<}�jAD�c�'sG�]ق �-��r���[��;�0����$Ȱrhs8+����B;�lVܝ�i��� e�N��A�(|�XpFj�B�as/�B �l�*��@́ڔu�����A�f�ޫ8$2�T���A�������MAdX��*i� I2sԻ`�3䭕¢.|�I�*}z�_�}���}� �:{� �
���M�s���+z�� 	RFۇ�!r��d���J��vJ�f��oX@�}���b���Q~F�?����2�0z��M�ǘ��X�摒����l�~t����+�rd"��<>ԏ��%kH��eL��a�=[F,�����M+�ș3ߔ���>�-� ��$#J�Mu9;��qO´��{`���az�}vXy��0/>�f�Z�v�3L�$)�Y�|$--#j��?C�AT����A"�r�:t��#G���p�c��92|"p;0�}�9犯s���C����U�Z�p�]_�ӴisV�9�[/%H%���^y�ϩ�ՔM�6�v�ܹ�~>|�zU�e$#��H��>΍
͆A�"���I��B����'�;o����`s8��jk+D���:��Z9}�t�YgN�4i�/��<�������0�����nX�.�!�[ R�z�(���P���w��f.^������Z�y���˝w�	rԦN�*��mmm�7�t�z�����}����%�6H&G�8&H���n��շ���y`��b��`J��;wQj~��-T|>�
I4���-[�m߾�$�Zl0�'�x��K�,I��B��0��L�6<@L�6��]FF���eZ�
����b5#AΘ1g�]w=�^FF����Z�xll��f�]�믿�uvv�M�)55uI�����}1� d8޵ ����=HCV:E��$A�����ի���t�"����;���W�?�:R���v��)�<���٩�^����z�;�7r{FDu�?K�r&j�0A���}<a呢T�Ϊa�<-Z1'/o�3��៮�p"[�v��y����%}�����{���Ѷ?r< F D`��c���I ������R&��`���M����q�.Ҩ���tא�33s�U���^~�5��Bz�*����I~��'�����:��Ml4�6�� ���6���+hX�U��ԐA����;�3%������əDޫK���A"���e�n����W����#�$t��	І>���F �bc=x�B�hxAY�����V��#�B}��сo���`���1��x֬���}��~їR�b�k׮}aڴi9V�����p�?���H�/�Ñ~3Ba~����P?d��P�?�Š�F��9���G�J3Fx��6��͍����ZZ���W�w����g�m�?����]��͔������))i�@�2��5�6ډ��^�o��G-/o�F)�G+BB&��}��������ϱ&I`g���P�r߾��={���$)%0=~DG�H�+AfeM�����*2R�c�X
Oמ?��^�����h���3G���uݭ�>0%-m����[����q�}}>k��>^�����k3f,�>�d���C0H�$ȵ+V������B����B�Bzp��'���*V��AH����{##���԰<�Y�
B���t�!�����c<���7������$f�ޢ���ږ->��/-ٻ��Wݑ��!m�����^����~���55�FEy������oѪ�۵�?�XCvU�;���a'Z�A��P��1AEj�����i�����F��k��P�̙3��^�������s4))uHȊR����g�7��C{uuɷjj�J�A���������x��O(G����k��X�d�v��q�eG�#!a�4�x����m;���F����#���� ,����O���b���֎=�����ڥK��G}T��w�����tVVְ���su�5�1P��j;w�'�|=�'N�r�����?�⇇��D�T�6i����0a��jݼ�-Ԉ�H���1���_2�_��� Gʝ49�իo�eÆ�^��8 �S�N$�~���I��-Z��������|�y�OFFV�ĉy7Z�!�$V\|Y;vl%��ed�߳g�'�V`I��w����̪��>m����Y�]�xEkh���m�佞>�V���`�&�p���Ѣ�n����`{�d�X�ɡ��T��rӇJ�u�ҥK����C�{�mCJJ�r"�	fa@,��5$=n%	l����ܔ�=u��f��3g�6n���7�:��l�����tT�P!�NHHXD�'�탯���Z
��Ƙ �c5"Ϝ2ez�5w�A���@�
8Y�6B������J�'U.�:xg>����&g��233]T������9��LT�k�{D��$�f�wRɻ���3��}�ʅ�S��6I3��-T����*Vl*��r\NN�d3��#�i9��d�4�ӈ=+?���Ξ�(�T��(ihٲu�5��X�UL#~�4j�ƍ�GSS�����#^WW��Y�<kvS �*Iw$A�k��9$��i�����y�����BF�9'��/H�Ӧ�!g��B��$o�ےt�ԟ6��[��������3A�~�����w,��q�F`M���`{���_۶�ᴣ�7��nݺ����|=�d}�HUy�������V����X�}���/�����@��8��Y33���8��US�����i�H�� Ab�����?��#�2(A�=���M�M������kg-^��'�A%��?d�![�VPpI+//s��E�G��$��H�$��I����h]�ͽ�����'�j� f꣭���@���?�q���t�9��F�#(�O�.$n�Y��~��۰޿���hh�q�UU��G}�}����� c���p�C��8�[zIc���Bgn==�ڤIS��3�i���W�8Nl���M�6��v�wќ������#h�+�4n1���D���X� ��v������>�r����Gs�=*5kvvj�رQL��@� g8R�S��fmϞ�h6�����>6���}��H9�	r��I���s?����Sׇ����T1J�F��T�pDQ ��Ԭ��s�S������a�xc6KM�v��I-?��+..�H29v��u���GGJK�Θ��DƟ�S�i��"H*�E���|x��T/@��OUU%���T{��Zn�"�^�(y[�ryV=4�i�S�i�vvy��_ʛ<y�7M���E$팣]> %s���у=���v�ث�;wnH��5k� $dN|<R��?��+)�8�#H�!¼\����`�Ç?���H>�JaM�ZZZ�ؕ���Ο��^��U! �J��('�����ퟑ*>S��׾KaIk�f��c@�VwȆ����a�ܥ9�ӳ���6�\+�VA�Ҭ���~<u�ԡ����.�y�������/^�8�#g�8�M��bL���D[�r#�~lўx"Q�^`B��{ � ��w9���_He�#G:;;�,Zt]ZLLt�C���lP�[�������V�v��4�2�QZ��xH�w�Mk�X\|�׮]�zܣ�=�.466�bSS9r-"m��̕&l��́@U�/�0A���0A� ��]fgO�/��x*F"Ğv<K��W�^t��R�QJ���ϧO������M��"��M��jN�ҩ!?�������@�	�	�\�d)��kEE�h���X�Z[[�����g.\����53���r��N�0r����l�%)2���X��q4�v����lai,�mmuIu���?@��k"Ȼ��������/���Z����ƈ�`WW��f���9a��t���P��IIɳ�t́���M#�#�,��=�����.]:WE�y�����|aŊ��J��'ZE�X�֭�S���7�b��z�jA�8 Mn�t����l��7s��Ldfl�c�=�ω�Id%���,L�n.���9TF��6%�&M��nX��ӑ�(M�z���U�|WWw'9�]��x�\'�]��juuM�s����Y�*��!%�a7i�Q���a�M���mLL\&����W�ǐ��8y����޽���~�ϼv�غ��w^����d�U�+0G��r�r��N�L���l99E�g���#6�I�,D�6��I}�������꠿�Y�'k4��ӄ�U%M�Ij�j��n
����r�+�����d.\/Z � ���.��~au5I9k�0��ӧ��I/v'��&^-,<���ܹ対�b���'_��f,:�dk�A���x
��11��K���L9Q;��bA��lY��͎����Q�A�~�$	�������T���条���� :��/Ε$�~@�K� q�t0w�'x�y0^���F�}�ҪeMl���x���	UU�/���'>�h���>$�M
)w�̅$�R֘���!%%�$��m� CJ�>�Ԭ��=v�ܩכ��L���)3H=^K���(���W"fta ���O/<�4J����̦<O�BԦ^�П�P!0aBn����񎗲����7�ۙ@Z�VZZL�0���~��3��-o���|�cEo�a'�Q�HZ�Pv6R��3E� I�C��:�IIYv��uITڰ��Ȅ��z�i���d�J^bfq>3f��**j�?��C���!{mM'��?���X�X�9�>�y�^�i�0��Ԗ�ѱ�f� ا>��m"�j
2�#�c.!0�_�����ę����T[�`�4o�SLvHU�IfޙJ��f����$M����ٹ�.\�p�T�� ��o_���Ǐ7��`؉Ϛ�p,9��!Hd�9x�3�g,I���CIGG'��1Քu(8���ސ��	RmڼL�I҆��i�vtIdp��~��_�xF+,<&�#17�;��f@I��O�����=fI�$:�����J��(�%G�$�$�8@K��A�\���%���CH`P�����So�����ޢ�+��c"9���z�X[Z�Hݜ���G�!l����5>��<��4�EM���ю'�	��m�s���ϚSYF���C�v�Jn��CN?d�;���t�q���'1n3�0��i�(.���b����--�~�y���Sx�䍇 He;�В��͛?1 ��&ɹ&�6'~{%+�@{{��#LTB��H��=��5�pZ z^��!�yj� ��=����->))e��M(	��[)��J�˛"*�466�R 'C�
�����ˎ|�x@�S�̤l&-��U������+~$T�k��=��h%%�UeF!k�#�<񗬬	Q�&'��4���=m*f�cur��>��5��L(���Û��h����\C�ՙ3�O��)�fTq��
��#�G��td���:��;�`"h��B£<�$b�.\�]�v�c���!�Rf�XH^�;Ţ��]H�s����կ~奩S��xk˗���fD�\y�U�_�U����גm��T�Y��׮U�&;j�?m�5H��H�R��Q���U�,&H��f��A玘�x��$}1��l+�����z.^��^��BI�+kj*6��f��#�z��Z��	�)==���HR�v��ƅ͎b��O���.1p�����}���s"I����׮����yfmS�$@�
�W��޽�D�9l�@�s�7(�Y��E���N 	��H#�[����\��R4%=bBPS���&11�� ��K�.\-))
�B�k�{�6S�D2w�u�yh��T�P���u����f�����^};�;����,�2 �W[�j�7|���P�X�����w��ᆵ?0��BKSS�#�R������x�=�a6 H�FM0A�t�M��6����S�;�wt��xA,��G����Z6u���%o�FZp�}�����9�ԉmBR��}�H`�!�q�{�=�h%���z�Զ�\j,�ϥK�>��c��~Μ9q���t������S�k�j6�ӼAj�t��Lpo����bb��;>�N" �F�d��'j�������~u�ل������T�����?����{�Ѿ򕯬�6-8Yc
Ou��t6��fEi�D"�.֡R���/!�˦RI�d$�\���w��環{*)R�<g=��SOm۰a�|_��E�nH�Ͽ��y����s�����X���vT��';sAA]]m��c���>p3y_6[�[{��i��i����=����u��""Y�}�j�ׯ'$J�t������߹Sy�
	pxj���S��QG�D66V�=�Nxq�߾�2Ӥ��k�f�@��B�V��$�����_�����?F����7�|�*W�ڬ��D����~aS��9����[��kT�1:�Qw���56q���Õ	�����i9��� �Ez������XاO�C1��i1+$-|C8n\4J;娬,1Q�BJ��'Ϧ��%� E=zL˷�6�&HE��@,X���F�"IoP�"� �4�.Z4����/~q��?���'�|��]�4i��5CBBn����n�y�������d�q�I��e��2� ����:��2Gk���;H�/o�ٍ[P^�؉�<^#��8�S�^��'..�/�L IIiD���z��S�״w��+M8IOVHw��%��jݻw���j��T�~��Y�;���;&Ǡ]ڋ/���GR����n���ARk.�^nNNj~Z��_���+�={NuQQ�g�ŗ�-[��%Kn|�ʂ�����jQ�P~�(���={>1�t�r#�j_B<���#�����3A ��k2�����N�2���cwK���4ZZZ�f�#���/Z4wٌ3�.^�H�� �X��鈔��#�7==�ȰX;v옶s�N������g�G;q�sQ���}��{�4��ٳi��$B���v��˯�	�f}}�:�V&��nz����r]8׬���1"�ر}Zn�$�?I�'�9�_����,� ��"3;y:8��q$�>�	�jDC�=�3u5775�t�i��1''�Ԭ�y����رQ����!"��z�$u����ո@2�ܛ�$����?��YA*V��:w��,擓�laK��PD��t�6�@$% ��\R� �A������ɠ��D�\k51�/H�EEh�PM�=Rl�ٳ��A$m"�h��6d=HߖVo*V�GG:�5��bx͍G�@�����������Sg�
c������6�R��q��o�۷돍�ְ��AN�6�^3�,�h]�TH�p?y��O��V���';�Ա$UnE�gAXVH�j*�������Y�ƍ�<��i�N���ԩC�i����򋲲�=�>#�:�%H�S#ϐ<�3�A�ʉ�y��I�܃������ݟ���MJB�\�HI��7�ef�ν�{_䤦O��H��FQww�X�T<$l��/����H����?��"3I	�� 	x[�~��hdA5Ҿ�s`;s�0y�^��@��?~��f�)�Z���ΘI"E&H{�2&H{pz�T��L�^`�IddL$��qA�ʛ$�|��g�O�>-P��U�DZif1�����T����~Cm�s||��)7�?\�r�)�$(�<�+�Z��<q�D"��Ҋ���
��՟��P2����a�d'�PY~�吆f�$�5wt���/E�4J[��^m���ڕ+E��S�MNNv����ߑm\ X�d�sf�q�ZI�X�����q)D�1{i)�F��C��e��+�=}��?a#Ž^Σ_��H�#�~����z���@ܯ�ަt�1���9��z

�76���p�L���Muv�WP֔�����r�����ʣL1���L��$���˂[-Zp��8P���y�=iFƘ@
���	(U��Aݸ}�������}������k����/	������`����[Z�^).��K+�綼�8}��"�٣M#�7$$H_��s�C���Һ1pKA@�2�tS���ջn��`+[�|-e\�ת��U��־��'~�bŊ���Һuw�T�&G�)�j*W��6m��w;Iz������2��}If弭j�oh��(�6�Ѹ����h�p�ON: ���=��8l�L�V�>���#`�|:ep� ;[3jC,���~����� �+�	�+,
T:)�g����#�}���~�-Z1}ƌy��}�q�SX�ZZ2���(�F�KHJ,�t_?�h�Ä�(���B�J�V�'����ȱ����=P__O��x^�z�7�	�;P��v�G��� ���e��f%"h|���5�B$���PE�P"ɤ{����>���yyy��"4u��;�|�]�.M4�e����+"���P��ťkii��kkk=�Ł;N��'ߘ~����׮���:��ʕB��<
����_۶�'u�c���4�a�G��7��Xy�F��F���E�	�Z<C�5Z(���
�濣�>=, ��8q.yE�d�WIb��B9������%��l_��>}V4I�NJJ�g�����/,<AI �:B*Pɢ��J�22�?��gw�����ov�a�?+���������7�ĝnjj������ms�#`\�!���;� ��>��L�~���۷���m�fԬj� ���-/o1I�{E���j��旞���2�x��g������#��N�[�궗��f=`EF�	ĆE+6V�v�A�e%%_7z7�n}��|�Ʀ���J��\�}�{��hE��S�y���2)}���⢿���|U���<_�b�V	\��аmQ��\W[@��D��:H!T�I� 5�PB��;�{�5(J�
B�*�� �A��k@ʉ�w.�o8{�W������;���¶R�(v>�SF�3$-�������~�D^�:ϐMj�(�^�+�0=R5�@���7�-*��@(��M��u�s�������6Y�a��#�(Kkny�7byEz���Y5���0[�O��3�����+Mf���ʊ�;��ui[򝬄�-'f�*����1��ſ{ݩ��=n藨,�~���A^@GH�:o�T-`Ol����m``{��͛���M��f�A|���~�I��3u��5�^(��m�p?����\%�ǰ�	|�*���_B�7y��pr�1��̆O&�+�ƹ�q˃i~�\ej{�G^�T�ZF�����?Gm���r��a�0���T��u$6��w��ͧ�|�m��*�IF�S��xW��U��;w������ӛ�)ߝ}�Jx�w�响��B�p+��N�3e&����$��=������\l�,:/L�⭫��܌�G���NP�9<=U�C��q���8-���98>�=��ڿD��
1���bήygݮz�h �e
��}
�Bi�TO���BB\��7\���o�+�o����ق��U�4iV����+$�(zݾQ���5���Y�Hw�R�T<�:�!��Ѣ��?zne�_��,����E�no���~��i/�-E��'�-��x���^Y�BKᮑ�F\��v9�ӠP1��l��8w5�+c��ȹNA���S�X"�go�ÿ�B�n��jQ�^^";���$��I�O����{4��c9����8]�&�sy��,��4=���%������+����ҭ�{�{�O��d~�k}���o"��w>�^g�ޅ̬�����/��k3���t�;5���Y�����T�6�d��g`����{����j����o�3��B4ˍ�v��PF|��iH?�9�"d��O�dkyc��L��l˵���8j�,���t��5S�=q�S���t��6�T�\I��u$��UR��!5=�g5�g��ޢT*&��f�~A�D9L�AGi��'�7�� v��MH#X�[��������P�&�������q�άy��˗�OP���ܼi�wf����o���0I!	��/�׍�YU�ؗ����25��<5����b>����ߡ��������tn���}My�p��gQ��ϛ�a�o�+��+���'���Ǐ��
"܃�n�6��!ɑ��pIY٠Ott1lS�vAuS�{�Y���؍�1�5)3�1�{���+?Gn�܌�w�y��x�в�/�>X��n����������K{[~�+�d����T�[}�������ٮ�{��F#�eie�m��{;�s4�wF���Y���FG׿x�����ne���*�w��k�#.��ٹ�#�G�$�G�R�0]���K�a:ß�Rl_\�)^�E��Zt�5��V�e���ML\љ��w���9�'�Y;[0[�+�>����o�:�����5�cN@��i5�5I�J�t^Yo��h��..���&ss�ʁ��ږ$ge�k�,�л�}i�V
�c�U�e|4�^i@ԇ��+ٍ�E�
UG1~~�����,�k�Xv��JO�����ۄagZƊۏ�͛�ᶑ8rN�6mt+B&��ɣ5l8�����t)k�����s�9\M����+*�j��m}QR���g_g��_�t��\��Ӱn��c�oڰ�>�q�����fɇ	$ɟ��kr Ҧ��a1*����qr�H��cr_61�8�&��a�w[ ��59?�	D�n�_�E�����|�7psu�����iȠ���^�+�j�nu�8�^A��v�6���+�X!����~u�#ߍ������?'Hۖ�s*�����Kc�V��/�� 8��D	�wum��oי�v'38��8�N,Ks��~x�-X�\���w/�y���ӳ0m���П"�Ho�WWSK�w���s�8H�7��NL�$,L��x���?�����V���a������[���<_n$_ڨ���y9�P�������e�T�>õ����D��m�?��M1X�Mv?,�S�ݵ�b�ӊ7o��ޕ�߀}[Z���Y�X�7[\�Fn7��m��KL�ȀO��ބ����>������̦s�r a����w(!Veq�B62}�G`��Z����eh�/���y�����*���.�S�1,̝�)�ЬA,`���],ˋ�ٙ:^:�چ�����馥6�٘~��J3|0�?X��p��[5ebb����ay�&��N�|��e�%�+u_�nig�SC%�����,�p���I3���C�X��f{'��i��Aq�����v�Q��p��WRzH���~�_녌E�6�}SY�`miy&`X��6̈��Ӷ�#�o��3R ;�"��x�(a6�
Y��C~�?uǼgd�)����AU��$��o.���*��77�(M�w?(�0���G]`�Q�pM̖�u�c������mY9qTf���r��)�(yT�&𻧄��Ё���\ȼԬ+j v��(�2�)ط��nc=����[Ü��>?�^8�<&9zΥm�.O�S��Ab�u�
ؘ(W��O<��FT�yr�;p�|h씥��r�B����年B;!^"�͠C��Cg�GZX,縰�΃�d�ihT�H��:��Y��.�1%��&c|vW�77�@�V��`O"�o����<*�i���89�J��Ӛ_��V���荍i3_G�"}7���(�D��ն��+}��hf �L]��ȁ���z&iɜ)��C� ��M+X�yuZʻA�H�������$�q2�m� �x/Y�|xƅ������QF�:��gf���d�L�����6�����]W����ɷKC-�,��=GNBr;ѣg�C�t�vv1�԰V..6M������x����e}��L�|��e6�7�-��2w	�T�N�fo�+K���'�ҭ��ifeu�l���۰�3 �n�);�h?WXH���$�	�@}�B���W�a���k777��!s9K��f��I��d����B��i�Ņ�ª��+�<wR�/.R^�7cH�cރ5�c�TP#ZT!q~D���t�r	�b�,�����	N��T�=����d��������r!���������~�w�����_B�N�s�35����Dw�S�����ǤMq���/V�eϽ�A��{�ͪV۔`]��Һ����(F�����$�����9ܣ ��ќ�}�*w^��':SD�㝬�~VVE�e�'�η�تm�(L<�׼�&jǊ��W��ᲈc���f�+ڇz���7�ف$�Z��<~yn��k��9?z./�+�8{EF�r�ԈOM�6S�:�\�Ǚc��SG>�IOa^�t�PPD�淫jU {TqL���+2~��&�����5�&��$mm���)���Uv���F1аA�#���5<�ߣPH��%\���"�Zs�����L�DW�ҍ�%��C빸�Z/�����O1�B�_R��R@\>��vyh���y���dd��j:ߚ�b��sq�G�����1E��v���2����^�p�>��J����y�AWJ�?�D"	DQ��k�Ϻ���q����� �|�a�:'I?��ӥpǏ����'(X@E��#r@2�/;$����(�io|��׋�3B�%Q����f���O�`p�k��s8��� �M�Q�v~յ{�}��,�/y���D% ^���p����J�<�ٲ�JM(UPKe�;C`��w'b�œ9!E�����Mv�mt� A���]���l]�����~��}�?KʌJ�6��|x�[�M�%h`��3��{4�ڽ��Y�f�� ����U�� ��l#���{��� �A���!����@`"w�^
颗tC"�ԹU:�U����s_A�2�%)@��I>����m	�����6x��_�`�)Go�����+r�s�g5����oG�u����9y�
 U���pXc�x3�!QzO#����u͸��$�"�0�R'y-Djg���`����[��aV4�-��p}>��Z6#�D}�Uŋ�j�1>˴�1�t�dW��T��w���`<©�2K���R�2����$CO�i�i̓ݭ6ϰO�/�?j�͵��ҢJ� &%�����T@v�;k�()..Km�	��|�yeHL�S�[K@�?G�7��~���{����è"BaŸ�~���cOq�e�EEՋ������"Hr��w�,55U�q��#�8G[��&L���Q�������U����9���������T6����oO�IO񍽚�Dq���Egk/^�8�c���Yqݤ�H�PE�NͰ/�qV�5TK������݋@��;�}��{e���2���tr�DZ������0dddVM�8ш*S؇�)及$��q����K	�!�1�2�\??(�,���fn\��_E����Z����j����ϑ�.n .H�X���~QF�%����x��Z���K ���8e/��{��G�c������Ŗ��i�F�  ��k���`��k��f�Ms���g���l�����9w<)S�Y���d$ J��3�j�I��Y����Vo�Q�KX89�i���w87Gp�o�Y������RN���x?{��������g��'���%�R�T�$9J=Ⱀx+��b�(ˎ���W5 �[���j�HY�Gd�/\�)��"�� |ʐ�c��NSJ�촆rA�Y~��u�(�8$3����T
E�ߙ�������N�n��(u�f�rԵ_ň� HSK�h����M9m��
��������z�;��>,y�lN���@�v�f*�WH����Aܔ�����UWW/tv��<C"V'���� ����]�LY���1f�\��1�B{�^��5ΡE6������Ih��O9�#�աjO;@�r�c�T�������YU�w�[W�,PfU�"K
č��{�(�p��s?�~"�H�����z�R M]VE.~��ڍ�P�jK�4y�Ϸ�qY�՜Φ��ݩ'có^�\3����5�̷x.��6��OD'��7��[��O��I9=<���#���p��$%$z
d^��l��!K����.���9$/��Q���GB��;x�>�Q��mX7����T�=���PK   �X�X��E!  d  /   images/73d4fb58-19c4-4d70-ae00-297313ed457a.png}�g4\��2a�Q�3� ��w3�`�.x��k�轌!z�� z�5�D� ��F��Q^��~��Yk��Z{����s��O���:�DDDD��R1���MT�ov&�V��}P��DD��������M�%@�,���) ��ϑ(88����������Co?�"�+������V�i��,
����B��Os�M�ۖ�!/�]�L�=��Y��<-�1��y�5 ��s�&,��a�<�ܸ���)?�<��:��˙��9v��ʻ9l�9)�.������x@Ԝr�	�B	4\555U""�fzt+�ê�NFJ��˫|U&�m�����5{;u�S����K�>��WW�㷁�����X� ���Z�����L���ަ8��K��QS#�^+�Vaϙ %�g}FՉsss�em����3�Q;r�H#8���ޕN}<Y>d��8��ֹ|O�j�3֟��o} ��6��.���˒�d*B͵�aAu�}2s�bܛG_�������6>˘�"~���9�8�9�8�|���q.4ӁJBI3	���[Fk��h��.l'�3S:��1��}��RA�5�QÝ0u����t��I �q#/��ςnl�V�_^αi'�i-�KL��<���g��Y��P.�j��.=;�o�GlD���\�	=�J�-���ݕ�Ao���7;>d�D����@b7r��(-< F�l���!�H���YG��J
=� tX�~sF���g�̯����������jP��w�9�LNƭ���4h�	˟�Z�W3��C�j_ڏe���K/��1��=�L!m ʉ�X�a��K���n�1m��b����-�O9i�УH���_neR���&�B�@��e�<,,�����ӹ�+ܤ�6KC#�i�]��[MM��{��eݟk��D��Pۘ~ˉ�~=ssAqU��)�L�Kݲ��I)�c��5�抎Y���[�E���G�-��3�{\C�������;�/Ru8]�PW�jQ
�{�J��A��C�l�f��U9�c��W�~���e�����o�^:@��MUa��u���M�~Q�Okt�7�������9��V�m�f�t���^��� �.�W���n/d�UPL,^�#嫅�c���W� n��BZ�=�O�KV^�@�q'��L�h����^%�d=� �֜h|����MVWdy���u��A�hh�����A��=S#sU���E�X1�9O���+ӷD���Y� Lk*q�_Ci�=6���8S��vݝ}ap1�l���X*��kj4�cb�����E%���!�l��8m��6rrN�252y�b���Q��}iR7���)��A��Z�&ж�)�G������92����q�����5PG���MsV�t�M��o�W;qߡD�!6H�F��P��x6�Y���lo�\
����U�8�
D���W�aS�mVIQ��,��S$�J�|ἤ^�iB�I�g#Z*�h۱>¨f�0f���}��t���k�9u���E�P���ŀ|�l�9;�V{��:X��m����nW���lSRuƺB�!,�A��c�4�t�,��tۛt�+��6�D{�E:��7��&fu���9%	ܘR�}\擬l@���*G���46d�>x�N�� �K �E� _�4T��U��+Dc6�X T9����#�W�.� ��L����jp@A�z$��(ؑ�8�
�7Nom�������� ���d=��ݠ$>>>Q��Rܠ�'u��U���5�K�W�2�C�#o�� ��$��h���D߬�^��g�z�nA(]@u�s�5dG�⼿�n��v>��� ?9�+���XF`�3��!�oM5j�@f�u��U�l����v%L�G�= �$���,i��S��ıɓ�r?�1�.�p��gW��e)hv|��.� ���մ���%��[5�yԓ�ʇLW	���ԗ+љj�p�e���y�'��8=�ԭ��k�>�K[�qr�42
�xM��m=�'�	��@�]�\�IJ�$'X����uQ�$[��lm�_H�k��tuy;>	A�v8�<a�]��-v��%��Hb[L�M8�C�&�g���(���(3R,��0�u����)�O-0Q���f(l�n$h-�*��Y(!������;�Թ�:�}v[�ž��Ϸ�����.��'az�q(
y��j���!�@���P�I�͵t��u��� ������X����]L%8&���D��Q�;�O2(�=�o�Bד����;3��b�\/�z�����yc�O��~���R��:���[v��G�t���7��hq;�~z���7k�+Dt�t������MK���u�!i&l�ʇ��M�Ö���2=Y$�ꏟ��B �	+��B1����t	c��������
��4��w�T2bb���,+}a������!�d�t/"��.!�T��ji�7�ko0��E�]�����Ŝ��l�5kt݁�V�6Zo�K~���Yp?�-S؈��I��A2���μ����R��ew�F���6:�h��myk>xmX���M��zr�=Ȑ%����g�::;'���P Hu�Q^��3�G�i{�28w,�51dp�:�;F�\ps5�o�l�G�"��J?WK������K���A�W�IX}�$g2�v��[W��(�D�.�~����y��n�u�H�t��˹��m���L�1f��'99q��m�s�{m�{]��<I4A�N�\�ֹ?��NS�L���_~��y��$�`���PGq�!���)˒���8�� ��+{b�8�7��
�c��a��Dv]t��\�n���w��MI�`�I�C�@^i���P*B�Q��^��������C�&��(���BZ&l�N���yw��հ)sK��_�=�ġiY�L�Z�҉y(�����Yg�p����r���/C!���̈����&�!���E�}������dD���#�f���Zl���	�*��w��bx�+,�GO�IG5�8����=����c!8��P��F��uv��H�����|��M���;�xʷ8����!�cM%Ş?���۞(��[nqLU��w{yn�x�u��<p �����0d/)�a�c��G����e���i�D�_�4�Z�V�Kv�
1�#�"��"�Bs�Ĩڒ�-�)�����j���g�հ�>�R�����C�5�7�4Hku���0��9���`H�844�9]����8x�1�Ҟ�T���4��|��_ڞ��*�Yi���X"���R��:W��ǡ�;? ���kJ��鬌K���\F��h�_��^�~�,u�����}O0ʑ����O���?�W��QW=�d�0�z��[�~un\#�.!�D*���׮Y�q�.-q���3�Ѽ�/A���+"�%$�Jo�?:�ת���P�(W�m���1k�8��8��}������j�3�*����]|(��?2@b)���[��|+ִ;6�)I��f����2���N��I8Ů;s��q��[��괞�.tH��p��K]3N�>&K�:3��/�P�A�ʡXSFO�i �0ԣ*W��
�YPf�fo%"����Eqs��>r�D�F��i��!�c�ўГz�)���Ӊ�-[�����nlq�f�1�|xe��}��t�I�#⁎���=񺤊5ϡͳnZ��r�<��u%R��
�'.�:�x�;B�nV�)V+՟��־dȭL�V�=�.f�(���M�E���K&� &�pjS4�3��(�V�� �D��Xv�R<�I��2��:q����BS0/��������7�+���!�b����x��)���"6��"o�u��?�]��{��d��`�Y�>W����Vm������0_�����"i����-�`�֪-��)z�������=Q8�"po�&���79�Π>.����5kvo���g����gԫ�M���l�/z�\�4���ڊS��@~��P�������ׯ_�O˝L�Ps�<�d��e�Q]~'�������X<o*l���"#�܇��T�4��Ç��޹�0ɫ?�لyv��/���6���X�Hm;?;IlU�:�VvJxʙ ��,��zl2��H@��u�|�U�=���?�e�\����0����,�>�pb���>�z��&�$�E��k𗐗�.*��a��c�ɷ(�p �	�ڊ�Y<t�2�S�7���;J�$���*<�n?��C3{�6�A�F'H7d�
ߔ���d;$��������u}�Vߑ}&�Ľ��j�1j�KB���N�	��D`�}WH.�MQW��d}�c9�����Mc��7��_k-�ﳩ[$Ƹz����&w@�Q�|!������
�X�5��dN�G%H���ă�7�Z�0Tp<ڪ�
�Ӵ�_;$�T%��Q�A#�O�BNY����ٽ�co�������� ��:l?��Y.1���#}UM�w�D����~�:G}�(���ξY��GQ�U�110Tp����(�h�xe$��1� ���B=ꆳ;?�gA��7��74���M����&Na4�0`	O�x%�V�w�x��k��Gط��*������Ҁ���PK   �X�X�W��,  �,  /   images/754cf6f1-779b-4e0d-9f61-aeee66719356.png�,}ӉPNG

   IHDR   d   =   [c�k   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ,IDATx��|	|\Wy�����G3i��h_-/��N'!{IJR-[Ѕ�l�<��P
�GJ�I )!����8v�۲,���e4�f�{���;#�d%$��{'����{�=�[��w�se�'�o��JZ�<��{�f��d�뒩,����A�KX���ݯ��s��{�8G�/M�Y��[��A�w�����~�g�"���	���R����f�eK�Ke�RU��{c�cQHݼ����4f��[��������(gK5B���u�w��t
�c��P�;�������Jf��ұ����gǕ���$iOP�)���j�~�_�p��]���JH�ϩ������NX���)�!��/�i�;Wm��m�J1��:���t&A�7��Ҍ��;=4����2�'�G��g���!�偎��0���J��/�ݘJ�,7=|�U�	~y�n��W����2\-?��0+ٻ[�c{�h:���{{���c^q�D�s�9�������P�r�\�\�9��Wv��(��-�]ߌ2ݳ��v9�T*���a}�8�2k��a�U཭�`��H�uݑJ����ӟ�Ô��,������'��0��KИ!�Ԍ���.ܾ�#'�G�}"����$�CUgVf��w���vܶ�����8��;uB�&fl�L�=��Ϫ�"�$-��}�W�N��3�zG�#$k*�џOŬW=�ۈW��8�4%� ƅ�h=��P���̄�Fp[��S�r'�_���D���a�'�^_׿�~�4�&�3?�֡�R�4��`&�;��_���2����� ��;k'�:����dH��f;��A8m2��=�����D9����P?���? F�A�-t���"��#UL����s:���!Dȿ%�a����>�͎ɉ�b�ٌ�ь"фT�`�I�c��g���qŭ8�����KR��q"��я�ĺ�!.Sr���(�aJ>Q�_��ym3�șSɌ�/K����j{��i�x�<O��5�gI���-���>G�x��c�Ȑ��Ԝ��Ø*��"����%M��_�3�D�Rb��&��+�S4e>�b��D�R��tb>|�LB�T Ig���!���]�5;���%g=�j�V)
��K���M����{�������;_=���]j�=z)��r�&g���
�L��JDx���v�[Ln���`��~���b��xF��SSe ��`1|q�b�g�.���ֳ�Y��.�)���p����HC�Y:M�o��B�)�s����e�	���t_Kq�h?$S�I�O��L$4zҋ����C([���`ʊT�d�IE�OĀ�؄�6�!�u�d�������RH�\����]�4#�ªϨɬ�5v�߾�|��Ƿ��CZ8;�f֧�X"(��1D�'�@�
�R��j��:��x��^6���G'V�֦�/���8H6�ȈG���Y��ck-���ߠS��P-C�YtM���'�T\^5�@��xf�����ž�J�1ʚ��'�b<��%�L~�\3�����7��x��Q��4v��67¶�Z�cL�^T���LI�ߝ���po{+��e�n�
>�5�U�~���z3��ĳrm��0���Lg��	pH�U�!��~�k��B'���H�NoD"��ΨC}�c�~s�0rw̸,ɔ�	a��p����[jd��d2Hȕx��1��dT�L�0I8��;Z�"+]��>�6J�F�5��zd=�n#�$�3ix\6�h�ޞL&�LJ���#
r(�������7ed����AP�$���h܄�P91���K��z�d~�/B�"T�#�*6�^#)��G�!?�p���I:_dq�w�<��ݶË3��#)T�Z�>���0\N���B��a"���d�L'��ʎ��L�����aC�þ8Nӽ����F��)��wн<��1\��?���6��ƙ�B~!C�m8���-L�1JA!�:r�|@.n�t�LԌ��	kPW�
�>������A�(��1����+pb�\c�N��#��㤋b!)D� �CI4�]���w�������[d��ec����w��r����)$�I��̈&��,1"��O�f;f(_㶐���bԃ?DSy�t.KD㹜�����fah�h��S���6QU
NY��6#�5�h���$F�u�I�B
�)�7�����W��2�UlYYBJ�d�Se�Dq��(VV�u�~�S�|"����k��D�#�;p.X8.��
���K���+x�_��*2X�}�e��UbL�h���Ւr]c�J�����'����q�%����;��u���$�1��찖��}c�L�����3ӂ9 3x��u��%Fז۱�ƅ�e.�I8rӁ0�'� R���ĸ��L�v�8��n�ȏe�%
p_m�B�4���{W5^�� +2���؍�N�f|m[�����>hƸw��k>s�O>���Mݗ�������zV=QM�,K�L����_w�7�����`�EIEjt�"X]����S:��d��d2���(�4��I�7���o��v�⤟�'1C\C�'b���5FZ�C���rԛ��Z3I��`�����m�[��k$�9���З鄯XO�$�L"z�q�����˄-�y�ct�'����fh��Qa�Xu��k�z!�_&f<���q�������e� �SR�6/97�%iz-u�^�T�u�Ý�$������^B�4:��bt����\Q%�r�|)��X"#�n%��nL�ml���'�d�<X�<k����m��Lk�� �$�
1�.E6ڋ��g��N��a5��t�=�q4�/l�G�ػ�1<�����	��%���9�7��U}e�pʇ)
z7��C���RQ��t:i�_/�����7�vv����XQ��HD�0	�K�TU��1$�dG��Dܼ�#L�'��7�����e�KI()2������0I�C�3�S��>����A�{%9�f�q�pI��UV8�I遳~����t����2�����;����X��BZ�&g��kF�	w��!���_��O�ݙK�i���r�7�z{����,�t����"�n!�R���vo_د�w�e�N,_��L������#h�F���� �HR?��c����O\_��<ݏ��8Z+���G+q��#k�����[V,�Lb���5ӆ1峕�̌�j�f�`�"��63}���7�vRܩ�~���
��#��Kf+�&����}��������g�gH�%�ȯuu������_�b6��!i��U��_��\ �'�c�7~94��{��r���,'IґoH�H~�\ g_���yFbМē��Q��� \v���H�W�p�(�g"�ŀ��IZ�z�����d>���w<I��l�Y�ֶ���Bg��E����8�>=	��Ǖ�7�NNy�&����<��q2%|pc��P�L�������<���C����o���2^%ĔH1��au�$.�A:K���{��jpe� ���1z��H��>�\�@�D�P[��LT�]O2�͢���|�(E�g�L��u��1F ����"���.5��bu�X��4R~��4�7�DN}�G$;�������:1��x�H?p4�'.��V�zm_QBN_�4�^�Y6G�>�K�-�+��EZ¨'X�5��`=����j)��LL�.A�Z0@U_KaD�2����w�0��Y�2�
�H3ńv8�x<�;ke�(���}���L��~~���or
��]:��(��rOG���+���F�v0�2��a� �0d�����#QՋ����	"����҅Ė�o�8��L����k$IAh�~�rt�*!��)<n�Ʉ���Y��V�.�䃵���w��E������w����KK8܆+����^ �9"�l#3�����!.KQ�"#��x%n���%���,���aQuPq���^����3�%P�.�%3��=Pl\�h��3��������4��!�F��f|}�3���7�MNvyI6����������q��������XCҙ�9��LFhϗno!a�I�$����,��[�A��+���e���4	6#��&d������ix� U�@��f����扟?2��r��tλ����]�����֓/�9[=n��EZ�8����x�����8�����,9H�#����T7@�h,��#�:�2�4�P&��kKEM�!B3\4T�0�OA6�-�"����8�^(配�aa̔7W�7�I��/s�g"�_d'�K�qd-HI#
�
~��.��b���a��7�	�r�;(h�ce��8��1&FH,+����_�S'Rm	ee�&'�'��2Kl.��� �B BQ�b��lݣ!X���fW3~v؈m�"K�X�V�����Q�;c���x����5�4qJ�ov��U3$�7�~B]O�4�u�i/�������(���3�r(�2(
(���.u�	L`��jw�(��Յ� I'�7�N]��H9p��e��H��[�B��s���ПH �`&������5$�QӺ�~f f
�R$>wn�l���$�w��Y�CS�����7��u��zq7N���sU
���4����4��^�/f�N�,�2�%��R����Jw���q����+�V�d��M���G�(qZQ]j�?�&bi�ȋeJ>¶�l�}�C�1�cG�-�~dE�=sQ�xk�)�#���>���Տ��{>ݾ�3���su�&?��<E/LLV�kE �=,��xN���z5���J384Q��Z�J����EN��#���H�p�����'��-~?�+����D����iY���k*A�ߋ=����t;���*�;o���555o	{�h᧲ m#���&����n�ԊCc^C𻟫p���8��+�FP�8�2����8�����b�mm�$#��Ĉ��0����{:��'���7� QLP_IA�헣#�ŏ��e Gi%*Z���G�G>��y�z;�	�L�����aם_��)�EF4,�4؆a֧�d̈́L$���^>��_���s|0R��&/�$�J�W�jpǲ�k�y�:Ȕ؈A���_�Q9"�O�k�o*Zu�2��9�7�!vSѠ��{�=�\��~L�9IM�3�u�Z<��~<��������g2ښ�[� �����{�RgAsc5�M*x��N���W���i��bZ>���7����v�6��7��$�w��¾o�L4s���j��,�4�4�!�H����H��63Cb\*
N#f�D�͌R$b�T"��
��1�µo����[w_�=�{���s��Vxs�����T�5���q��q<��sh��c׮�"(dGΙ��Xi���cU�B&:��jo�'ު2�M�����bi�,,%s	��[f��� 7l,N��Ŧ��_���pى���L��C��v�|���	{z��x����KX���'s���c���������@ |�	
�+�QU׌�����b4�FcE�c��%r�/^���@ʊ�%)y�M~��b�y�-H�G�&�gK)�d�0�ݞ�F0c,pp���!G'<b!�h�We(qR%B��0Q�e���90J��5���R�������|b�C�A��=F�*B_8����B7I@cL[C����X���)lru�n(��\֥hoɐ|%��F�/��4�j���ʘ��˽���5�n���)��_�v���|�0�#N�MEЧ��r$p��J��N�i��L�HP��gUQtk�}J��\�Y�Ɉ���"��^c��y�#xO�A��6^T.K�h��vc�E�7}P��l�Gއt���ԋ-c��F��@m������y����mp�S�L�q���k��ヷ� X��M9$*��$P�%���$1�����$�+���KIc��D�(9[�;�X��6��n��8�������
]���Bľ��h=ǃ$Sb�����ɴHZe�ʑ)_LĐ���N컘{ �5���
,&	�N#�&���I�PlU��e�X\d��eV���p$:a"�[Dإ���5F0�닇Ajˬ�Vp�/�2{�4����2ngl%�Iv4�G)����l5��b4QN�V&���0nl"+**�1ia�}�Q�6��-�]Y�)\JJA�UoI^;n,1'*]�ľ���+�Ӏ�d�X��5r��nhr����� ��9�c�Œ��XW��*�ݶ~���Q��0��0a2n���A��c�y�i$�Y.:L͐���e��v�0~����gztpИ��0��?{�<��!L�c�*|�+p��bہ߶��=a��\4
�F�o�n_�qST
��䱕$"k�a!��8Aݞ�Ǽ�6C��{�k�����zǔ���J��ϦSf[�v����<�4@b/^���L�3*�}c��/$Vj�gq��k�Sz��T�cx<��Q�����4[�$\���r�L䩩)��o^���9���O��"�6������fKPD�������9渓`kr�HU�Yά>NH�q�0.J�g$�%�Kz��y~{X.o�WrN:�~1e� E�SW���������#���J�%���,��:�P�B\���F��ch�-!��
�Us�Y�#���Ήq.X+���� �eէ��=�OoVQi9+�~sBT:Ie�Q��OpR���g�D�>�P�r�TF����!8�iT�g(��R+c1�X��Z�D$�H��b�Ia�I0a�1bz8y��,ք���8�4Z�7�@r�Aɵ*�beP$���"���êH�\������t��w��Z��N �U�,�l�k�^�`�w
e����(���Ph��St���u��E���iܶ݋��EB��6:�"�E@W��Ś���}/����')���Ʈm�s�|��.��gHCJ-	Q�2nN��6��(n��^������"�g�y��`�+9�T�%ǯ#Tk�-�����K�l��G>#�'%��u�˫�02i k�,�
�'����5g�d�4.s�� ��IZ`$ع�݇'M�Kw,�x����at"�����s��������%n09�0�-b0�����nK�\wJ�?6�!�l�_o<����d	=w=�j�4Ӧ�����S�9x�;�͖�� n-Wa��E�(V�ɿ���\_&*8��ict��m%���,D�um�C��2��m�+�="@6�#�!DD}��ؑYt���亲)��RoKC�ȫ�Ӱ&��٠F��(��0�ּ��o^�t B�̢v���Ҵ�tm�ʔ�������r���Y'�V�j�v�y�!�Ru5-LG���n~~*#�A����5tn�ԗ��Dr[�ԣ�x�aL�e���e��QK�b/v�����xX��(��0�K�pKde��X�ȼ��rFM��-H�g/�B"�����T0�ȉ�����Ag)Ǒ�*D2f�HQ\L����|p�v���xn6����xn���x��$&y� �JG�Ba��Y]bJ��$�΁�*� ��ݹ�5��Lx��ˑ�O�Ł�;V�FGD�	�~��F�I��[��pII·ӄ��4�(���S �.�A�⌰8�o�Ҡ�@�6��===-␼�Y}��������N����F���L������ck�q�va�pSq��CN�+K��7(8Qm�����ϝDW��
Y��v��𓔯-��W��g�_0�I�N��8��C����Y�.v�9c6����:���~Dɒ�2UlǷn^[���V�&H�RB,B�N3j��E�L]�VL��!�w�80�㏵��/,A�u�;�JE}Օ��b=��A�^�Fz,�]��S3*ڌ|z��j���L�"�qs+��R�&��T�p≽���_�Nǵ�����j�.t���φ��"A  @Dψ��XZ&�B� �Ә��V�j��6�XNZub��0�kmS�-
aZ����l��ͻ��\�t^d��?�u�ia҅K��u˨Z��RU�����\�D:��8��v$3l�%�(��0�#q�(psM@2����$��8#	�f�r��x^��ΩI��\�F�� �ތԖ=�h>���Le�����<T���C���+��������(�	��:/i�*R�ٙ"a�6�o�?N��],`q�PgG�X�� �_�$Qd��B�e�:ǙNPVM&cŉD�8��q]������K�zƸ��)�,+�ۡU���<wl ��h��{v��>O9DJ�A
�@L�W1��:���8?O�8I�pĆ���B���%[�|�^�T�a0����'Q�\��Tl��$��(��4I1��K05c�!�!U����S�őm0#Š�Ɛ�:����D|E.�L�iY�a�3?�m^�(~z���5Ý��Z�y���/Ӑ
�w��'����}߹��jx=��z�+�����j�������my�p�_{���P�A�&�Rh2#�x��]9�I(s�Qi�(8ס�4A�-�dR/�.�K�s�LzYH�L�w��ň"�-�4��V�o�ׄ��ہ�����SJh@�_p��ky71bd eŷn�H$�3�����y�����K�45FL�go�8�Ȓ�+��&���Q�����(�Hƒ�t1:��ڤ8�j��6z�$���Ox�$�	��R�˖�Q�0���ز��$�|B{P��BJ[7.Cs�]���T�A>�-�fm� '�\:0��巔\Nk6J'�]e�G�S+f���%R���Zg����wO��'�a�wm�S��K�)e�Ec�5��#5x��Nd�=V��3�
�91���H3O_��׹��a9ce.�Y����=��fB����K��3�~�h�_޾��	�Ə��"�'��.���w�����Z�FV��W�ñ�F�L�?��$�0�SW�y�,޲�%�����޳�B�b����&m��ߑe��Xf�'�%QXH��)h(N���H������4��j �,.q�ǹPU�W���aL��p�vyO�����;���nE�z����+��'�^ۈ騂��� �|����o����
K���ϡҒ�$��=9�ud���w�d�����,�Ų;~rz�`IhB(�C\�
��VƓV5��Q����1��-�p�U����Ƙ��;tُ�~F�$'%���˨F!�!���40k�2"�@����gH��7���Ë�'pm}?��Kb���:zK7�C��S����:e��Aq iq=�ӆ�d�_��~�i�=��Q	]\����ѧQjW&m�u[�ӼJ76c���|�\�o?q�'�7�hy�:�/L��SlF����|Hp�ԡGK]�q=C���X]�d|}��)Ǯե�v[�i�V3WЏ��q0�����	�=�΅1�⪳e@��Xd�_)d�v�ˌLF	WV�X��JJ��1Q���U������e���c�5��Ft],d4f˜�q���,*<���E�5{����M�`���\�f7��HdM��N�x��)iKk%���"f�M�.}�� �NtZ�\�O�-�����x�@'^;,�kƱ!��`o/����"���iF�X^c������k~�5���N���1�����̹��z}�R��re��:�@|y-�D�q�z(��`�q�D?�yr�@a��P6]#tW�+��xN*<�d�Ro������ɧ^��{)b2`7���$n/E�i��(A�Z'T)zB��׻G�R��V��Q�����,�#��x�Ss�{�Ln>���\�$�;5Dc���n����0���N|��Z���~��/�=1��_��~��>��&�y�U0��5%�d~�2�X�H��`*@o|}��,捃��Nۜ
��%_]��%SM�q��"��Z�Y�>�wK��0D[��\	"�|kG~�_.^2�L�ĲG�Z{J���t��W��NF�v��؆\��*����C3ȕ�KZ	��ioz�l@l���_\_�7�8���ǧ!"���h\�<�����xJ��WO�s`
'�"h,/��h���HĈ�i�J��(���MN��C��T/��Mp���h����C�P��� ���w*n#+�����@\8m���
�k���ɧLFf;���=.�=��RBp��>v�޵�n���4�O����>;t^���}#��r�E��x����{k�ǂ4�/E�^0.!�.K6�K���$�z>��ݯ�y�i��M`�c.Ҧr�o��?�	��x�|�O�DOd���^?���Mm���[c}�O���SL�',�,���̔���-8�L�(�`�p±��3d82WP`7��R9�+���3e+ó$=�0?��̌�v�ra�_�t�	��&~'J�MJn�u�=BHk>Cx,�ʸwx-6W���d�����t�r4o���y輂���a69��!%�*,)�8��ڡ��E�����L�l94�8�K�d���|r���V��\�!��c���4�c�ήS�;z�nK�����#�jN� ���G7j��P��2��0>������w�^W���F�`gU8�1L�S$���:D���C��v�.��Y+1
�b8)W 1�T���:�J��s�s��؄�mҶ�+*o}L�bD[ʒ��k�<c�p���,Z�>�N��|N�9�<.Ac2D���{�뱿��*;��1<v�V���2��u(oZ����,��/R�u���}7:E�h�hK� �^w"��˖c�GC9o����AU���o~�NP:�,2d�����{��3�6��t~�H���$�*������Y�`oP�mt�E&����2'�-e�%?���A�D�����M2K�4f��K$OEt���'�biYR�Jp	�H��<~�Jdn��Ý?lkv�ؼlJJb����}��b���ֳ2��I)n����`�#��H#����ȹF<�/�y� `�|��}�JVN������Q����b]�S�5H�r@���3��z	>�/��p��sO�=�\3�ߘֈ)���躹L���߸����|�'EI��wH[㟡k�H���5�3,Ut�4ӭ�g��l���:�ź��f\�H�XC�#q'!��B�9�Z��I�	��ȱ�{�Pl�k/�*��H��ЖE���9�ǻ��F)Hf&2�6��k�Y��ɲ���C�la�x����-��Og�    IEND�B`�PK   $��X�,͓�u  sx  /   images/7a575584-996f-4f1b-8f01-a278e4b2f0d1.jpg��uT���9��@���w�%�Cpww'@pw	������=��|g���޻�o��WU���tu���m�m�^VRF 0�wޖ_ ���i��_CBEBBDDBGAAF�D���@�����}��������=�<|||�w�DxD�x�x�y¿{�А���0�������
Gg� G�ǁC��{�P  pHp���-�����߀�� x8xD����_��~ "�G1�*�(T�x���<Tj�|�?4\&NAh��D�$�t���yx���|������U�������cjfnaiem���������=$4�GxD|BbRrJjZ����¢��_�u��M�-��}��C�#��3�s��K�ͭ�ݽ��ã˫�7�w����@����?���<"""�|����g "�Gd\1c�T���x�м�4j.�|�?�4ܛ�����_�����r���?|� �p�^@��3���Y�V z��G��O�9����>c,}�,v}!�����^���O����^���
l5Um/�*gFͮL$O%�ƈ�f�h2)�#9��B#��C� �B,���dl*���9�?���1rR�+�:������>�@��S�~T>�ӯ�{�}�9�;���H�e��S���>��
\ݯd-�<�@�zꏚ�]{��x�
?�g����g�K�W��>���^1rI���wi���Q�L�N,���S~�(_b6�f���?�k���MG�0wc8ń��ȩb|in�u��X��*^=2�vp�*B{�k�=/I�z�׬IB��2�f��t�������0����$�vl�v(�� ��|����Tf��C�\��#�}��S�|6�4!N�ġ���y�<.L�c��M��kW�����G�3���Շ 2A2�ٙ�pVo �
�y2���eJ�/2��a��q�x�RtT��'6m�gx"S�6̞Z���,��.k��b���m��t')7r��|/ip�Ɨ;��y�z�}��$Kw�_rE�-g� m�!M�t��v��a�RLv�@�¦L���q+���/L�l!��|턘	tEţ,�i�b�1�1�F��+L1EY�~�d.�n�/��G���|j�\�#8SK�Aj�S?���[�fݳ��x��r�Hx*��j@PӮ�U���I��TpYk�h���{�_�����Nr�Cc��a��n.��g!��������1���J��8k������c<�7�k��f��>�e���m[��RM׈̸&:bi�M]�޻�{R������=h��-��9��!�;���F���mw�Gf/ׂ&��lM�Z��az���"rVO������F��:q����Z(��t�=���KF^�y@�k����4��	��X��@�B�AA�dU'/����� 2ﾦ��h�8m����_��� �R=#D���kI[�|:<�VM��C�H�M�&-���ߝk��x�F�>�>Iq�m��ݦH_����P��͗�F}��]�$����aއ��-����-�gXR9]$����q�I�0!��p7\θ:ә;���uY��v��V&ؒJ<=�jV�����b7Iw�g�?���/5��
���re�(R�c,m�+��eX������a��!�H�y���ڡN��f�j��s:�����aX���H�	F���.բ�Ck0�,�̉��S>;ۇ�����5��y+�2u%a�%�lD���1��ދ�����̨�Mv6��(���ֶ?IK��iۓ�1����v�������
�OS�^��Uw�=ɫ�cĹfb�\�_Y�B6�hO4���i�@Qu����Aиn�8��2SR�b��Ah�T�����,�J� G���>4&�/_�?l{�N��u��sJa>+'S#
���56�@v�I�iq��ҩ�p�d�2��%��؎�f��QE�k\|O�H��Wr>YfӼ;�}� �S��j�}�{��ߓH���8��d/�l��+�	�b��B�_�nٷ�걼 ��G<T�wI��R��]�7��g��̈́ٽ��DG?�;FC�J�'Ӂ��7@�Pd'Y���R��:�Ll��kN	�8��?�6F����vąR�H�~�/S�b��]�74��ള&3D&|�]��n���dnWJ��^�!���3�Y�15e:^�/���!��_~�fn��|yG����NO7%=i�A�J�i~��Cn����߇���K���K�}g���/��(U�Y9�ݾ6���"]=miT�dA�c��Z�,�2-�Q����C�]����B#�:G�d�$+�Q
>�~�8fE��5�.1��D�Owkg�����6��>�f�*�F�6M���V#�E<k���[T���Uzײe�)B]����y�-M��M>����0M#�hO>�j]�bbO��6l�:ϰ�H\����j�1�V�R��������k�7�}����̟
������ɕ0q�}��*۵mg2��z|h��lu�m�.��.p�K'Eqڌv��m�W�+.(϶3�/�>.͹���N��F8M�/������P[=q�k�ʙZ�Eg����3m���Vm=ɿ�N]���]���}���y�b��kU{=�������J0����E��	=!!y*���(ђv�u����N����<z�Q�r�V�CP���8w|�=V��w��2�[l����Y�]��U�=����k�y�e>�ģ�� �}o�����b�����9����=��+Q쪒��Y���͏x��'��v���6w�k��'����8\��E�]��*!�����ڇ�K,{Ʌo ��"�p_
j*�/.Y��D���)�U�~5������[d�\�^�M�4!�6|^�1�9x�.uQ��� 9��nbۿ�6-}�z��H<7'q��NVx��B��{G���mG����JO������*��;�S&͎*��G.
uΚ�@����\z�)Wvϥ�:뱑8��äM�7�-})�|�f�R-PAW�y�#�n?�)6K�@�̩�9K^��p@-aGTb2�GH_N>kP�����Ed��3C�F��N�'QqeBv��dG��O�]&�hf��߭��uf��+�����e�ˠܥ�V���MYV�S��{����.�0�J�<V�v�ř��ŋ��E�+��#���SQ�se�a�a3e<������zt�D�����0t�h;�ڛ�����uhM�8Q�%]^�&`i��\�Ǎ^�h�o{�5���S� �ⴘ����ӓ�����De����Ñ�?�˛��:���W�ܻ"��0��V>�V�V_��(*_��<ý���[G#��q&�ZWk��!�\"2Mզ���@��ZB���m	�~��kKf).b�Q]�3�����N�1� 6J��B�M:m�K�^kv@)�����"�>�=׷6���^1���Y�D�KI�)ꩌ�c��I�֙� ��;!"�w:7�<ų��`W�YV=�w
�����������O��W���	�s�gC_ҥ��(�A���ː����;�U�?�\`S��YK�]g��*}зtbdU�E��12ۋ��7 K%��� C˿��,�B����E�m�H_�	o��Xj�e W���D���DY��\� }��H�]��L��>S/d8ކ�Җ�?���u�!��U���a3�St5�XpQ���3TB��!a��`E�"���Q�ܬ��9�4�
U�'i v���C{e�`�vV��̩!��=���?�E�=����)p$u;﯁?��cd�o���'��?	�[��i?��7�}UJsY���y#�Ҍ%ҿ\���{�3Q�&m֖<�K�kJ��cX)��v��d�+�i�!"�b2�YE#���2��Nijen4��J�[��2^*D��lˋ̶��dA\�9$�)Y.B����q��X#,'M����7V�;>��Y@?�j@W���Fk/���s�8���5��������0�uI�u��d�@�n�8Pt���ڃ�JѺ���~1��Wf�mؖ��M��߶�6��*0?���Z��B�Һ]�$[;���{t��8�"�"��n��}Jsgl��$@	�*�}7�[MR���3��e�&��,�"blPǮ���q�vU��R�?��cm���s�r�Mr�fJk�<��k��i�h�̂�+H �)�7�&��������4��&�)� ��Y^���=j�^f�%�T��^�|�}�Nܡ J��ϵh���w/	%Ø\��NCVD}~�t�yϝ��
�)��gz�$�?
b(�!�~���E���D�M9�1��1�r	Yg�ϭ�~������Ȼ�kV�zG{�3��e�(�R�q�5�f}��:��vB���G��R���QbhQx͟�G��ѷ�  �8�t�g������ѱ����
�b�\��Im�T�T �C�.�b�&�z�ࢲ�t��J'�Ǐ�J,��Uq��~�N6��D��j�~�9Z=�&�I��������9�|RHq�2&�B�7�(3HD��=~op�(�^ф!n��\���}bm�X�=��Wi��&n/n���pK��?B��5��/A�B����E�k�z[�\-^�ϋ��(�[�-@T��Ɂ��̖�U��4`N�w����<�-c�=CK����٠~yaH;�F�&U����ŋ`��2c\�?��M�t�Qi�IG�v�TT��`��m���o�$�b���1��F�P����$��k��%��,��;DpO
�[����Â�!Q����$���g�E�s�/q���h�`�a��T�o+u�W�w���?��L>����|јȧ�����J��	�
uU+\�&����6��<�*��|��̫I(y�������?��V��]�7�7�>��2.Ϥ����=ކ?{CǞ��#�>?�_�Ĵ�X��,�z\F�g�F5�2��O	�?A���j�����G�o�"��6ٖ�6�͍�<���p�����V&��e12+��!-i�QP�Z&�^�oR���P�Jd~�W�<\+��O��P7�e` �N����Z�X�O�����������V�(CS�0TR˄�{f2h9x`L�Ccm��)��������c[��lw(ʮ��T�=ɀ��٤�tXT�� ���3J#w��з��,��կ�u��ȟ�	���
w��
E�]8�%j�,�кĆD8������AC.!AT-��\*���)��y��J�ey6����gM,�ĐyĹ��
����}����2
��;�ma)�W_f'����w��.�I�ޅ� ��'�5����.e�y8���G&4̏�����h㷃���OgS�h�m�1g*X΍��|�<,uE�-|���=)�Z�Üi���d��`�>?��>> P�˪~Tcq�3�h��#V3qRW�lz�`����r��/Rw.<RFs���;�ND	�Y�[�:������Y���,c��F�3x�*��$@k��P�m���#oZȰ����S���T�[7��@]�!l4xoh�7[B��^� ޺�����Tj��Hx�yW&�>B}����LY�䍚m���]�!h�jȉd�I��l 7�#u�}���`��q�;Ye�JY+���
{]j��+[�2����d�w�7m"��:�#M#�\�'1��|���^�I�6��Џ|ެ��Hf�Ԫ��{%:�8hqxx��g��eu�x��)r���|��1��J�.D�#8��wf���	ӑ!�}���[�kt�f��t��J�8�w�A�hc.�L�h���?���N�Y��D&�}H�s��i�s�w��$+AC(Lx�:�P���'3Y Z�����Eh:2��~9I�Z&}4�م���}Yӟ�Q������"�~v�~Gjê�n�M��0Q1���&:[i�;�%ݨ�@o9Xw{G���i�s��6/)�������yju�Co6a�b='[�L�[v�+�h7�����l,��q��I$���O6l.c���~�I����K�Z����_���)�4�4n4O��V�O�#
�.���Xb'��ɑ�#Uf�<ɋ�-���W�L��������<9��:�)��e�[����B�]B]̑�4�%4Fh=#~��u҄��o��!t��
��,QFG�(��crr�|^}�1��1[ ��XL9;��t\�D�
�
�e�� .�,�$���GKNk�>S�*�H����(x�� ��x��GxB7��I+��}�=���]W�1��}���U~��Y�[���p����S�o��m,�G�)4������&'O��+L����f�B3R�A��W�p%��7����*Ũ9���dX���[{�
7����j�4Iд��E��ٶQW
v�oᳬ�X{�m=�7ڣE��[�ݟ�X���G�L����Jl�r�r��/wC��s�i;sJT���\�Y$VRi�(�Zgq�T�ͭb�,��k;�Z&�;��u�����R�n�`�-.�T���(l'��Z����T�,�U�7@�@	��B��c�e/�,<���HJ�>��A4nc�a!�Y�����@�Wa J�d�ˉ&��'�s�LV�\�!ËϷ�D�?,-��n2�X�rCI��4`�y�s��3R-3��
aQ�M��l�gE���#X���dB7���@�d�������U�M�E�ن�g��n x���#�P�xE�]覩t�2?sS�m��Sy�m�w 0�J{T�a�ZV�ML���m���KyU_�,CN��r!
r�`%��u@Va��0����x4B3���@ |��P`X��:��\|C��R�"��\z�""����3sx-����P,���D��P^�S
.c�Q"�\��}�׺��,�;���% XAkgs@��ܨ�H��!��J~�sɓ�P�X���YK��6񚝘6�@	b�@a�I��~�8j`��yb�Q�λ��3������Ex�ı��#���9�������+�K������,S���J���挒Ɔ� f����i���~��j��{��������ǛVT���F�af�MYe�b�����D�r��
4ac)ݼ�1i�'M�����",=#N�ԹD� ��ֳU,�p�$��]dE'���y+"�@���>N#�'?���r�٠���vYi��ؐ�|JӖ���pg�h�g�v��R�*Mmg�f�n�ڿ5*9e��
=�[&�\�ƕGO��~�@�t�?����y��7̻l+���ޘ|�̩՗tg��yK�ү��#�<{�ӑs��'�8C��X�����Aʉ� .¡˴J'A������;��1���(�)\�j�W��#��u�_n��TAL�Z#�������p����q�!��3n������zڻM' a6��k7�[V(���Y�%�0�蛣�2Ee�3���9ȏ䀺c��Nsj>&Пqy��֌�X	F�T��YO$�B�(y�?����Y�����+��`�Igs�<�;A�eS�4���p!��.~F�F�p@��˴�����z��g(�ۍݰ�I��ɴ="�*a���VkM�Q�AUQ�\����|爞�w�n`n[&��� 4�;~�%e�����V"��mB�.]�)��E�".C�0=�eJDj]޽*�"�L��
~8՗A����Chd���j�����H�KGz�&�49/�CMT�;��L��R���h~�o��Q&�N�\����M�P��(�����w�L�6�%[V�.��d��9o7��H�ѽ"yl��������/��#�ۼx���W�Ă�4��ĸd�HHi��p혹p��i� ����Q]�dOK������].E�tD�dӯ�}�0�Ć�,5^�Bh�A#>�2�QI�!��Sؕt���]$�?f��5�	�<^u���団�k%��@�������_���5�a۪i�0��&�oj{�OzG\z��T�(���(�o�`x��s�p�U��i����i6r��W	!��j�:oNh׃��f��zh�$1����K�1�� |N��Z��g�U�^��˽���ڥO�lm򂶟���]��c4_�*���(C�6��RX50�Ό>S�F㖒�շ�a����m��RmuFe ⧎	��[����e�\��a��u͜#��:#1E=���N6��������`�
�&���.��ЪX��MfDwM�|At?����5a�A�S_��~Ǣ���^�t�z��!�Qߣ��Ո.gL|�5����b#�2��~���xw�v�)t�'L��B�Z19zQq\���-&�n��g��R�e�i���b(��s�����q�wL�+��{���u��egWCc�	"���ϗ-r�ĨJup���c,�+�%3� ų<5�����o2���S��W(�)�S�g]���@�O:im��5�.^fg��m#�Ը�Z).�hr�äh$���t���X6�[�cـ�6��c�B��$
M#�������2�b�b7��G�һWS��-1�ޚ)@f�I�g�^O6)��|�SxT�ۥu��<�����'aF5��%�����휩��� �x@���U��R��T�p:�J�������T���du!��at�)�ҏ�k?��F;I1�6�m���GI	n���r��;���0�`���q�b���$ܰY���-_k`.����koܷp�D��VgM+�pP�,�`�*�J�{W��/-�SQl�J00�yJ���f��Ƌ���d"�-0^�72W�<��D�NR�s�t|#�������̤�4��uĥ�kW��D�D��{�~�9H+�0o{,�)����S�~	X��*�NfWP 8K��{�G7� ����v��r�W�3Vւ�0��bW}����i	�n_�Z�ρ��W;&6{e�E�CW���
�*�����K8�P}�ǧc����X�8�,R�����|��y�Y��rr8����?�'�R��kم͸d${`��BF-;�ؕy��L>�+��D��J��1v�Oа��kv�����-F�@���/�
�_�q�M�B�h��M_G���Y;�|����Tq%!��^��Snj+�]n��y�~ �cq�_�ZѶ@�r�I��2H*���)��7'��w���x�0�'�R�a�9�}���H6(���)�oq�T�K+�$��Sd/���]�,l��7@�O���Xq��P�iw5��%4c��d�[Gڹ�z�p٬�wVVw�z���e*��J�a���a6g٤�I K�#��w��D����p���Y�=^�!;ؗTb����`+ئP4��+�ajL�a2t[�q�tC�΁��?:� �7QP�Mqx��|̨X�'ʼD�ȧ��r?���33%Z���l��bLTox��h;P�8��<י���ȟ�J�Е*QحW坕��w`��ԗ@�����o�[7�ߤ^�Fsk�k��� l����@*�WШV�h�!���A%��I�&$�{�J���v������<V�ҿ�����ܑ�h��#+ۣ�-iܭѥ���KQ�yF��'���i��=����&����݂����j��C�S�F�G�z
�&�M��y�,�V�f�`V���>*}��H=V^�G�m�kw��3�����DM��#J�=C�!����\ c*
���}`*�X���29P	_KgU�$-u����@%��  @%0�ր,{��K,zbw�n�q��L|��� i}��a:��s	��8�U=G�����FYOg��&�=�k��$��+R�X�Y"�]U
k�84�����]C�=.~q�z�9IGG�\�*��$rP���k���{�����3r���O�3�o����`M�oU��V�ۃV��y��E��f��{�x��;�w��P'2P&2��������pm��i�Ӈ���Β��&)��S֛��>w<����;\���1���k/3¼����$b���b����ap�J+ލ��̇g+��I^����V �h�DY@�%Y�sR�P�H��?��D���`u�m.�Ȑ�B\Ʋ���!@�&H=<zZl�I��P%nq0�}a��p�V�����R&��	5�-w��T�[�����TXL�6�mƱ��q��m�[<��t����7'@� �AK��T��l}F�ߕ�ӭ��n��e'�F��r���&�ĮX��t�`z�mTB�Gm��H51���*J��7������=�TW�L7ɯ��
�*،03VT��x�j�cr��� o��F��ϟӆ����px����6}l3��<�gf�9/���:n��)[�����q2�J:���jl܎��!�z��c��U�m}^ݪ���1���\j��$��m8:M�  O���uR�
]F��>L�b��fF�n��kɘ���'z$,��ՓϿ�A��2�ki��v�a��<�gܤ�U�胏��S�%��'��3���ʢwo������|
H�˶�W�{���_:�jҮ˘㗞OJ�ƙ2K����1�#K��%��u>l��b��.ּ�W�?��:���s ����2(���5��U�M��{�3�H���+�!~��l�ɫmz�|2��5��V���& �E#`Sfr)�A)Y��avp(@�c�������L	�5�e�1yN�A�HG(� W@�M��l�^Q09�2���7Ӎd03�(2s��g`���m��0�T�շ[Ep�Pt����.U�pʡj!��k䁙�L�3��#M�B�$�cn�#�J2]ܔ����d��,'l���S8N�wm(ug��3��Ͳ��4:�
	EW��|F���]p%Ĭ��*s��+&�^YxI�7_5���~-��yuC��ƨ�Vv<�(�6����o�6׃���:3�&��+W�|-�1 �E��W��w�~��U�`kte�{g�m��V���foNPJ���Y�/䙉T�6(P�)bU^�Ӹ3 �x�����}x�5���������d`d	ww���oڰޅ�b(L�������MA����c���͎�6�*C���Ǳ@^�$^��3��,	�$��*l���8�Y��)Z9r��I�E��*�����}.�"����ٚ�޲�����%��J��xOP��} ���\�~�(
�rF)>�-?h��0�BPX�9���\;�|�W��9?(-��q<(��,�E��ٺ��I_�l.%��ޣ�����O~�p'�h] ?�1 �O���+�h=*�ÙseL޲$Tя����T��b��f��҃<tU�t�DT
�(�c�|
��G���-�A��G_���2�Tz8]˴�~��
/t��sE��<ت�	��Kd!�`f�%al��⩛_4<�Eu}��RI���Q��[��#�2�`<Sa�4W���?��r�9��Q�?��~U�M?�Yp1�)��G�ּ�5�=e]���@�Ҡ�� X"���z=IHK?;pR������9,�vd�A��t��ء�	�<����&�88�����/�-f4�*�1�䆟k^2Jơz�!���JI��K3��� ���.o F��;�N�a��Oa�BX����e��)�ЍR.� ";��!:���_���j��� �F�B{tYO]W�:Z��zr	�Y[m�D��E]m�y0�v'��e��I��_j:�^�P�֮﮼��T�24�^�̎Ԁ�����`�j�!�{��ʼ�U�B�>�֮��]�i��&y$�� ��_��Qd%�6)af-j�j��g{��@>dYZ��	N����T�F ��!G��j�r�H���2^q�YO���u�3lĊb�����m�'�+(���#KҬʪ���mdFhS������s�C!�`��mwh�L%����:����@�ƃ��t�t����֊q,�nm7|��$���>�����i۳��2����P�0_�SeƏ����:)��1�*�d~٬��~�֙QS������R�b����B�ǽ��D�I��P����*�T�0v 5���F�Mq��1�G��j[k!/R'����#x�h�#��ͧ>��$zl4F���d0�b��鸓��4I"���V.ؚ���R|�H����p�M�	�iAL�i�����ڶ�q27�_2F�1 ��j�e��ZN��nsNn�>���NmLܴjl�V$����Ҋ��e��'u1�PW��kcO�7_�d/�b�m+�U�ËV)-f�P���r(Z1��e ����S�zG����s�8�C�񃖺��@��� �x���U$��$<2˘`LA���T���CW��)K���^��N�����D>���5�s�;~{�wPb�4�*��d���b�I�9y��bmR��4)"x�[b�qp�9 �:*D�&��Q��m��&\ن��!���ZR:�˲4�ԑ��0�U(; �9jT�e�:��c7�`o�,�����YnCn+�Q��־��t`�;��Ԝ	�&OWն;��h0{��Z= �S�
6&��>�	�b��+X�r|l�R��ɋ��8NԜ�I�R�?Et�c�yx;�����Y���n T}�I�y$gjp%��B����WL�bD|����N�}����Qü�o�oV/�;����|�m�
9�M	{!��n���ڢ ����|+s������	��EL%,�:eB�;���� ��� ��<h$!��l��#���y�2ֈ�e4G/����s�N��#M\�֛;�(�W����^m��]�>�7���f-�K�,%��!#�lʻ�`��4v����������kBR��=j�,���2���m�s�h��B��ß[M�u*}���R���B���)���ьa˷K����~��馌�.{����R\}��(b���9n��y!�2�����Ͷ �ܔtҔpdٔ��e�>t�[�*bX������W�O�_�rE�=��3Ξɕ��#j C�B6ս��m�Qc���m	���H��g��)fIb>�B��J62�@�9�uh�Q+��4si��c�=�
�l\�Y2�'�i�@��)�L�Rmn��@�^�`>���u㾀q�ֲ"��_��7����i�S�ቂ��¶���q�ЮL���Exs�X�W�&�vS�[Ä��K,ѡ��EE�-~gq*�e�H@�#=��FE��o�}�̷%��*㿉7g�C�Z�<��&eC�(�BO��.��ZHlcY�/��H���icNIU@�!������U�P�i��%2�<���P��l(���=�Lun�i`?mh�S>֢4���!޾�kn�4�Yz|)3���N�0<��d��� ;ZIH�I�"맏Ќ���`Q��L�[4�*�sl<(�v���_
�Ǝ��8����/$A��oƐ�q�&�	0��Ax�$�j��T�zf.hib����!�(�� m�Ϙ�1EA�R��_��PL����cӡ�Z*W�O�����4���)�ʛ]�c��'.e�6οϿ���+��ɷߝ�z��r��i�q��;5.��TE|z|�9/l�S C���ϵ"�Q�3��W�NE�z-���e��8RUǎ
��.�VAhNC�HI�NFd�*� �g�x�d�ч�ςZW��%�B����E�j±�3W�(���zm��>x#�n�_g�N��1N�j{t��~�&V�64c춀�+��`�3�7�S.�Wz?\�t
�kUv�5�s������������23�E���噢�X�ad	��)�%��j���N�]�ٴ�u���Q�o�7�wɐ�ͅ{��98O����;�a7� a��d��i`n�Ð���]&�8:��^v=�$�E�eM�7�Q�Gٷ��4����`��m_���܆G�c�L��{�r�����Ĵ˾�
����x>_A�>9��`i�x���!�z�y�a&�;M#���+���� ����S�S^6��}|���1��΢,�o�����(�1�LZ�l�ƺO�fT����U���qq}x��&aBϱ�/�3� �.�X���U�6&�p�P�9��ZT��8@��c�a���YH���@�I�!�y�ڵԺ���ʆu�~��2�*� ��H�]ՕFӯ�V�V-0�(azL+����%��q!A>����2F��5<���&���m��q6���3o��^�8�C����;x6�>(H(@L7�����ʖ���_#�m��̨q�C����11�컑y����A�S��c̈�佇�g��%k*����e�����%;�:0u~���l��h��v�26����^��ƅ���c$�.��Xv8�4 ��7F^?��3���Gg��������E�򭯸Ga@�  �当SU����-δ���m>�/2&����I~��� ��T �k�uD����[�+��!\�R~O��6�/M��������Nf�L���9"�������*�9~#��(ʩf�UA�{�9�I��i �S��z�9� ~��%WP���fas�I�Ѳ0nQia�Z7YM��K�'m�Þ��
�֕l`��O��z:�/���B	��AG���՟6�l�ڍ�r��r�@�^�&s�2=��0�d��mp�&v9����`ږB����c�S�W��PfM3N#�� xiN,=H�2�5��`��;�K��ZV��qulF��_d�)-�Zc4}	q�I<%}�n�-`���Xi0p����.4h�4�usG�3Ʒ� ��x9���a}g�(�Ir5�m71�Ү�0��W2��߮Xػ]�Ge%,�
�rfO��ԘtM"����Z�F��M�6�K���{]=�lH7��Hjx�q�nq���O��[a�t6&��B���tT��e���ߛ���}���9��-_�� �n Ͽ�pz5ןP�P�@�+���R�C{�._�����n�3�u|o+��9�ˮ�IVǎ�2��&�}t�i���ػ��<J�����N�h�T�{�����M��F,5�G!� !��6Jю<��m��ݳm~Će�F�c�0vtFD�i�J�ԗ����.�ib�fN�#_j�eƞ�]z�hί!\L����7]P=+�R�9Q#�Q#�0Fw`n5�����H�����l���ծ���/u�=>��D'*B2M4��n��H�D����,tG�9�g�l/c��\����4�Rc?F64��I�::z}�+�p�r�@pD�Gge��`�I��:��bT/�]Ǜ�0�$xDO�r#�ek����Eb����TTp:��"Qp���`e�FI��Z��fո]W��(���;��Nr�늤;�1bN���s�=(l�PgL�d�";�
z46�)����q]'�~k�/@�d� 0�e������a(����[f����l�5��1/g��Ƒb�*^E˖$�֋��m���m�Ǌ�H�5߱�S�����4@���9��k� RQ�&Pwl����d�`�/9�ޮp��?F�A���"�Q�P�ׁcy�+�L9L�m3'X��<��/7n���]ӱ3�_���,l
屘;I�������፷ld��#k1��
��0��PѴcaQ�En��Em��V�#թ}���*�UZ�dX�"]�]�쾽�r+5�����Tt��I�Y����X�A�-�/��	�M˕!.�c���v#�����1�4p�F��K*U���)���rƒX�Y1�&��I�ݒ��x!���Et�{��%n�4��9����C0�I�G�f#Q��E͇@G�2�/ZIg�/���1�K⥴�6� ��_�+��A'%n���,{�~V�mm��G:{� �v �x�d�-	3��c��mt8�=o��Nۘ&b�X����6�����-�{��<j��.%�~>M��v�9-�LDE�!Ę���]F����C�!vMX�%�N�&�K����$��T� �\�H��taag������)��F=*�6"�<������lr
�}:?;ʛ4Rnc�X�ƱP�0��y3�%k~{�O�O��$n�7�Z���X�aQ�)6h�i��s����ۦɘ��!����s��|$��y���Y§���r���x�A-��P�Kx#���co v�&k���L��+`I�(n!Ӹ���͠��W�Α|�f�Nb =\�L������_n������7�Tu���:���ZW�A
�sh�� ED�!�w�iW��`)��r\U�3��7 *���L\.M��h�n¶��y�Aݱ��i��A�Jvg�GH>�M��S���K�E��ڐ����&�;�X��~��v�Q7�#0����p�e�@���0L��9�#�rW�̧���n�k���-�%�����l�!N��H�ڟ�̔���l� ��_�,�e�?x&���%�p���v��H��������]_+��u���cxP�����  v�O}���^6���\�g�8���M�1�AQ�L="VS0΅͎�t�HG��pz=�r����o��CqE�a���۸�?����qwrj�6��]�5��'�!ᤇ�-C<�*WGO�|��E���A�qOXp�H����=O��&�[��*��X�� KL��ϒ��4���u�VAq8q�� A�� 	��A�Cp��6�	N�wwww0@p���/[�Wu�w��y����JU��zR_���n-���a9��7:j��,K�:f@U�X��]{��{��ܭQ���
����y�(䮖ޱ�-i��O�7]���塰1��[J��\\�`l��O�i�P��A.����ܒ����AM炞���*C��p���D�l�Jj�w�~�D��̙x�
�9��f9N�Iψ�	��#�,�-�nk:�!_�%s�6�J��%JZ�g[Yy�O���������]���7�>;�@~��͍^�-�!*�d�N�f�LȱӦ1��k����ŮTR���������+���B�s�5�+�d�8nڹ�����@�����?��p��Yu��vx�.���vձع)�s�]ce�B6�QX�G��WVyB"�E��b8s���\�蜇|3̎�7����䞌���%kt�O2@�>|���҃�`�����Z�;N�1^��+��v8����m�X�+e�"ׁ��B����W��c:��s��~�7�'=QӼ3NU��C�X>�!}����m�O��`�M�B%������N;��Q�cOw�M ��ׯ�$�E1����P햞M�j���5����8]�Uy�CX���|�9�� 2�����F}����m3��7}�E
�
~
�.�} G0ʇ,��D�C�?kE*��A��U<��PZ��w��XCR�[_�oW�+�<D������fv����z���6�����H^�ё��U�i�!�e��;��f�g��q�޷�K��~>|�a���DT�K�s���݆L2�+���~��47����͔Ckx�Ge%����l�>�6��2���g3�_��L�ς�o!
��{���8�/�њ�0��c�ݎ�`��c/���%�柙�8�J��Zp�or�Q��x̹	=�bd��cm�g��!��	�C�7iR�W2��l�M=O��6
�?�*����J�Z��#�L�������>��#�����O
�6�C��F�Հ�s8rm"��
wsj�fڴ�)���oOZ��S��j�6����[7�ܨ�]&�7!T��7N�I�b�qw9������c?!َ�y�E�K�$뫻�D�g�������b�����f�Nm_�r�0����i�~�h-������ʏ����u�疛2۶S��rX�2��m95�j�K�
cK����=��h�eʛ�)���ˢ��wp:9���d����en�� 3m���Ճ��랯 LV��L�ިr�q'�Ƈ�R�$���/Cڔ��-����߼����(����/�y�zԇֺ��ۏ�ˣ�J?��@�H���3q�v�Bc��)��Oʹ�=-7=�ǫޱ��$�V�KT'%_ʞ#��T��,�%�z$S�Z����y8��}���]U͑1F#�<G�w���[�!Kx���^l�Q\���L���W@c] �!������@�#`bF��!��YeF�-���<��:��`�mm�n�3���]4[��Ǵ�� �	-T�� E��,ߣ4�AC3%4����s����w���-�}�!�!4�os�,i�4�W�'���<m}��S�-��ʦ�5{b���v��_N��4�#�FGͅ�w��p`L�M�e�[�a�ڽ�4���;��*���[{��z�ж���k	���j5l'}U�5,��|@��������`[���P��1��n���UZ�8��7$*/���[��y_�bC��0L`n�N;�|8.gb�X+;�n����s�Fwi�8�����`����5VE�I�?@ܹDk�вh�ޤ+�`O?w^���n=B�b���w>�`4�5�����V
#��p��1`�qͻ�и�o3�i�,:dݥo{���\�4_���k�:�+�o�\0��	{�	0���K[��~�v4���������1�����6.ܣܻ��G9�iG�_�m���+�T������܅A_'&���m���m���T^k9���t�j���єC��9c���Ƹ���B��cp��"!�`��}�H$���}D��˫��%��G{������b�b'�J�
�چ�C�])�O+��n�� ��u���`�X��Q�1�VdnNR��AC�/mm�W=ܞ,�4���)5ĉF�I��i/���
0 �4��6��Hs���ώ��fN���s.,��<N��md�i�ƹ��(��k�mȟo5�I�M2M*U��ll����"*�D�]0#����IXNU)���q�>����?��t�%���-�IR��)�퐑=�O̶f�J���HJ������$X?;/6�r��
(�웾ڲ�i:m�Q*0�c�({��(�{���շk�0`��B{m��`(_��M��c�Ob�x�Z�
4�GB���w�e/�ԟ^�fW�ڈF�v�D81]��[�p�}t���jt���6E5oR�K�>�Έ�4�}�(ыP��8�Uԡ g���%�� (5mc���l]>��l�Pf?�U�R(���K�CB��nNF��d�K�h�D����J��gꦟ��U����0g�i�Ge�A$���̰�A�Z�c����z�+^#�I����g�eaE�^T�z|9	tS�����u�S|��s��-�z'�WkD���2�n
t^w�/�׿ES��W�=�,�-�+�v}�U�N.o2�`tSPm���8�[�fM4|� k��׫�e�B���\Kn�0�X����w�SYQQY/���=1}:����(�|͘i?�f�|Xgx(��<�&Bv�f�䙴k�h��s2�̵c����y$y���'įΓ�TP�"�Y��v���q��k0R�Gjv�9�"B�"'W�K��)�и�L�W�����^"�����D��T�,�4Am5�;k��'}2|#��K�s��R����9�&b��}�4>!��n�L⹵sq�}�Ye9�.��O��C}n�7�@M��U�>m+Q��2wY��4aS&�!�:n
v�>'�N�M�vch��S�I��S3��u^�E�U?N&(pzN*	�;��3W:�_y4��Oݕ�8þԡ^���|�����
�b3���o��4D\���g��N���O�~2H�ܑr��D��a�����v�|�@,k1kAM9��h=�Ƨ���z���6�ފ^��̹f��$E}ֺ�mf��Ƞ��.}M�,�u��.�+����Ǜ����q�G���'��8�L�� ��%�'��fv��d�+��!�:���,�L,鿩�����^�<?7�����Z�R� +�����d���{�ϖ
u)��ю�4M>��~O��UJ0��$Zɵ�P7��wWv&�� �[��1�}E�;s}�xL^l#�3�+��Bl�o�b�P�Țh�K)Zo}�g�T�������%w�k^��:�<*���؀'������:)s� u��H\A�-%����dC��3�J�86�KDb9tT�.s�`�/,։�h��w����4	�]k�y��.����֚���o+�؜��\��k��n���V���Ӭ_+#���W��,'ߑ`.��^����U(�챂D�1�qy���K�e�D��#��B�,'I��W}(�,�,f�<=�/�0����|��;M��$����]��([4fڈ��ӟ��o�gG�ʦ��k
��7��5�,Z��&�(��3��Jh��Ժ�JP���MR���H88{��K�-]@���;`����o#�w� Z����X��p�	�ל�t[8l�>����9��a����d�{{���c���G��	[h{�Y��'6 .�jPL�p�����~N~!�/H" ҵ�5�m���l��P�̅����#��B�l�t����a����7���܇-2(F�;%{:%eKy�h�z$(�g?�t6O|4Ώ)ʖk�IF[OD�F�y�a�.�*�+�3�*w��Zw�[8_/I�DGF�d#A�eD`Z���Va����;Eǝ���V)���\�+m%+���8�U(.qx� �K�d�EOI������R`!�բ��Tq<H�0L-ԗ�d�c�<��+@ƒ19����9�V�>��z�ܧ���"�l��Ah"���(.f!�H��� ����%�=������*CJN��gv�Z:F7~v%d�����}��~~m�1�Ʊ�)�R�S"A���4)�O�/�q4��g�w�cӲ�U�bŊ��Ⱥu|����4E�b���R$AdKÓ��]�-j+����;���u���4,H�X~A�3]��)���ۯ|��X�y+ �^jք��L<�#�i��M���$1RX_&�_�����P,-����Q���|��w�F��'�+�K+�#D�Yk9i��d�,�'囂����'�9���ߕ����^L��/���.h�g�W�0��+��0�llNT-4����}��1��X�4L̽�/Fe��?]���jz�L~C�Dӏ����L��e��<9���f�:���/�W�I��`%�j�9C��3��.u]~x��/B}P�9h�#�K)R�<ɬ6����g��N�W^��W�U��5ҩ��a ���,���Lf'XI��]�"*�÷����o���������51��;g7��9L���@����0� d�@�������8������䲮��;�
8��N�!ڢ��M��#�rM�_g>-i�a��Q���M��W�q.���D{���E�5w|{�����#ѷ�S��ƕќ�2���F{�K�-{�4���R��� ��M�+�	������ۅL`HJwd���W�&Ns�0��֊̨��6>2�����}X}F�x���`�5�s�Ǝ�"s����߱��CЪI�̌Ɛ'��a��'~}C؎"o[ډ5�bd�=�c$Z��]�˂x9.�~Op�flt�>g�b��n"���K�>1>��!Y�N��^���T�B/��ߑu\b��0V
'��\�J.g����u'�#"���/�h3*�D�֮'HݶnagɷO��v��~��K���J�\q�:V�5Do7ޟGRU����&�t�x�y�)]�7C��[���b��;��Pu�U�>�cy=�X48��n�Nߜ�s���.����_�'?�F�	'���t�Q�_V����A���:�?�*dOmV�n�T$ f�K�$it!����T�(v>pg�h3��wg��� �w��h��1Ⱥ+�i���CĈ�1r�@�Z���lp�B�ͮ�C/�Q&���;9D���%��?%����O��ߕhb��@��eiA�AN���)��B���5���gu��%�������%%�!@#I��J�t_�(���~u�� F�jb��:M�l������G)�%�TEZ����,��\�hts�ڎ�
�z	]�d"�^��rB�u�q��w[�1�*��.y��n ��:.^!���g��b�L#Y��֓����ã��5�$*��_У��������zx���\���>O=��!d0[pkdХLG��_��}�2��$�q�c��;��z �����ᨵ�㦮#<w�L���`��曩%������FsZйrq��T[m��8�m5�2aa0N������8�/�a���)��m�CY�U�\~�׶�ӑVv�������D_���s��ƪ�72�o���P&	��7_��]��*����n��f���E<��,k'���v�{����Q�CJ�D�.-w��
�ۖ�nm�w*����X&_����\�%"zjF-�`O�@�݈�!��k�s�]��gLu�Y�,��6Rlo�l3���%�����䍝и@Ffq��āSύq�>a����P5��<#l�Y��Ç��:�ɿ��o8�� B��lxp+�T�M]>Az�Q2mG�3仹���U%���4���X�[ڂ0�c�����Sp��G�����_��
�z�zn0�K�2`����B7@�;d�du�0d�� ��xqò��Tܒ5&JXa.K�mH�'G���齐�����~o��)��E;~h�ę/~gM������P_�
[?a+�|Q��������ިE[�c��m��N��S�d�
 ��C���%+�)Y
e�v�m�ɑ�w�T 8f���_�Z�bϳ��,ߺ_���Һ��U�҆;
�eFL�6M��?_&w{�A�CR����� ʉ3":��x
��L��2i�6Y:�����m��ޠ w����n�pIq�^��\�n>��׷�m-�c�llTln}4�����4�K� �p�Fu��)f�Dh��)�\�KI�8@��a�QR�e(b{;��ߒ7����$|*��jXBN��&F����I��2�z!�ϟ����J>���l>U��k��gAX��D�����I��-lR[ʾc���IX���7�L�^��7�/�U�5��.0�nS���[rMI�Q���Y�1��������ii�}��3e����u��
�2�,�di|&�n�8���FzO����Ȧ6��j�).�Ϊ�A�(W���}���|����xF��h�.�u�%��b)����C6��!�u�����U�����(�Vow	^�i�G�&E��z���{A`��W0���s��V�9�Ȅ�۾U7~�O>E9����ȌR,� ����΀eB�ɑQ%�%���m��yp���\�c�:�K:��
�Rp�I��L�"<*=Ҿ�F��mM��w&�����;glc��)�/�m��r�z0֭W�-9���Ӗ�)]�bb��-�NaUn}�J`�A��+}���bL�ߡ�I�ˍ/阓��q��7Ըσ�����1e5�3��9gkh�>G�
o5��Q��ω!�I��g��)��������ri�6��n���Q}�|��	��-�Ng���|�a�t��4�ȝ��������K���¯�Ԑ���w��;s�nZ�OU-Ћ��Ѳu�����RZ���\��<�h�=�@�t׀��-���,c����A���"Zp�w�Rf���8PoW"#�,9ޡZ�`���tO�72<��6&Jc������o��E|��5�����KA��@Z�ł�g���qK�e��Il�ݞ�u�cN,�~*lE����0̵�'�����U^���?�G �l���k�gj�Z{�GV��3�A+2�=7�,ߩh#��7|W�zÀ��JH�x�m�,��w�i�o��~7%�sK,t#�L{�MEg!|C5	�`%<�|rI�5����i��E�6,�_;3f��'�	����b%]�७������sz&+�S� �g`8��]z:#��uNE{*���"Da�k����c��򧛑� �(8�Q���i�F�UU@�7�u#�����,�Q;u�B�E ���7Dp�����=��t�p����O��6H��1�c���.�^�����!>����	{�ח3�����OIY<RbG���<�R\P��&���A|ŭI�����_�&]ޒ���j�W�r-�wѧǑ=��0ơ��0��U��+���z��k���/�\��U�)eļ����e�
uP(��7�-�!!�Ve�<���˨xm��P�C}�����ʝ�@���)3|.�iP�v"�NGPR�H���7��d�'k��
ٱ�u`��`������L��ƌ�;N��r��<�{>����>�
J�H�O�kq��i�9���A�J)�AFm��1 I�/1n�]��i�~�9�qr�1X��>9���6!��ȝ/��Rʗd,�m���P��$��w�[�O�~B��x r^J��B��\2q�ZX�B��;1l��O�G���i��)��P�T,����'i����~�}s2�p��%���heHC>od#H�|�&�Rp���Ȧ�~U�L*`z,�Qn��)FyΞ�q����9�3��ԁ��Gub�$�p�cQ���s9�q���,yϢޤV�2��d�mP5^�p�Y���L�
] �����Ɖ(z�_!!�&��^(>�V/1���\������MELwE��l����G(�JA��z����\������/��7	������6��$���?d�b���r^H@����;��Uz��L��P?�G�'B�6�??y�����0�y�-�Ꮵ|�tL+4�k]ƍ�?S��޹��� k��c�I��K%Y9[�/�%P��n���ſ�<�}�76�җ>�NPd�T�/�sld���T�ẴvFV���)y���a8�\�ϿP%�,:l��]���	3���[����!��ce�_)pxs�Vc�e^��K�w��p�U������®��?ʹv�`.b����MX���;�� \L�ێ,i��_忓�s{�j���_�Ô|NM�!D4J�+����z�7{3-៩z�l����y��H�jH�1x)Ͳ����̆�xa���N�ef[�P_��go�!#ղ� �Ok2S�(��<�D��0��H����휭]G��II��)����U[��?�:9�ڗ���������ۊ�G:�E�de>�B���Aչ
BS	4�Ұ��-/']�_��[*���K���_:���q-�t���Gz�ņI��jl-��	����[�wx�bO??��1�q����Az�S��o�q��p����b�5��-I�n����D��W�;�y"�y<֮~1��f2[pޔ����x@��	���w�m�'�!�[Z�b/���b���n'4r$���h���e�WG敜����y1g��#����h6�EL$p�Q�bڄ��@N�蟛�e˷! �M��ܵ��ܵF~�(��]@ �oD�G��=�M��&Wa n\�k�d�/���\��L��DK�z�E`�2����r��	t�M�%Xr�킞���UGp4l(v>	K/����*�it��v�z��fu��;4�SV&7��6�<E�P��w���%�%:�ܧՍ\��@��-ڰ��zPT�g����cr�g�`����=�=�	~��E`������P���8S�&�k��>MA\D�6�>��4'9j�,Թ:gJI�*"I�����d�������-8� ��ѓ�1�Py������e�@�D��q��jL���Gq��J��>�u����Z9O�{�i�p��b��_� �8z?��x���0��P�j��2���Dڧ�j�s��� �5{r^+}��jM9���3E&��%��7z~XL;���.���z�^΃�}&���ey�?ئ�1�T0s��q�K�L�?0�]Y�a���?��������/�}���Pr�A"9+}�jC�oꛝgp���� ��`��n��	�Լ2�:����}�;+��s��������@N���m8�|b�w��O�b������ӗ��-��G�� d,(H��>��۠�s�����F���3ts2� �0�ܠ���-�U�O���XO�s~9$E�����Bw(��X�h)}_x����녓�&g��26s¸�T�n��4/<:fb8#����4V��l) E��%P ���"����O�5�%����o|�G��:�a��!;���%c?�����结G|H�F��W~���ey.}B��b�X��Y�@�b(�s��¶Z�%�M�٩W���4����P��Ri_tgl�����I��[��\������d0��MZi1R+������fi����<Y<�=i!R4|D��m�'��� �T�3\�٨('G�ܤLc��-�?DLϑ{ϣ�<��^Vf|� �bQ"¹G�ũ�s��f[aq}X�Ŏ��,��R 6�%�K�V�ఠ ͻ�LL���B�w��mQ�����B�j?ȼK(xN��b�k5d��'>I4���d�Wq�W��wV�Y��3�:�KD�0H��*Paw i�C��Q8&���>,sX'+�%P�~2��JZ�F��=0F�Kʁ�Σr����s�U�]�+rTqӼ^�M�TԲ�I��T��5=21O�o���Č�{�M<���DS�hq�Ƒ�������<J�����?�M���9òeۉ!w���N^sW8q|�ɂ�;�"w!�5��\��eW��e�Q6��S���Q�Ta̘�H�L}������6$���qǻ+���X�*3�Ckyܙ(h�����1���B��r���/��Z �!����c�ּ>�n�u�<�v��<O�c����I}�i>�;��l>�d�!���dF)��O2�k�^��֞кH[��7J�~�!䷷G\�ċ�N:�^���S���fMÞc���o�Y]�T�m��Z����TÑ�Є���զv�Σ�c�Er�N��뷘���fr�TS��D�+�7/G��Ѩ�]ؘ����j4��~�t��V���Qv]�Z$O4ngR���)�ŕ���Bf���.���T/���+`&
dT� �����v�p2���L�����k���]��#��Om���[�t��-����B6⥹b����$Q$]�����8Ke5�V����yޡ����Bu����+�@��ґ�6��hd��+��.�NNyw!h�<�;]�e��V.�k?�ծvp9s�?
z'f�R
�>A�drM���0��$���Y�Ѩ�D⏦h�KԢ�/8�Ʋ�@�b��;yq&�u��ҡ���+ ۪>�$	��w��,o5��<z�Ձ�^VB�}I�=��Čy�s�@3��괐�ːZ~�,_cd%��i����,e�=xt��N�K����T5�sԻ�-�]4��JHB ?�E��r���rPM���[��n���{SaӤ�)T�o���rl��t,����l��$$3��=�q�j�������jO,�������Um&���ޝ5���V�{	t`ХJ�y	$�0a@�>�������H��(�]+6Nq�,W�'���q���Rا� ^�{P5J(]݅���V��� ]���jw�}��$�d�.���]��F/F�&-B7V*d.�iP�k~��|���r�:Rۧ>~�����ԍ֫��C�=��/՞��	,o�&�]����1���� t-<t��"�#��D�b�a�������oY�[S����/o�7��MD[V�^,ّ8/m5����E����ܥm��ۖɹ�A�B�oN^K��O��P\�z�c=��Af�Tk�~R�5�"Av���;U�O%�\M�`?�	��R�Z��"�L������u�b�n[�f�w�����fG�M��(?x&�9S����p��V��KH��kN.�Q���k��qQY�����ψP4��$q�ġ�l��h���z:X��2�8d̂`�L�O.�wkcIZ>����Wm��I�(t�^�M]q���t�Qc~x���լc���w��d�'͐�5W�%��7N>k����l�����q#ǌ��^Mn����=��HYIR�(/��$����g�Kv-�����(����Z�uAЮ����t�`rZ��z��APr��;�|����%�� �<G��=��Ì���G%tM��?n���Ao�b;�c�)�-��������/�m���s��;�2��P(�{�
0��F�� \�2fF`KV��n0w%��� Z���(��@��xI��#9�k0|��+`V�4�VYqN:5̖@?G�XS X�J��=H7	t+nF+���^�(t��x��࿉u
t�t1b.�>5���/0��ي�;�����ej**�a����7a8�x��m��V���h��l<Vĝ�����|��0�ݽB�y(#8@k��;�"\���$ ���h2�B�i�B����|g?������i�ić��ns���������	w��K�g���WU��t�64��S�]y��쟮�
��f�����=]"#��d~�+�e՛���	2�wG/������:�vĀ)�o��33؎*��V����������C�$A��B�<�h��*=|IJ��2�ޫ�w�����v���'��'G��׬6�-���Eh`W�.��Ü?�}�.E�|Ç�����>��B��&��9D&@�0}�Af��B�����|��1��! pg<J�֘�U6%e�+F�v�7���ݹ~	�i��4�AߍK{�c�ȭߩ�B��5�O�]���1a���k�-w a����_���W@`'��Y�~�}���?�u�C�q>ǆ�(��L�J�
,��O9�D�2��>l�D�:?'>}8�\гlP�3辸f��=�h����|����Pe�IM'�o��Tx�l��𡏨R�S�L���ݵn�M;N�M��?�o:�tyX<�� �+�ܝޏ��:Ďe�f��lw�T�6��4J��BA�fW�w���3{�Ȋ�U�J�I�|s�����ߴ$����g̷�ns�x4ӑ������b9�)�^�Z°|���"�|�eb��F^)�Y�d4r=���9�	����p7y�`s>��SͲ:KK��������x��!�
�g�3@w��v+���v��8��*>�s��X)�w�^Ivo�a}�Y��-9��I����+���P���-��OjB��BA}ѻ%���X�+�\��HA����O�B�%Z�Z0n����ǴQ�xoȖ7�d����{j~��BIlYܝy�T��$`B������W�\�ӈ����:�u����M��H��F�u��~\�;�ԑ�;W�4+��U�xO/1�OrPuS3���S�wu������������)W�+1�P�_Gvp�Z�)���n�.n+Cq��S+��՗��4�!:�k:;wwս����'.�6ʌ��(Y��@�0��d�pH�58�����қ`�~�ڋ$ˌ��)������F]���XU9e��y����^܍���]����#Ԡ�QI(Sɰ��(C>��4�ԉ�4*�̬i�.�o�z��V�J^��IU��MG^��E��)����^��Ib���-X����������)�<�ľ��
z�:���
���ndҋ�W!ب��6����s�vGpʩ�l%�:�'0\��c����1�y�m�c3^>Q�g-+k�y����8�!x"��M��yeHW%Ӗ�v�L��o�xQ�a7���R�剬m;�e^,%�o~+�,)��ŭ�㔭��K��(�n��~�`�ʓ��eܤ�v�-��%[�O3�6Ӈ���L��Z�rV� Q�J��έ�q�54�����Hy���{y��CL�{Q���z!e�M�ޟ��Gq��ݣ�,��Q-�w�h^8vQ.��M������p���v;�.RivJ�]��o"2���8�6��f��z?��[s��NexK��X�V?ɒ�t�e��(����,ٽ�o���&�x���M	���p��85M�0��S	�I�Kx��+��;���() 4t�h��&l�������jp}9w�A沸�$g�ڹ95�Qq�N�W ����ʹ�����G�&*S��o��/7���6I�H��M�]o��
�AT��OLJ�6JF�3ұ�IN"�:8c5�����精t��TQ��9���*�Vɧ����E]�� PK   �X�Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   z�X���b�  �  /   images/84b07818-b924-472b-989c-78bd96a030b6.jpg�WwX�Y��(B�* �B���ܕ&]�D�C,����" E�@@�RE�ʮ��4A� ��|��������{��w��ϼ�̙3�w�3�cM�&�& ����~`(
��_0���	g��A.n$���@"����
"��G�E������������� ���9��89I $���j���=`��H	b���  }'���(�BN�y0��f�^�`�P$�免����m���ǜ�3�m�6�2�W�����;&�p\M]CSK[��,��������������5��uO��w��CBc~�����F���������
�=}V\U]C������u{GgWwϛ���Q����6=�ivn~a��um���&ck@@�I���d��� �������P�Qe>#k�����*Q�gRW�q�TmV��8,�F���C���(���߀���5pC@l�A� �~E���xN���R���I���P:>"��J{CVϓš����>�1j|*_n%��WN��>AOn��^�۱	�g"Wb)V�kN�J�\/J%�I��C��,����טw}�X��(�y��p4��&�G<X ��ᓆ���~�)8x�kySϝ��l�Hd;|�����ķ���ݮ܍|� ^����2�Gb�̱ Q�)�gX���v7�fή�����Sr(:���y���i��"�����b���6/y(@���X2%��
&�[�9,���� �`�.*���E��ҹw�{�������n����r/n�C��:ֺ�$�W��?ȍ��kP��'d�`���[z�Ioƀ���$�.)xN��`�[��B\z/L=�K��oJ�� ���1M��_�^BSė���һ��,�Ҷf��ߠ�\S����t�>�ZN��F-D_�"���Q�|Oz45��u��wZ���Zo�x��Lڍ�ω��0��# �u`���g��z=Z�_C��v;آ�(��Zq�����m`2����Wĥ�F���(:*U��^��2+��f�k�|�(��q�0n9��_e�KW~|,�m�O�Y;�W*��?�G�6B�c���5�y�� �0Љ���&�\t���fj�~�'G�Q8�&�dhZ�yj��F?��g#�up���w�F����.������zw���[hƬ���]\6���vx�SD/�9�6:��-4OIHO��r	a��
�v��bӂ��`F5���ٔ��Wo��4o�DV���79�v�|���9 A��O��ޟ
���S���J�7�W�G�nl�����!��2�o�
��d}���
q���=/+@~���y�������bl ����C ��,�S�D^�H��ѓ����j.[�p���=b40gJUxll6l��kdV#�#J�;��vG�#�����M<U��j�<�`�|�*~�<��?�Vv��X oMRģ�&Uh�緇4z������������tW�|{�x���;��r��r�ܒ�Bb�0��˒�p���X��}c�XCO8t�W�[��!ŒFɹZ�"9Ų�	���9�t]oI$��=�x��Y�G�^7����J��Yū� �AJ���&|;�c�O�����ɷ��j9���o���?�uDr� H"��&��g�?�jt5���`(,P`#��]We��?�Ut�J�Td�?sjhٍtd˽Lo��閵"S�4�5�[EP���%yP�M���&�5���, �����a�g�	l��g׾�9��v�^�ͪY������upI���;?��_� �*0O)�q�P�_v�a1۱�ѓ.�ƪhgyak�P��ds..1�C�V=��6Ti����6�o�A��q�)��7�?W.x8(~�kM_9�sw��=�k%2c��1�}o����s�xI���4�"��dz�ۥ�$o/*<��N�����S�2����3�\�D|β��#�?���M�=H>ed�$�� ��Uue��������G�����¯e>����#1
����ȩ�о�f��;��I=�uN�w�2̶Rv��ɹ�	�"J��MhP�/wd�Xec�6��\���_�n�����O����V��3�Ŋ���ZhmڙB�����>�j3��]B�4#�$z/�)cY@��w��o��E�c�k�ҷ�^�h�4K��1bu;R��,7�r�lF�!Z(X�z��2-�(���=�s���y�=>�HMs$6)} ���~�-�x��B3�j���4��1���q�k[�f|��c����W�tTr��ծ���L!��:�m�W��ǹ��nL��s�-��oqv�؅�~�Ƞ$�L?�g�H�L\"wJ�NgS�¥�UE��u��i�a�ҫi���<zt�����r*���\�R�;l��?6f��6Ca���;h��孥Ң�Q�m��ܞ�?!ο�X�, a��q/���xo�o���=�g��k;�JI�_�[�u���sh���'ϣz���C�+����Ή��_h�=�gfHd�k�<Pl�Ѯ��gp�k}]�{��B��m�w?��a�X�S��b�}���$�F�G����� ��+���J�3�:��nϦ�%��p���+��R��Є�*
~`���G������.�̯c�݁R�
���Ը���T���x���C����>nD1�
�m�>^�,]��R��A��v���浱�E�4]��*ءM���@���{�שk�j��t��hx�~�T����y\O���N/���h� ���r�M����s�/׍��wϟΟG��	=r�R���U�if��rߋ����q����!L<Y��.�u�#�-�M�4s����E�[Gtgh�#����1�uȃ�	��?rtЙ�, f��=��"q�������>Ʈ~BN�bc-�G��Z��6��e���T�DV;(��ۈ��^���u��8�*�حde9;*���>�qqv���h(�7�b9�Z�����ծE���
��(���K�9�}A��1�kK�#��v|�$�"�-��Z���;@�ʬJ}���4��>?��,|��O��
�?Oed�Ck02�C]�>���G��K8�R��P	�%�E�tf��@ja���j{���e�`�Y9+��A��$�C�~���p���x�[��[�,�.�Z�� gp��������-(\q�D��f	��r)"���;z^E�ϕ2//���+YM�%�{=S���>���5-f�/���R߄��}�p��%!��TY���J��B�O�1�;l�P[j�b[jv^4�����Ie	Z��M݈ ]3��ݿ�1Gs9,E{�I��E��L"h��߲�ZRcs3����L|��f4J.�O}g����l�����}�6˜c� c ���Vˋ��ϭ���TU��S�Q��c��7�崓I��[cF����y ��\�M�C;��-�̚��xSS�P�ܕx����&%��%Ma<��P>,%�@?�4W?�|i�N�ǀb6���(������0  �����C����|>hB�K�˺�ӈ��5�����D����ᗸ��''�ݍ>����F���t���q��r��c�Л5�*��0I�m:�_��y�<���˘#O�,�K�U�m���z�{�)9�|oE-f�7�ݵ���Ŀ��́�N˔Gl���^���U�Ց9���݊7X�(������f�<�����Ij3Ջ���Y�;B5(��u1��B�N���w��ó��z;#����'uW��T_�$=T]�a��h�{�R�[@���-M���ᓚ��uu��{���X����t0ɚ�K}�\��As�f�V"�R'-��K�u�5��C�	�ڶ��]%����+��:�"��K���nP,`�Q�}�G�ص]�`���%��`��!]9��X ��_hY��!n�e'0����<'��駘<�M�� ,Er�*�����:ٱa>T�L�wB|xM�F&�ܮ� ᩬp�����;�|2�Ա��4�q�삿EsHƿӪ����9�H1⑬�8�=�Y��PK   �X�X�ԴØ+ �{ /   images/85110ed8-4773-4cfe-99cf-d6f3d0ce91f3.png�Zy<����~�H�J(�3s$�ز�]ֲ�]�Bci!"ٍ,QȾ�e�nB�آ��32���{m��������}�]�庯���}��i��PQQT���KE�g��j��{�3;�.��vWP������:8�v�pٝ���5�ߎZ}=��Q�Kz.�Ыn6TP(��|��ꪫ���.�(}������9}���AXl��ͱ%?�A�sN�w\seoe�Zt�����BaǏ�߼�<�P�U��Q���N�����ۣC��>o�~�P�?����ʽ����"ۃ�۴\�z�)ۣ:N��n�e�]Rj̏�"��!�Yh����v��{OJrR���o��={gfY!���J������m�6;���Uy:�
Yu�֗z7��>���.�@�*խ��N�vqj����zw��u_�9q���KK�4�BK���d_�3U��@\ڣZ���˰6�iKwZdoү�2t/���T{�C����,�6�ڤ�P��څ0sl�ʒ��[��'��q���Om§?�������i�����zxi0��M�]��2)�|IBtϯ���!����}��qL�6#%+�О���@h�]Ӽ���x��O���Q��O?ݗ{�|�k�o��u�L�!�/7��������T�}�y�DI�/��
#����?/���x3�~�>� ��v��?n?�s,���}(�Q���ä���k�n]����= l�D�֑.�d�!�Je��V�_^��k8J� �y�{+l��ɭ����A�[O^�0�b��-1��I��;/�u�)5�{��\PEy�����߹q�P��		v���O����өö��kZ�}��~Y
���� |��|T�=��H�@�m�mT��-���l��
`#�9Gh�/m��a� �����T��L�)�ׯ#�^W�u����ځ��<Fg���7}�`��_aد*#���SH������%���ff7�xT�ܥ�;l����0���պ��W�1 N=ܾ��n#&9|gϟ���e�4���{XD�v��
��}=US;�'6�k�^y��0��=�� �N����.��\Y�?��E����٩IC}�j34?\�o�|��fa$ʟ��ױf�}hU�8l�At�n���[Em�V�L�Ρ��~�� �뀰�|�w~����u�����%�u�&:�E�R����M�e�o�Т��)� �F"��_��/pc!hy8���C�@�gԉM;?�k�){Hp��q�=IC-�U���b+@����<J���Oƛ!yX�o(S/�p���ڤ7�Ֆs
���N -�x�̔x޺���ko��Q�=�p[Wn�������HTF^(/D�E�I�@_%lb�E��P
��ݬ�+J��f���Fǐ�g��v��$�8�̎ߨ�m!�=�If]4@U���	IJ�f񰆭��_n�k���T{���mh��ڈ�u�FI�	���A�H���G6�Q�f�z0��
 ��_k���`�T?����_���=Bk}b��~-����	γz3Hx �������ڵ���}��'��N���J�W��ļ.���`�C�ԯ���)�hK�h�_ �!���Es�I��aJJ*����������������6D��\��:&@�����/J�)�iZU�ƫgfeȊthJ��Lz[��i8e�[��#���<R��(��V�@6���>��"y3���2�ou�B:�_$|^ˌ�ͧ�OA�	�NY�l��n��@��ԧ��*w�Ξō�+YX����������ƪB�_[v)]HX8yc-�[=#:�ecvXRecv����ǆ���$�����5�l�}��@�t��յ��E���7{���n�݈�,Ne����d��b<�����,��k�+a�!�Y �I�,�����9-�m���Y��~<��e�
Nz�f'n�ŧ�c� �g*ue��\�6}��2R{��A��[_?����f�o��m��ph"͑�f��r(ڬJ��ȉ�#2��Q�8�ܘ�7p�E]�Ѩ�Pf~AD5 ;���~�x� ��鯍������ۘ�7[|�e M[�)��(�,�7�?,'��t˫��t^�%�Ojmy��ɒ��z7NL����o��$�{mVhއy������-�a�X:ʵ2��ٓ�=��ڵ�qv~��<�S���j[����t�1
F�aZ����w*ߒ -��:xV{$��x��{j^���cD:�\J�Q������4n�'��-�c�e>6Q�>�n�%:�֠�Oe C��ۢ��~��,���!��m���0^F"[:� �Pѯc�b?��J1>n��{Z��w-�0q9��o ��0%#��p<�����'vl���WƽS�7�*_�Z��mf�g�c��ᱞ�b�����d��`�b�/�"Ez�k\Y ��U��	����b����LM"�:�P~�	P�Y:HC�*���LF^L�~���� ���՗kb�[*a�^�Ա� �����ݧ/�h=�one�7���~)8x��rBR�"�=CxPy�e�=�kl��m�ڠ����7�N*`�!$��>�X�m�f34-���J�Q�U��t<��{�7�bQ�o��S��$��*[��8�K��tt���$���TW�s�=XfaX�@p��� ���B���FQ]m�iȱ����z$<�,%��[�71���۞}C�p=�$K� �ζN��.�7�L�a����'�^�7��ݘ1qsg2ZH�����8��W5A6�gSVnBXpBg�)T����&���LɎگZd�a� ;�r��4J�l��/x�<O�KA�Go����%�VS���ޏ�4���������@.U�p߾�ikdP�E�4GQ/Ԡ�ZH��o ��1ص1Z���0^��7�B��T#�xNa�h�r�E����}�����͋x��J���3EB��
U��d��;D���`���	��� ��u����>���C҄:FK�D3Ϙ�����&�3G}��6���vQ�@����2�1��+nA��9��"Р�Yb����J͋<���iC]C���ə�?!lG��]6V�9=J��٬��n��w���6٦�/?M*�Ӭ.`��c�I��T�fbʗ�Y�RYq�b���?R6����D�˙ bk.�q�*�GO��i�q� uE�6�Q(K�R��[��
n�A��뭭��~.�+��7/&��Sc�+ר~}j��7������U��f�!��+a�ChJS�QE(jic���I�]O�*���l�u��e���`�_m(��%Mj�+{��\�$ l�3-�%zzcW�fm ׎!�����J�v>����L��!F��s�XUa!o�|3�_��w ��S*���e�#u�A��A�<�%�����n�]�P`,��Yig�e<ޠ@��%(�v9����\����O�hP(_��'= ���?�d&��g����m��7.�����P�ܚ@DZR
�aX��UFb�� n>�_�F$�����g�8��W�N{���&G���䋞њ-R� �`�*K����@��Q�G��F�Ώ
�Z�s�ҟ��O(���b�v���(�@��a��T{�om��e#��ÿ˗2�`�p����̄�-���Dq��Y�!޿i���y3�u�Z)��,kk����h���Z�Տ/X�����n�aX�#�����e��	a��8);҅s���<1Ǿ���os�,��^聹���\Ua�q̀��J�e����E��͋����I�I�+����А_u2v��Wu�q�u2���[���I ��R*�R��\h���>#Q���d���}'�g�k�fv�:�X��S֘$N9\t* :�
&���9�I�{(X2�G����.��)l�����
o�TW	�L�f�D7���6�"b �Fr��D7bpF�E��8�G�B��6�l��{w�2s��i�Ӌ�`�J/�����><,�os���N��JB�s��
��O�+k��y�
}��5®%;�Z�����}�l����Űq=ʘz���rH��E'�W�)�Ϫ�'�K�H40�!k�ل~�׽ a^9�d���\����Wa�Q���4�cn4$9�ODI��a���$O�>[��:$R:��j�tWd
jy���f[�����}�t�!�EBXL&�%^ca�߄�� ��-.O��';��o	2���&3�W�~p��H?��l�^������9���!�R����a� 3j??@	ɰ s��7���F�B�_Ɏ��I\�^�e�T���ё��<s���x�ԭ��^:�h�Ꮢ�U���Yt�K{����c�vQ��I�y`L r]Q����]��o�6 oQ��$`�\�����a$
z�<M�HX&3̱$�o2��u���cF�WN��->�Q�!3S�)�o��2ǝ�T@"����?f�P�,����У/+�z�&`,�O�V��0r�4���咥՞_�5�j/����_����2�^��n��!�1Ԓ��:s�ǲ,�P��������O+�l��l�NT����Q(����:�<"���4����*��ٰp���ʛ3NMٳ�]�}������`V�j�=�{{�\^�T8 ��`���/g+��� �MC�Sx�Q����t��vƁE5%�Ff��Y��<k ��b�2K"�B$,�)�ŦOҟ`�,e,\�U��X�|�:�U����~-�M#�,�g���+��D۾�Uk�>o{��Ҟ��OC���� ρȠ��AGЛ�8��ڸ�X,Пh?�V��̜S�Fީ7�2���SÚ�`���.n�#�i��B�2m�S,

����@�j�����`�͋�DΪ�/i϶���5Ʈ}�)�%y�4�i!���2I������IC@ܡ�?+_�/� 0I��vs@��%�s�g��+�G)4rX�ME!���̒]��T�}2��Q�)ed�B��GG� F@`�]I��Qͷ%���gܯ�Z���w�,'��p-�5�O	|D8�_��ʝ������b���G��� X@ -�� ��_��U�n�M��1�=m)Dg?��>[�9"QY�Y�(�[Wq��zĽc�j�n�x��nK�E\�cVG�l�>L��D�^;jKɬ��i�\ �k��-�:4?@=���kU�&'��.{:}-���a�ݛk�΁=�F���~Z��KY��٬���o8g�iSVƀ��s/`�Q�$
Gw��G�7�`Gh� s��9-��L�-���Pp���eWf'~I�^ۂ�_�vJIOx�����HcP[:2lYf0Q����ԣB���~���w��/d�QpzZy����'�"f�t-�B5~����l����≪��$������Tn���48@m����T烐p0"�K����,�ki �?���:��W*${��mz� �$1�[/�Oa�z
�+oNY;8�><.��	�%j�,�:�_T2�mh�|$�d2���7g�H�㒮@����h`��D�K7e?]*P�bý��3_a�cD��.,<�\M�K�phY��N��1��m,Ձp���JG&u0����r${Op�Uy���^�.�?�j����$
l���ѡ��E1��K�.m])K�J�v���䆙�u�iG���xI�j��ű>�Q���1�����c�mU�?��M�B���,#A�m����O�uv��J���۬}��;�� �s�1�v޹P^S=���n\���Z�k��#ͧ��A�\C�����r�����)����)t驤dh3C
V3�A�$p2����n�g``
�9deeٸ��]T����G���%�����n]� ,�)ٿ@MN����"�nm��b\��n�;��Bx��3���0b%Sh�[�I�3f�SVI�NZ�r��s�	��{]ĭ�KR��� M�g�E�ۨ�/f" �X���I�YJ���cIL�Dx���dY�Y�+^-U��C!����K<����
��,�T�K�6�~��W	d�<Z/G��Nt��ñ�e�F�t2���-�oy*���#s-ظ��;��s\1���6BB'{͕����/%�M�������v��`����c*�`����E�������	�fu��ɨPO�$�}[߯��zs�.��5��"�!��:ql}�$.-~8���,x�� ����0���j8ΐ�?��E��}*z�� ��hK�43�R��@�qt��j7��m]�Vm�a줝�l�	�>��Gح:�t�oj@�wm�:��]	��7-��1.�Ue�d'��1�ߨthߞ�,tL+�5�X<u,\E���P��5Z�U4IrNLudi��ϋ�`��J@r�;�O%�Vq�w`�g��d����{�C��l�ʚ0�ts�d *��d����V���E�V1oBr����R0Ǫ;�����!�x�@�I+�G5MЦ\��-����W�G������U�y�*e�(<�n#	�$8)W����E�"�f��v=j�lƇ@n&�wo]�˲�i�_�L~^�ߗ�S,aV�e�9��|�����U���ƾ���L'�,ծR׈��d��7���[J�X�#�2Q˷cA|��ڰ�g	�^fXG���Y��/R:)�F&�� �5��E�����f,��r�$n��|LCg�j,��l`�H\}3�vp>h6��i}�h%�Ӆ��Ȏ�*G��7����*q���������KiJ�Kg��1�9vP�j �&�͋�@~��W{\�܆a���s�=�-F���a�}ޙ���o��_�J�-}o���]^l���-a��ME��J/�q[�����jh^u�7�N	B���[,�쬻��U^D�5-G�c_�G���^r�2"Q�Ʋ�#5��/CAS��-���A�����qS���U�,Oi�wRA����O�A+�g��4�W�m�<�f���]������Q3�@� '�Xt�p��_k#!��D,3QY(�g��!�_k���P�~�Tb?t��+�Sw:d��p����"�DS�P�.�9��k�8�f�Jm;Z���g�F=s6;d_�'[qnA�Y�����a��ٯl-�~�-����G�-ǯ� D�������%��'퐨�����|!�΅
i�bN\�K��≯��:I��ݭ�| �H������c����ɴ_ɉQ`���He�c���Փ�d��C��'wI��.neB��q6\S�]�D2�z��H���> ��
�%s�ǀ�f=sq<vm���Ƈ��W#��#��9�L+�	�w%���i|�
�a�=Hܲ#��0l̵3���(
f�B�� ��ڦ��-(Ax�H��l]al]����������U�̹��gs��||�Wm �M鰃�Y �L9U��Z9)e)M �l�!�x@��ah/g-�b�^�JMK?�$a@���.��$R�E�]W��	Z�&�Xx���[� �y�a���Q芘��L�`��_'A�9F����Y ���~h��KK�+�va��:�_)$_Ӯ���;<����s (���������ʚ-u��(��%�U�5�v��o�YVu.��yxu�IN<���)}_�U��3�/�!j���uih��k[W���B
�y�i�Z$��Y��pC,:�yb��Po����Ԇ5��T���g�oWӶ`)X��BT�)oY�(@)H�S[��2]�4�|�%��X� =�6�5q�#�����*�
���-�ݎ��˟�� ��1��Kr��ދ�����|�\�)��ƢrP�,��eLD)�rWN����ך�����;��ZEyS��'Rݩ�:2����$��Ժr{02 ���&1��zc�{0�
�C5�/L�켥_�4=W8�.y��(� Nu��iU�Ն���4N!�?%,��{k&��������1�������ӧk�[E�䞢����oxNڗ�v�m�EE����!���H������a�{ʨI�/b�����~92���n�	DY^�(3�n�x�������]�ޫh��F����R8��K���H�Uo/ޚ#�ɞ���2~D����x|�KB�Mԡ���9n]R���|Klj�}���-������;c"O��ș����e΃RAp���j6s��V��9��q��m�_�_�$S��̑-czI�T��nY�M��Qrծ���|}��/�?���	L���i� hNZb��v\i:Z���.R �/aW���n��R���"/����jjjj�����D��q)�8���$����w2��5qOd�za�_Y7���Y���F8����R������n���i8�-��N@I���F��`6 [.��Ɨ9��w��4L��P꿶ܑ�z2���4?c.#�a�y�?"�CF� <�0�1xbO���R>mv���Hh�!'�O�[�y�i��cX��Z��[/��v� .ͧ��බ��%��{���n�6-�7�dv��������l�ƛa��eN��#K�����}n�qxu?[�Vգy(�q-$��z���Xv[�p�8��$�cո�*o^���Jp�Q�5|�<P~��	r+m�E�رU>��`����docs��(�Le����\�舙���]~���v�]���oIt��� ��c�[wej~ ���7p��n7��[/

x8��j|�z�KTF?*���"��O��Oh���^�~a�F?�0�V毞C8�!<�p�v�wԗ�I@�������-���T?�����F�H�]����(��6�x�����w�H�5{�Z2�.gA��N&^���S[ft
�������go��	��[��
k�k�B�,\�S�@y�}�����3��
%����pz����w�`��Y�W��|mބ�6�!��I���)N��������%h'�� / �-3qߛ�����6��� L�_nH)]��*O���o�0�(+��U8��T~,�
�`� ���7/���}��Rs)��z���#/�� ��/,8���+�]�<)���C�YYs�ta��1�3���>$���?�`��^Yb�'���ȑ�́��X��-��?i��:��q�^���r���)���4m�9	�<ls"blhl�0��-q�0�I�X��ӱ|�%I�Q�׀�X)�8Ɩ֍!��������w��r���]������s�����7���x�D�@�l�XN0<0�h�(Ƨ�e��M�.�ػo�s�2�d>��.�����B�9[�]��YfB	�����E5�'&����^0��p��;�Y�lϸ�A�tq0,db)&� 1}��g�I�J�m faHZW�V9�����"���@YZ�������(^{P�Ź�
�W-�6�t��� ���y� ����~6.[�F�-/'�X�/L�B(Q&:�	P���S���*Y������[�I�9SWrD^B����yQԅ �/��~�*#O�</7����7�O% c��fwx�0���YQ�|���<�J@%`�V�B��/F �����q;i6��Z�?���6�����w(+oh�D_�+�����ť��CsT���F����Vr+��>���"���\�b�C@k-y����/����sFF�Ve+���V2�&��< ��J;O����:���F�Dx˻�*��e1.R^��I�z�籸�ȩ��­����E?=N㢮�k	xP�hf����N�3�RR̀?/��eΈ��������x@-��N�c���ψ�);_E�N/�[*�k�f�i�1���Ə��`���v腓D�ܝ�x��4D��l�6������J �|g�*��db���.\��8��z�D�l���9w�מ��cã�%�I�����<��(Z�\u�r��(��6�0�MJ�W���ǏGY/�+	ĩyV����s@_���8uz���qK�n�d/�B�W���puV�.>�[^Ii(`�~�R�IJ?&�c1�@�|:�L�j��%�&����!yTjߕ�]Y,Uk3)$��sd�Rџ�~�yUw�O�5#�# ݤ!e�c��t�]�	R�ߎ��㬗���bW�i�`N�Y���k��7����L	���mMm����Y�I����"8R���0�c|,�3]��N �$x��G�h�v��q�L��}��j���c������{;&̭v͝�>�<7���=��S�D��Sŭ���.�o����J��=N)7\����ϝ��S�^�@�Zy�.Z�r� �P�d�ة�Ę�T��+�]����)��;B4�OǬ{�w�_\w*VH��,ޣq-�~�'O ;O1l��K;ggbk��
�E�}t��%.ò�;��������|Wep�~,�3
*���ӡ?KΜM��{��a�ʞ��׻ ;���!��t�F��]t�i�r^CY��^����3�H�u1�?0�$mڵ��5���pE;8�fJbL���b�����O �)1k�|�� w����f�G�\���?,'(1$ǻ���z�߄`��L8YY/�TM�-w�{P��Ba^m�i/:3PS�sؚS-\E���Y�鉬�Ouo�'yU������m8���Z���[���~��g��NK�)��_�E\��՗t_ԍ���a��r#e��\�����K)��B�S6#������kF�Rd��1�������N�3�V�3rn�?��J-����p����_�pr֎��]io̥#�F���b�M�}�-�6�Xӧȭ�{��#��P����p�S��L�%�Kp���s��+����X����R�l�5Y���2c||�1m�ٺ��`���4�]]_J�����B����zV>[L������/�d�m��
{ꋯWj�?���Vvл��<N��R�z��z���"�f�(�D��d�)���c}�9�e#:(.���|���S������Wˈ��h߿�z�����}��"��d��af������ �ӧ;� H���bSGG����߱��Q�%�u��3Z��6����G#�g�bgP6%��n�$��1d`.Ί4S��g;��Rg��1auj���Ne�j����ͽ�ÅSn��0,�K9��/��Wh���㣤dmm��k���fJ5����)
����������b��; 3���ceN�p�>2��m��[�ԯTb,l�����ڊ{�������=�-n�֞���{�իsV$�X�=?)6��v"�u��w��9܏ Ƈ��/W�}�{��P�ŗ9R˰��l����I�9<�c�i�Q/��u�Z�3����|��(#G���Y)��7T� �2z'���L-��o�����@�OY=��/�i8.�Ic�il���%������-bH�o���$|�6�ē"�� t_x��u0���­YO����Z�k�.��ʸ����2����'�FN��Z	4�R(�)��I2�ɋF:�ǧ�!
6m����&�މmHd���%Ƽ�1?L2�oL��L��\�Z4���{�n��h�$��F�%0Y�Pi�×�.���<�4^��ө�M���"=d���\_�����a�0�}7w��,v�`_u�F��(���Y�)�^��� �Y6xf�@2P�Msl�����~i�t�}�Wk�f,?�~����\�/�-y_�	�Y��f�GBf�-z��9M9���J��,��~<�s&��.����r��>�P{U@�D#��K�� �������}�1Whfуt�M����{���0�V�u�P��������B�3�:��0��a���9�!�>�ORY������d�-����O����-�uZvm��hx�8N��j%%l�<��8%�����հ�gB�d CAחF��45_#u�����ֹ��P2+F���ik�����߈���Yz��MF�Ǳ�~�E�D<oꕁ�u@Ϟ7*ŏ�1T�t�ݿ6P�]g	1ś�b` Ԫw��{f��@�ɘ&Y�*MsJ��	��ϗ�k�ᴍ.�H5.�i����?��v�Y땆����rj{����>v��~n�+�m{<�kR�)��e���h�({�JG����A$�s�n��y��l%L�݆�9.�|��r)��BU����@k�޽˞ӽ"���ID�du2��gX�W���8Cd\��p����s
�?T��C7,ɿ�̍�vb����#G�'�B� �ۦ�rg]?r�-��i4��zl���w�{��;�)�2���� ��k��]�E5ˢ⚒��IN�88�-ʗl�(���%nn�sh��K����)ВOж���X@dee_Z5<|�{t�ӧv������>����H臯�?���*�n6T�����������R�u/ ��m�<`�&4�xpn1�R����d,���b�� �L�6�[����w�1þ�g(o�o�<`4����ה���P�����Cj��o��e��X_m(�n<H��t;f"��jc8��\���P�y�n�����_�?6+�~I'v����U�!���_���yp>�=y	u!]�P)cdW�)J�T5��  �Ꞃ�.�^}�N/R�2@�=�+Ѷ/b�*L��6�~k���KqS��R3]�E��������pz��p�&��� ?�)������ޜG�^_�p�3i��&�0~�KJ$��U#�~s[� �D����P^Iǥc �W.��}��v�m��i�PiL)�)��;�H���$�?~rN�}JyE��4Z�E��j�"ᚂ�0r;Ю>s����a�x{׾�2��xo�<��L�#y�7S�P�~��cRD�@j...?���������L��7j��F���.q���\4��8�[4�|�S�g���@�(�~�)�����Z�n�Pۏ,�~�E�/]�F.��"REM��Qb�{t+]v��h�
��e"�e�u�p0����j9']K�I3�#A��y�oea�-���*�LxUe>���b�{T�g�������s��ii�����B�^�h��V�ПC{��ZGp~��t[�K�jiO���hR�D�Yug�0���e¡�n̭w�������3�
r|����?L�5�|�R�G�]���p{�:�{���
;� ���5:�H���ϰ,ʔ"���e+���m��Gk��c0��(�3n��V�x#�g�8���\o��P�Z����3ZdvFDN������k��X�٩��>/�ۗ�#��h@���u=�Ǭ� �ⱖ���EB�����6;;q�m܇WHS"̬����a_�%�T*����N����lc��'��w���GyS#�?��pxݬ�O@;�Wy��_�j$�9n6�o0���� ��Z�c5�c��S�J��x{%*;L��)XT;a੃�f���S�:Y؃�͜ ��wH�t����yxy�m��x�1:�[SS��4BV
:ZGM�V�[Y1tf�`3�KH�� �fOFy�>.rTne�'y���3�G�ҷtDRJ�1@Z�!�xxU�j���Ud�=��je1W��v��^�8.7:9ꠤw��K8�2f�Qﺟ�� .��{2��I�r�X_�j���Zb>˳�\���CtI��H�}�\�'8�8l��q��T���A��"��k��n�N�3 ���Z,iWKw�����x3��E��=3���.������p5��oa԰j���ZC\Q>|�V~����k%ƈG�%=~����6�T��̉kW�A@Z~�&Kİ0��N�QWؠ������h���4��֣��Y�2�Hx	�f`&�W�Σp�έZ*��=l���a��O�qk;��2fw��{��e�v�>P�{Hn\��V?l�<z
��UΟg`b���D�帔��l��_m�,ɽ�5�LL����%5q����J���a�qw��A�-f`C�|���߱�A6dğ�\�߀i���_#�1��^E��'e'��G��r��jV��)"7�y�Ɋ�髭���I��M�$L���\�)���a�dN��"�̽-�/�9i��}ծ�$i*���	��j[��s��o�b� zo�>m���ڗ�P({7��o�W�b��=�j���٧��B��d��'f�x�YA����1�v�d�H���E梖��э�6�!nN;��N#��h�,±�I�s9�JE�IF�=�(KJ�n?Ԡ�쩏u�g��׈����5�u(m���F�d���+;QM��*<z�sjjJ�81)��l��ծ���#�����]C������S�^Q���?O&qT��zO�-{ؒ�B�ҧSO�TYh������TS���G�>eZ��gS_�X��h��ɘ}3	:+ٽq�9$ψ�j�S�ɏe.�� ��2�@�,O*B��
�%C�x�V�iCK9sF���6�s���gߗ{Y���u#h��-�P�R������̖;ɲ*([[�;p�����.��t�����X�U�B���G���<��W�34�x�� y�P��҃M)��'�?���zW���q�]}N"?|F�AL�V���\�i�CQ;���x��x	�[m��+�M*�$`� ��؋��B�)N�6���)Q .C����G��
�Y_���]�;����pY@T:���-��Z�	B5��ud���ѯ�Tt��j�����B�)��hb��~CϢ�b�����ԗ�S0�W�n�!���φ�@��&���b �T1΂��ĸ�������6�+9�����{�cJ���L}bh��Ј&L�P���>jv�P���`�V�yw�ŗ�e����[:�T�mp�|u����~J����;��~�{���LU�d�Y5vz/���'N=B�A���9O��Y�R� e�5���Y*�(�ޒ��^ȼ��}[�y�q?�Q�t�kU�/":�Mv.�-@��<�ޖp��&l����� x�c��E����mx�(�/e�����\� w���-�JE�H�w�HNO3���Ԟ|1���u��Ž��n��8Z��ԥX�MY�^;i����X<P��O92���Pd�)<�{>|x2p0q��B��͈C��V�Ė��*]۵k���HTFF�С+� ���<��R�jG��N��]G��-�ʺm8ǺB�X�����n,�ͻX@V4~��+�k��i�?`�����`�ո�230vO�_�˟���ţ��Ϳl�� d�����"�d��]���nȀ9���n���/ɎT�p��� ���}�|�-�*�������o��Mi¤aI���n�r����R�����x�n�9��[�7��a�%�B��]��G.��+<rR���ʎ�p�H/�)o� ]��r������|��PO˫���SV\���|��N��1���G������*��H���*�X��=�]J{ �l��?cPz�58�8��P��* )qS�e�l}�5��f�(��3t���0�l)/��x����`�ӈ��L`F�O�qv`pߩ���"��lC s����B��w_�q���b0s;<�[89`��)��ۋ��A��q)�ct�;�T3�}א���|�n�quа3b�X�O��pR�w�nu �R�Fxkâ--E`��g1q�/��z����t�z??.�#� ym�G`�+��>�9��?s���	���AG)1�hD���L]kQ�;}�����Xr�0���]�	ǄZz���#�)sU�I݈i���8��.�J�g�;**�Ᶎ�Qy:", �%z	`�$k���RV$D�4s�W��"��=�
xQ��)�~���*�V�J�l~Xg�m"	��:�6v����$���d���)�fM�~N��WNҦūe\�w��mr2A���A�[�꜀9��F�5;S_Jj7����7�y?D�9B�)t�JV�\�j��8c*1���BߧN��2J!?݀i�;���[�B3%\�%�{j�`�*X 'Cp��=P�m�hm)�#I0?0"����Nym��s��Ō{����󢝳��@�m����l�#f����Q��Wh�Uq��W���$nniAZ<y�1zKu����l�L]�H��8����i��b�8�|���H��K��F�w����\��p<�,�I�.�-I�C�1O��맔3*){}�w���P�
2�a)�'#Q~�UI��y��؈�HM�za�'�<)���Z�\��P�$X�Đ�/U
<�em~D��EZ�;�B^�����U�/ �QBg�!W��K������9N�T��	4�����i� ��~�<��;�MA�V?0n�)��F�i��ж���
�0/�j�1��(MdSs.b߯6s�SZ����\�Ĥ�	K!�Őё\ה��1�֗���D���OnH�5��</Z;�,|�E���V�����e�+S?��k]I��y��ϖMi%�.F��̳��<DmfL���'^	S�#,,�il���А�yp�l������3RCcxۛV�#j�n��w��Q�3qEEI�~�Ee9�9��V	QA�Z�Z9���G�v�
vT�i�����s�j�w��W�_�/��V/�F[>�r��7,dzdX�O��a���M�b�3Z�Ʋ�X�nq��,�~�!�z�N��g+K(�/��?߮a�`��T�ls�7�&C?�xD<V�zJ  I������>�8�V^�C^�Rsm^�6�s;!�>3�?8{�N�Hx���S�}���a�$���jq�7����0�/!�GEQ��^��O#��g�4i����{��}Lj��5��j���v���0555B�����\����ͭ��z*����������2�@`��Ocg�����Ri����.�[�\�?S��r<:]�4�5�j�6(:�ϴ!���7�D�_ϝd2�5Hetc�����a(��h��B��<a2���!��É��ڣ����
U��Ya�Σusu�Sj�rF�E%_W�>t.����3�*.d:���;��t��C'��X�Nj�����LA�{;wB��T]��s@�s-]7�ܩ?�]�|Wh����3R뽻����h�c�$�w��qyD�'����ȍ�g��O���	\tVH?$��Z��`��#�K���򟤞O�s ��9��]۝͛�?��2zzǶ��U_���9��`�֪��?��zW3����Us�h�h��)7U��|]P+DcY8� 3p�<�9Z���n���gt��X� >s|=9�P� ����e�S=�;Ϋyᘸ��På8�v�.#s��Ŷ�WY^�7{�`_b���Z���?!|`�F�c�>�;�&��Z�U�B?�g�)?���n0�E�"<L�Z��� �W�"&�k;��-ڋ�`�#�H��b+L�t@���h�?i8|�&/�﨧+L�%Y � W����0v7~V�1N�A���6+���b�VC��>��(���q�q]mㅴ�g���O/^�P����pR1��RtSz�����ϾeVTy��W�|Zu?�����,hUcˡ�:��l���m�}I♎��?�`;�ȕ���7����;�=��X�y��G�-�©i/i�ݻ����:�7n������u��$�i��F��S��t<t��3;�n�W���3���캳(��Y����naW;$U��u�^Z��71���4cS���H������y�̣�z�vd�ܔ��
��S�@�ڠ��G�r��o�E� ����V|��r�����6�9�*�;�}�¹�: �sGȅ}�
L����i����8�V�,e"��~1�_�\1@	V�2*�,7���q�W>x��� �]���ڒ�H��}pp"�n�d��7�Ot��U9b���;�`I�+���̡�kd�?Q~z�&�\]��ĸ9&ł�#����6!�4HIJ��(����"����	iD�u��]��HH;:�G� �3��{��|���9纯���@�5ȱ��qQ������	0X��Z�[Һ8�E�5�AJ���&�6;Td�@d!Bo�Nx\+0 �O�D�C���/�яJ<��
tCG6)�a����h��w���藇બ�ˑ$�Rޓ�M������� �ge=����h���}�@���'BDb�y����P�N��FdO\%�A;-;�H��L�<��B���B!��:��L�`�n���96�`N >=�O҃_�C��!�y��ܫ��gKT�T-ai�6I ��3���V%Q9ܼ���=*�����Gj u��rtmoOUʼ�⫰�M�E fZ�YΎ^�&Ԃ��{x-��C�3�SRS���%<��W�r�6f�Z��b�l"wj��w<w0�I����5$O�;�G��y��瞹��S��7I���O��5��SR�~r��-XH3�L��|�*#�*�]��fzg�ݞ,e�(nMC�����@�C��Q�QD����ߖ�l��y\$(L�C��o�'�%�yW+y�宜�7̖��}~6��������y�n1 �Eߕo|s�V&�)�i�^�J�Ʃv�o�+v�S��]<E�PP��j���s`�D�?���L�y�g)�#��b9�YY1ל��Vq��xw�A�=Ǟ�����+Q�$#gL8��'�eK\d�Y��%��`88��jl=�'L��c��tX��iY�g������]��.��n��9S��K�����W�M,��v!ʆ��Y����_=�wE�M^�w'����H֎��U�b�,yF�{u:;M3`���a'Aޭ����B���J�:���!���^2!���U��>�L��(��ps_�ʤ�h���U����eB�$t�JG����H{��1e-�����O��疈d�k��HՓ=�uUjT*t��y"V)��)#^&�{Kq���/���/��+��g�^]֩<>��S-m���u6����:��K�w����0}��5�bk��s��'��3�/�G��E �o���������W+S���k�{�rx�����U�ׯo��1�f����ym\ EL��A��`�=������SC�6e�ؾ/9j�*���x��[/�=�I�XA�k����u� <\��YrY��<�D~L�[g9B�.���%ɒ�J��Z#��.O��@1%�����7�aT�sģ�Sž�x���d�%��j�3��7FC����ؿ����o�Gå��(�/v�5B�洝 n�0k*�H�e-�
ƳzF��O��#^��O�ɬ���	k��ID�(�h�-V�����h��X��gӤ�ux��<��1���pF�F�G���y�'�n��/�T4���!+�օ2,������=bn+�M`RFq>��v4�2�_2s{��b��������$��{ud6L	6F������o���Yd� ��D@����Ҥ����I�+Z�⤔=pT�7�ب�E����9�SA�*Y��w�:!��<T�(�;<g���號��F����y��j�6���1-��L[$2��Z�Y�mN�$�Z�8x|}n�7�+Hrj�_#%��F^;׭=��64]83(�����]�l'�Y@ >�̸ ���CGv�Kf�lVe1�fQע��/yä�m�3��.n��,b=��I�|�?��{�C]yO�[`�;���F��?X��ć����?b��LAKNS�d�b	�~��ሗO�CS��6��
�R�4�)+�uE���[�ӛlA�	
��:q�;��q�Ada���U�f��
�	ƶ#��RZt������o}�����k�"�a��-���t���z�w�W�[��@:
w���(�?Ti�&0�ޜʒ]����a�#�����U�}�j�ڧ��Ơ��M�5�I�vL�߂�:���\�E�m�ko9!K�HB���XLN����7�{�u��Pd�}'w������	0Nu�?�<Q-�Rwzš�*���b�w��m�v_������/���B������	
�b�����`@�-�˧��KlqA�5�4\�&4�Q��LR�X�(����-
Wp�J�s㴚��+���F��1��Z |g�:M�� m�CZ�E��靋��C����dm��B��1�J�}�����Ë�\J܄��f^�|ز�A%�9����#��#�� T�7G�x���U:�߁c�����j�S/��M�U�Pl�3���[�]�ݔeU���M�6S6���'���!�p�� �g�|-��av[x �Lh���a^F$�o��4;�V��&��ZV�D5��N� 	����Y��|&-@�.�B���*�)���NoRP�Q�d�i�� |�U�E��.�ְ��u�g3M��m���S�}�E�Ȫ�^Y�d���ыBO�Ҿ�-Iva������;�%#�����
��2KN���5�]><�A�w5���/�����P����͞F`k�tD�W��CH%�[x.���:���H�=�Ǘ|����;�;k� ��l��X��V�YL�r>�~��0�-6�2І���f���l��)�R��` 0uY���7|��_�]�� e.�>��	ř�:��c ��G��� i~tF�j���#�v�m��♕��~i�z��L�eYh����RWa��9��g�*�/�{��0�`�=sr�!���/��-���ĩ~���Y�5W�*JC�.kw�E~y����%�ֺ"�r�`�c�a�(?wޒ�6B�I�HƘ#}�g~�p�h�H�â�h���=���4��Et]�*J��XY��m�	�I4ضu���EA���@�*��u;&M^���8�dA��|z���PF��l�{�ˏԤT�U������U(Y�o�W��j�X]������J4�q��9�5껋��b��o擇	�h�-��v��F;9kj�c�H�W\ʟ��^w�*�Tf����V���Ci��UAb��xt�����|�ѽ�v�O�	�
�.������ᓀ��t��_��'k�B�
Tɩ���6-����5𾶊ߍ�z��+�9��8M'<�\L`� $`լ����$��`&I��f;X� �L��#��2�"�w��#���
z�X��r?� QQG2)a �d�׉��㸗h���ZϔC��|�ݕr�r	.'�}ze���$:uP�s@��~�<��Q��맨�	_〄2��(@c�%�
,?�}$���`��޴�[���ݦ�NҸJ��b4��pe����W�9\ξKU�܁�fN�_YP?�2Upg6K��ۼ۪� �]8':=ζG��$Q	JW{��H�>_�(�1�2�7��5�C����x qi�l|9�c�Y"�GL(��������g-���{y!3
Nq��o�*gi�=�Ԩ��i8�h�h��&���n����C�^(�DU�3��)�3�l��?�$M>�we�	�W�&��m��0{��k�2b�F����Y�?u��g{�� �˷]�ű��"�Ϫ@�`Z��:u���E�n��J	�d�[m����Z���ɓ�#S�Z�"�����ca��݄R*[u�t����0^��p��"�7"�V�Jع��}��YĦn��N=A�3OM�/o�����Q��]����Z�s*zr�\���C��zF����(l@�]u �y������ �3֗M�G@�E��a`��7�ԭ,�����m�1��Q~���'��K/�UR�-!��&�0W�8(��8'�f�Z��k���WM��f��;lIFF6�+K&�I�xJ^��RY�kQ�Y������7�O�>]�q(6P*"1_>�߰��4͵h�Z�f]� 5����y�b���..����đ��GLE_w��v\���KI�� ��d�R.[���)f���~g�-YB��I:���`���ٯ�#����9�˝o�RK׶p�)U�_,5P470Kw��d�a��W�lr�;��Z������~���y7� �BykZC,����(DJ��Z[o���lռV*�E#��+��R�o�i��2����ɊD4��s /�8<�o��P��/���7q�}/��Qk�#2�YD8��MU c]LG'����j߲C�Z|i����f���$n�`
��I���V�צ�8a1����#&1��S�F��I���V�T����C6��<!����Z/��iA�+�|4�� �I8�]��{�Ae*��ݑ���&�J�4=�"����,~R����H#��`J��w&�[�[�sl;�kc��0������^Gz����J7�]*������n{ze�p�D��]B�@.?1���8�2��
@]�T�Q�L�qS%@���sl "U�[X���C�_�yW^o��6�T@�k���w�^�hM�B-����4ؚ��X�.�sD�C��o�y�7D�D�B���,B]13pZ��@�	i已'������g_�	��8��2]��)�E:Μ	�=.��پ�4���ꈋum8�P���8pZ� ���G�#��u�DI�����*���0��2�\����Z�zM�5��qsv��	2�՝ .O���~1i�)D���zs���,�7�_9mI���S�����l�(l�M�/��E����򆈆����\2I�W�!��Q�{)"gr��n����G(�E���PO�2w$Q9-���ץ�t�5u5�?�2F�(���0�v�l��������)[k�D��R���V̵k��>!;�̾������T��f�!��q� ��|���;����4�$����; �>��3��ؕ�
1Q�������'�������f0���`9@�	�k,l������E��u���nP�f2�͂-&�#I���yL�4�����@#ɬ?��C�rP�}׮{O����V�aY����s��^+�R�	�!�]�yX|i���uO+�<�G�#��1n�R?����C~�?+��ul�'�F��GZ�I�dc�;�{O_��xQ��N(o7t:�Ԍ!����Z{�+8C�zy�yR軵{8$лL�0O��E�t"��~��*�pt�|P�r3���6C]�nvs<Ǵ���<��Is5C��V��S��(���Q�Ȧ/07ؔ�np���/�-�m� ���jv[�QN����/�J�G���)��'<F"`å'��^���_7�B���/血���D&�MM�`4�s�+��ڷ��;���+]]iq�>�oQ�[�0|�4Xo�.�u2���sF�P�Ip��|-�赅ۭ���^2�hPA�t��	��:�ސ�7O��I7Zj�w�{S�G��4 �Io�sm�s���;����%J ��&O0Y�^�?~/'	��V�+1�v��N�D�=��� Ϊ��iɔ�%t�#��c��C�� o�D���m�����!�|�h�zȱ����LB
JV+u����cnW�ǒU�t��/�����ܵ�����F�`�.��H���#=���6��=��Z��"!Y(���C5��a�1��>`y��8}b��3s�\�]�y
gMR�� f2��=���e#?fl�PIE7�
�;](�q�M��P�\䟏�O�aǒ�*��/�CW��b6ࡣ�x}�����Lو��Έ�sGfi�Ieچ���<]$�������}Y�u��{9�QZ�f�!���6��W�0W�tZ�0hbF�7ۭ�BJ2�E՞����^�R������c/�1"��b�Ǜ���;�5^5U�w@x���=������C-��ݧ�_��/��aҭ�ia�t���^߇��NP��>�
��B�O�e�8�'Ōk��(l{Oݼiw�^�$�$�{Ҍ9�.�s�笕L�pۻ�:��Kv�/���<�`zQ闤����U O�9~���k!��ǀ���]�B"��Ú`_;�M����s�Մ(u�r��C�{G����rG�\=vf1����`J� BR�6�x|,�Tr��9j��[a?��b��NТcD���SkP\�c��@��μz���;b���e��^j��DCK�=z@�,�E?��^�[E�t-\?��Z���`�Ѽ;p��h�%��@���fg¹E�R7=«�g�}N�=Q�����i���g��c��n$6c��R(*�
r�	��b�m�����0����]��pJ���cEì���TY�ٛ%��u��\{z�k5�w{�2���zA#��/'-`�px�@�ە�p�	��U*���#	48�cxp�Aq���қ�EF�D�j=�z:�ag�ְ,�k�K�Ȫ�`�B[�M�k�|DK�^�\M�v�'�KSO8)O��Ѫ����:�`L�� ~�bį���+^ʁ��_?�j�m?�(��wѭ7�'R?�N�ܞ&���ie���eVK�5��-�J�R���A���q�=��{�m����1-�-r�J[i���(^�{/�J+����S��֖�J�7+��0�~���#����^�c39Z��HV��=>�
�D�z&��[6�(y*�c;�]9���S���V��+��P����m��sW:��h���
&�dD�ٳ�Q:��"��;��f�� ��� ���qį�$\���g�A?.��PN���{o&�0�;^��_��&��<��0�7z@��Q|Z�A����gҟcu
ͻ�8�&���܆':m��ŃO���L�|��sU�z�����b�Jfk��b��!�]�"�����#�b�St�uByo�Ƀ�%fVM��������b��-�` 9�j�veX�:�(�3��⡻e��Zޭ��ϭ?0�.u�������t�L����F�8�E�໪G)R�����_?�ل��`s+'V0�`B��c�,������xY��>_,�+���'��ѽz��ok��BL����l�&{#e�̭��e@�f��Њ�i�\�U�@������3E�/��g�i���5���S����#�SmY�<�I��p��Ì ^��.N���Y|�r�ƿ���m��ǂ
EF���ƬL_ͻ�0A�zP�HF{�!�Ĥ���h�@G��u l���7P�EzI�+�ot}��U�D^ Eޛm	��F�����̿F%-���Loֈ��d@�K�G��+�����A
F�u��O ���6�g��������MdD�����B��O���P
��@��7g�|L�@P���|>�%Pn���C]NQH�Z�ؿ������q��諰�9'�?'n���F��3}]w!J���Ο��G>@i�_)X�����)	�T�v��z�P�!eΦ[��X�s}9\��zO�����Z��r��D����=���� �]�̦Y?<�ts�/��/�Y>�b��Xb�3|��5-��W@�kW��a��5KQC Z�%�j���oM���{�&|������Z��#���.���R�U�_�\s�6 	�~��/��3��F�s�rdrbp@ii���C~א3����\߂GJ�o�:�|񥢅2��i�n73C�Gw�iO������X+c���$�[��*��4'o9�c��P�>Ե��Z�sP�PW�áEZ�kc��!��d^2�&�q���|c�x��(?1��&%���=t�����~V�7�&	P�oz�%X��4��]$b,[��'(��xh�I��w�.F��i��1t����䧉f��'�J�������D)�����-��,��Y�������+*���C7����͖��	ഒ���E�?��8AS�2��AS�b-���e�����iPPG�O���]�K���"�j���?�]�Zx?��ߊ�sb%�H /r�I�Wօ�N�?F��D�'Y�o��~A�o
��^�-H�;a/G;�B��K�򈁯�*��[l8��5 ���@�� �̊�5���ӭP��I�j<�S�ͯ.tq'g��G�aO��럧���D��ޡ�?<�z��QP>�����E�p;>�nǕ�@"����E4�޼caqh��yȓ��nB�o1����'�%#�z:93� 7u��� ����sߡ��(�tF� ��F@�َ�r4���g7�5�a�2�����Ӡ��a��3��(��'�%g1R��(٧zn�c�~���p�}t�4,�FV2��b\%
|>�A-xyu9}�X�h'�B��fm��J�f5c�,�a��M��j�=D.�Df��V��d�ؗ���`Şl�,�!J��&�*�����c���7��Ǻ�e�'� 4Zs~�w��~��1h���x}d@1�0a�gV�e<�}��9X��'	`͠%��k�4А����ܟ�g�n�rr�f�Qd���
%�36]�������w }:'�j챂�H�“+���KQS_��I��4�IP+�وn��ZL�y��Fwa�����\� �� ��-"uۃ/0��%�R�ߟL���ý��*Z��R�$��WC���Ƃ�`-�;K�Z��'�Rz+�+�x�I��%~���=����7��[	��e�c�|�p.��^�:��G,c礍��FL�d�0��o"�Vْ�Ē�D�����&(�sK
y��ޱ������:Z&]����y�"_���
�IvW��=c��֮�~x�p�	k�"?/'�XP"����@��%�{�Z��
37qL��� t$�%[5�ȸ�BXG��a��ʭn&�-i��W��0����j=�,j�Ё����T��!ڤ�k���Ld�_*/�
�Y}����!���8U�?S�- C�R9#�C�ڃ�; ���H��~��,Y�b�'�K !G�#�]�&���#�^B�S��6�G(��0��� ?������Y/�Ͼ
{�@�.�|�}%[n�Ш�V�Zdd��^���������_�I1���\�����I�����a�o\�����'Y��Rh휦J�S��@d$J�nc\��:��=�4�d$�%�����&($�	������\�>�hG��{�d@)�R�銿[���ì��g��4��_|�a��S߃�ƹ��#�Zr���U�{H�w6���퟽�E� �b��`^9}y�U.[��k���G�y�n1f��򋭏���$i=f�Y0����<M	��;�OO���8�WJR��Ɋ ���N�a�ymYSn�Q�%4^���}!ٞ�l��@	�j�f�2�t��|���p�"S
A���"��?��$�T��|��k"3��}�3}�YhzR�wyV�_�8�IӭS	\[���+[}�q�?�4_��Faf�p�3��N� {5dA��#�Y⻰�ʽ�@����Ҙ�I���k��q�J�A`e��k*T�r��V��:.�=ev�~9�{7+Y�?�b+��GR�%Qf��p�Y�	���0L>�?�)�o���5ūI	W��H��K����\y�lXR'\�ђ&GQ�3��O��.�+��&M	����I�����CS���{.�-�m�y��ڐq,�w�S�h��=����公FF�YٗS�0���= D]Rr�AB���+�����q��F�̟���P��n��Ex��>�Ȋ����]�*;B�0�&4*!��?�n�Դ��N4j���Aikښ���o4�v���F�)�a��#�{7�4b���6���̷s垃��@_�9j�S��K:�0+�*ـ�����Ԩ��Ҹ�������L���e���ty�Gd�V�4Vo��8�`�1p{����;l�-o�2���l�@��������W�+�&;R��'dsQ�ր�f�6g��f��\M�7�^+,V�螎G�P�B6�j�Hs	'�O=`�S���������?R�^SY��?.�m���l���c��t~��R��C�1�ɔ	������Z�yS\���5{�)/2���GM����lOOϟ���;#��%��P���w�XU���)�cq/���b�z����(�nO��S���h*�R���$�Z?�do̚D��Q׎]M�����;�[Z�c��5MM��n�����=-I���.�ajG���\\\�i"������zE9���4o�R3r�Gژ�x���wv�j1uD`�{9ik=��N;�n^������zs��k��\Q4���b{Z���7i�4��;ssrv�5�{R��zE�**<�8����9G��^?,6k�4�`�N?99�GP�Z����/I�����e����xCI��t#[�;�H�<RUu��M���aܝ�Ss�S�ʳ����j�u�N#��\ثc~� �r����T+������x?!\G�t}}=A3W�PO_�+�eS��7^����5��k����z�����
���H����3Y�|��ze��_��Ck'k��\n�H��H{!lS���(�/*O���^,'�3a��~-�x�u�+��zӯ<L�W�?�R�����ء����}�{F*J=_�ZSS��{vgc~�����,K#��QTF�t�'�x���1��oiG�;(U+�4%��������!k������F�G"�٢���C/*w̳_G:;u�]].��	��o�i��,M瑌Lv*��ۻ�ƭA�_�~oߟ,0��q�Fy�����y�f-��|L�pd�(���:�3�DT�\�h2+�MKN��FT��-���7���b7�Y�E��߂�-�S����
/��8��u3��;;eHlYU��R��=�����KT;�����\�VEk��f
���x�s�T|�_:�i��.:uɎRG�z̮о9���Y��������*)zb��xN��j�ϴ�� ?�ϷQ�Ϭ�Y����0�rL/}��^�n�G���6!u��Þ�줞��f��k?[[ۻ7ꩩ�#����Yv��v�pÈ�4���Z�K��\#ێ��C�0y�iQ��*Dȟ?��&��J�:�:Æ1�w!���,��薾�t$(�f����J�J�stp�o�j���#	��@�
	UOLL�>*������1�Lg��`��bN�77��DD�~�Dܥ)�Yb,::І��h�:�" ��?b����8��%����f
�_O��ͩ�C�,��^��>S_�iQ�y�ض�9��M���Z��m��EB@󻪄A�WB[��x��V�B���W�ߩ��N��>��P�z���,��EEE��H��t�J���Y���KP��Ǎ��{��3� ˜5j���]X�t�|���Ž������;1zo ��k��	�9����TM�=��u��Ы���������\�!x�������������{mj���.�1��^�hVY��k�Au�c[1I�!;�e��q�dnnn���}����F��A� �חzڅ�a>K����(����]/�����߶���g<��2��_�j�[�w�9�>J�^g�����^�BzQ��?��{"$O���&&�'FG;H�(�/..�����%<f��/,��l�ZL���gs���y/��bk�U��Ht!�E̴��}����dE����R-1j�(��M��	�D�����o�ބ )r�:�FLL4�.�=����P��$���	{1��R���3' !u+�+O,Dvk�r\%���cg����o�}�|
uJ���[m8��K�q�.�-O�Qg��ã���++V$mn������[Ӎn��=I�o�*�n��9�	A^��Zk_F��[�*��Er^t
�U�˃�p<����G|&��Ferr��6�#�����X"�g����EVI	/]D{C���_�ۙ��b����1��_%\�Q�Xy':/^ܯ���x�������������$b�0�gP��}�[LN�����-zx8��M��ҳe��l0`j]�/Vx$V>[�A��VNHH����TQ_�ܿ�Y���b��ITU*\H�0n��G��j�D�d��f�uD ��À�@,�����RI�׿K�������z�#9���⥯��a�����%v�׷|��uv����|��BƦ�$D���i���~\ZZ�7�HKiS��i�!���ו��d��sa0y�qWz� s��uT'�I����;��*�4�b�Kc�o��yֿ���:R4�u6cţ��ы>���#s�o�x����Tw:9h5K+�]w�d��C	�>�P�����p�̩�bf���u��[���Ww�����������:#-�X�;5b���=��%cBW������Ħ��ϵ���ݰy/&���cP��W{n���m???W77��>����v�~�ā����Ǩ�I���{Q�M�� �V,�ݴ��G�w��ޔ�~�6? 55������ꖸ=�'���,�d�Pb׵$�ؗ�_���5]l�5��vR��vd�,�92j������N؜pf��4�"Dy�O*o�n�p��෿S�8|�>���>q�T�@EW�uoMQ�Ҋ��v���ڋ��Ĺ�eKXv��(F莛��@���HZ��+ۻ����XL�|�p�"��1��S�	����[T%޵�����"�6�ޕ�n�(S�{���H�9��;�������P[a�f�--Oߌ^x��<����WW_�H��a��ذ��������E������2i�v}�D�:�������v5���ZN�7%��ڨMRb����G�]AIIIϮs��^�z��	��*��;�Og��ԇ�"7~W�M/�dSW���b�kN�f���-i���#O�k��K��1�l����n�Ïxf�h%:>��1��I=Z���3�:TL�=^��\$���Jl�۴-��8�����f|q�6{m��mq�H������Z�q�Y�S�E�l�|ee�?@Y�x]�Y�?�(�ξ�8ۂ�/�=� O�y�p�a�p��;��N��0���s�T�����ᯆ�>vS5�$��q��tǋ܆]9_},ݰ3�v^4����_@Ș�;��d'�n�S�a���f�ԁ��KKK��k�𞕧x�G����N�t����0e��>�Ac�6D+`{�ݻ��ulz1\��b%@(|" ߬�8�E/�$F-�W��f}mm��k�
��:�+�1M���rG}��ŃzMK3��^��ۦ>��l?5�z�:�uHs���/]5sd��,z!�w���u��r�o�˗u5�I��E����cҦ�\k�����(�&,����7p�r���~̳}��'K��0r�疐�9��gd�C�c����-SEB�[���+�o�74,=Y���H����������]щ��W�V�g�`r��ͬ��!�����xԀ�>��<N�{RQ~~�YGGG��z��y�yQ�r��W4y��ӣ)�Q�^�w�%��5���ā�)�ی�Dy��i�F��aBb��/%F��P'`����+"�	�%I��תޯ_��M���;�?�}���uC�U�&Q[�W�.v=��6t�@�x=<��X��R����#𬮬�����_�+Ab.l�vwb^�"��� �;�5�9��ƖK�w΍�T�7�AW��g�6�"g��2��$����
��kn��LMO�^n��l��"cb�D=j��w�����6��;��]#{44iMT=���zw�F����;YdCr��ǌ�����?�>$�|�����:�}��H�sQ=�4x"Ax�
G�?�Hs�do9�D��&1=�N�ȸ	x��QfnmeE9U_ݻ���Ѡa9+ێ)�,6�Zd��?<��^~���=�2�$d��o��4x��z;Y��j��y���)~U���?k�b��/��$w?�6_d�C�ﯻ�yv<&�,*^��s�p����ůѝ<�:}�SR�"�L^(� ){�C���6�&X�>���9��aϕdw��f�y̷G�,�g�xBP�P�n���?��q
%��\`��n�.��p{��?����XPP&  p����1��*<�����mA�v����稅�F*	���xû���Ƣ��3��� p0v��Q�M��̥�y�Y�&��������>���!���\y�U���͛��]�|�?�ğ�G"v}���@�d*�ÔQaOD�7v�T%��O�|Q���R.�G~����\(�s����N���W0�z�={�1^���VPP��s��$����۝i�lm����+�����5��'r�]���?w�+�<P���V�'��Үɳ�������C�1��9��-t��/�fsy2)Lf11Ռ�Ч^܃C�m���O�i�˹�d���|��[����F[�B�<�(5̣�閈��&�@���������Bn��7�M1��mD3{�I�3�+���&Z�u[d�*h7�⻔�ݐ�bN�r}/��X�)7\N������x��y����D�KuX�
4�֏��g��@��Yh��!d�YG��G�D>������M�km����*�}���=��kI�)���e��	��`ؓ� ��5�>����iE�Pb���gӪh������ދ<����M�-/U����Ov�Yė`�k�B艂y��_����_`ee����M��
�E�E�<^���.�`�!WNwĶ���'���w3~�\�m�x�|K�?�p�$^:��C��'���߂V%�S-�"������[Y&��<@��vl'�NOO�4��dz+�'��,
���O��\<��o��t>���A���Ai0ڧq��J��\�-!�0U�A0O�ܪLI��:���?��4<8�A�ac��Ǳ�~�}C�Ц���R�D����`�2#�J>�v+G��e������62q��F�ʞ���G ���h��?5�C�d��ck��ZG!6��+�ܒ�z��'$&^"�u�#:���3LD� m߳,�S���M(Y3}u&��B"��Y�w3�d�����c��c�"��Gý�c�C�om�5B��ɪX`C�c�c����,�"��@�{�\�8�I��^=����!@ή�ԏ���������[p>��NG�Ŀ��@I�w�B�����JH�~�\��H�$NF�]�ѱ������#��\�/�����g��p�+<Z�J��%�y�9[��O�Ͽ�Ύ�"W�-�1�)=]�W�ٙy�#.V(q�	[k�m�ıKٰ���tw�qX���ޞ0�반�<u��z���	F��ߩ:�!�`H�r���ȿ��=��=R���[Z����?�������|Jp�l�%��8���|id�P�2�۰��NΤ%����V�]��]
����]�^T`��F�V溗���!/>BȐ�f��j&�v�`b���>D#��`�}r��$e ��KX�݀��Y�tӣi[ȇ9F�=����p􂊪����;��f+�ED/lO�\��s#��<�I2���f �p�.��oN��-���qه�_��Ɲ�M�w{��r������U�M�um�̛8j�Z��ɷB�_�#��)����b�Vu=.��f�x��r��1_br8�\�pZ�-x_)�{��RWWW�5���޲��a:�e�$ԑ+�8���;�v�4�Q�.H6���RM�俔�X<\1p,>G��!Sl5���i.BBB/t������ ?#��q��˗s'���I�y�bv�?.:b�u����}�u��}n..
^��.*?�����ա����D^o�-FF|C 90̷2)���<�9�U��s�}����Ғ�w|�=P~��݊�x/1�P�J��1�� �V��[��l/��E�EO3.�����y�O���h���:��פ��ػ��?�x�=a��/��]����H/�^�[A����*I@3 ���,t�#'�K��3,T���r� ��cgk{%GQ�:9�5���!k���0m���Y�ǢN��>>&�� b��l�1�S�L��:fU�����z��AK�0V�7�~����q��0�a���V����")�+z�u"�Ez������{�F�ܡ��P*y,��Ѧ���)e(�ѣ{@X��C� ��U��Q���5W��1����������袼y�&(ʖ��{���=�bAE5c|�ݠ�X�89�*���ыh�O���>�K*����17�L�^���߇8:�wkP.�O���볛�%�c:�����}%�b?%�x>�k:9|�P��r�$im�t��-�t
� zEY&�A���L%�<��k���L}�p�J)o
��p��OY$u�~mZ,�����P��~el(R՞���b�6���ioo��IڡA\B����h��ȃs���*��h�+�:�@�t��ks���u�"N�l4�S���}g�P�x�N�ק㋶�"(�m&�ɥ��z]��h^^��x4�����M%vJ/c�q��	^�\��Q�=�� N�zCu����l����O�L5M���s�o��2|v��4M|�V��p���1��;V�$�����My�K�H~ܓ�@�?@ S6o�	�_G�N�b�m>9��ASj�g��\u���Amϵ�k���{�빹(MU1xyCCY_y0kF?�4�{8�jg@߹���H�S��5����W��r������x�Hyۓ�{�������Rsh�#@��x���Mv��t}���M�� _�!�I�c��]T��=+�O�"������xt�l9E��Pw�k�l�e�X:�~�����^�)=��nx��x�,-N{ɓD!��6!_��8V��D^�L�0��}WVD�/G��=��)\�!�91��ʨ��k{�~�l����&���}}����k&(��RE�W���/m���ܠv�bi�}u�\^��ٟ�3���1W��!T��j2��7w4�e�޾�r�q3��������L�����X����*w?,�zk
����	n<ī�6�KZ,-hw�E�qUii�4XM_�b���8��w������3B���U^���L_�&,�U����`p8��S�ǖ!��?5�TT _��9���d��Bk�.z�ɏy�Ĵ�6E�D�ͻWFy�t�G�).;'D�6�I�k�ɾY�:�G�ܯ9z�.�g�»���r�����|`bb��H�{��f
�w;pPt���t���72�������3��6��n�4co=d�g���h�Hp��8��T���o�l�}���)�R��euB���7����&��	.�T��񞄄�z��FLP=�������:��-�PSh����Lo�y�ٔ��i՛}���>�<���M��kaU�/��s��&�g�a<�k�*�N�;�tmԻw?b�Au?Y�L�3���N.Oz�Ԡ�LLr��nsS�蛘w�-o��4i�;��s\�> �;�}���t\[����Tz�v�DyW����}��Co=�P���u��Dٚi�:�
��wWFtt��ʊ��ވ ��<*��A�����>��oȞՏ�w��"��%�=�Wͨ�P�f�A�]D�>��V���}��⏆����'��R�ξ�ua"L�E[ƪ�l���̞ؼ�\p������
�Q~�~.K��ظ������1��QQ��ۿ���7��HI��!�R��� ��JJ��HK34]�"10���()����������w�������y��8�k�';#4��rg���;��:���ґͧvq�|f���R��8�  �u4=n����/F�{P{��1��Vxr���o��ZT�GU�PHh<C)���у�{�������?�¹m�_�9{��i�?�����ʟ�E���w�)��i�0��d��i��V}����SnV.�H0և��5C��}�Ў�������o���E~�6u$��:`.����u2��uJC�/,Èl�̽8}GM���vﳅ�lu�G�jۋR��I�����1i���S��	$2I���K�u&m����:ȕ��e�?�4)��`03XXA5�5��Բ��?w :���f*Nkq��+hX�/�����H��_����c�q��by�p����y���w222b��h�$
���p���g�J�z�-�9o�κ������h����3m��2z����|#S�ϛ���I�%�CN�ց�翫DZ�o�;�>���(�͋�������ᖨ�X�%�����l�ǟ�Y�A�X��%�t��q�?�F�o�7������aC�x>��Ϗ���{��N(=�'`����rRd}�zcC�9��pa_�@HN����N,�ٙ�Kv�j!T>��k�ʙ�x��y��,���n��!n����K��o��8rw�D^L�����jq�\gSSS{BBB, ]��!?\�@OM�A�͒>�a�o�j���b�bK���'yȏ@�6��|�{{{>���|�aY���hMjn(�"""0�g�s�
�H�����Q�Ǟ������4��崯.�0r.l�4PDt�6yM��N�/������'��n�it-v�5��26��.�k��w�� ��z����}�Y�+I�y��N�n�g|s�o�ɬ��'�6j�C?|ap8����i�5/��b�f��a�F���Z��.';���vuu��Ș�}i)?�0|l���MMK3���*+/O�`g�.A�&y�{%`w�X�W��� 3��+O�)�{��uq]lM�bgտ17���co���ppp���4�_hQK� >[�w"��l��a�5#5ՠiG_��S�G������=콜!-�~��@�F�i����f�q����:aG�&>k�KcF����_� ��Y��oo画3N���\>A�.��9y*��㧤,���PY�L��^�~gl�������i�������[jߗ*ֺ�)������W|o��|��uR����O��K��K�X3B��3�<�ol��~��Ѝ��W������YdZg��s��z�v;�����|eӊ�0FF���1��\M�R��A�U.��
Գ��ߛ��b��3B�	ZA2-�c��tӣ�v��ӯ]B�lRG?�rOz $�ڟK�;:������jk�����}ZC�oj���0M-�fO371�����D����Lod�~(�E�@�px ?#����&Ro֏@יkR�P�GM�n�8��ӳ��᷇�����`�ݬ#5j7����YocYx�b���%�4�|�F��5�}7Ǔ/�(0����L���@ԖV,�2<D"r�k��>�����w���g	���\��V��J�t� ��6G�i1ҹ_���u0�����.@����9J�V7�ǎSm��o��%ٜkmF���s��4�""qOBZ*�7���X�Lx�q�SSC�|^��X�Y�'��U���ke���>3<x��9��4+�uY�;�:(��˿tw��z;�Ʉ	�7N�?��3�6��;h��a������ۈ��T�^g\��Q)oLs�%�~�Jzm?�fOT,�O#~�?;T|P��j(pY��� ӝ͖B�A�U����8��R-��Urf�Uh[P�.%=��)(5''�͕�!�}Ú�aEv��x��d'�a�CJӣ�#�k�M��}q��沺���^�9'����'������p�ƠOm}2�]j?z�-�N�M��R�QVs��Ɓ��%�������9e�e9p�Hg��q?�\#1��W��ME�E8���A��;�K����� ���+�����S��y��ڙ���o��v��r���#'��%� �kt'7����� 5�>D	xճ��PR;���\�hꯞ����7mgt$�x{���u�=�����A}�V���yo�^yً���ӗmf�S�h���Ed���9��ÊJJo�4�x��Z�i�6�3<�vn���Z����q���r{�! @ ����� ��57:�������G�:��#g�����P��K���r�S�j��7F����m�P��LV�tx9,�% �^��S����3>e����#�>��`m��}{�=�;-�¨���
�AVV��J_�D����L1��p���,@��N��8(���\�v�O��}䍚�[Z��y-;�Zٝ\0�{��i*aWĕ����%���,�aU�ZC����y�W[��P�;�,~H^gO�ɲc���⑵+�>��f�nB���8a�!\�sL
�����:R����GG�=	�=��丝j�![��&�&����1���S3%+�*��ߍ2K�m&�'���6U�[9�}�m�/���>���w9�]���0ͨ)n�%�G���sn�;��D7�Y^���d$$�c��,�E�zK�-�!fx��x����H̱�ܴ٢����'���ٶ� �L�:"�ɉ��q�2�B��-�xH��;F�l�l�/{,�ɾ�Ş��q�m�d��w��O��`���p���[����q�������=׸�}��X���9�W���g�T�BS�46"�D���Zc86$��E��o�tn �=w:��b���{�y�`�p�+V�/n�,�J��4��ը ̾�����C��\������9b��n�Zh}#�:�U�Ӟ�A�3Y"�eC�z�[�=U�p����I2�w���g{@�q�	.�x���M�X���{W��neVvF��s�<纒�y��c9Ӟe�"�v�j�o�]5V4��0M��l��zkG�����6��e���F���E0M��
�	�,5���>�:9�f.o]n{��K���删�����ި@8s��[vv��w#!���l'�E�J]ړ����|�_.��諕!py9M�����y��22�WJu��^�� ��^��~��� �=O��*p�d��Sw�՜���qg.~k>�I�1.�qȀh��I`����\3���^{������ė��W�J���&��Fc�9k��f��e�Ɉ��u��q<�w�hDf��F{\�>�ӻ2̞����득���+�6�[�1�iy���C�j]XB�KqL�gH��9�c�c�j��[GG��_��"lu�'Y���f��ެ"G}����v�sY	|#�\�;a�߳wr֎|74�j.� e��r֒7���7J������l���<����>���>�ē!D�7��}5�su�g�w�drȯ��i�T��6�إ�S�j�8R��8��L�ƣ�Q$�Z���K��ǐ+Mt��Xo�E�՗`K|V�Jlo�:��ͯ��g�El��6yl7�p2��(]S���K�C ��yW��<.��4RE�DGCi&�Z�z�@�7���R��o;&�\�'�1���K&k�A�i"+0�UI凯�~��,To��{�7;fM����m4�q`�VN�M[2��7z�]�[�O����cUQ/㝤Z���5��@|�8DMP}O�3��vc�'�l9p��b�j������r�R.�������:ј�1�H�D����Y���B,J��$��l%I89|0Xp��{�A��d.iC�[d��<����J����y�R+a"W����?.&�4ך�(��B&;|�;ﾐ�Ȝ�	~a�HGi�<
ʍ݄�����!����%� �-Y�9}�L��ua$xe��qDn�c����?y�}�4%��o5��g`��4�N����`]�=]�~u�o٤.v�>� �w��lCc��bH�O�$o�"Mr��T�dOWX{_���"��T�HQ9$���]��	��f��IS�,B�	w~=�	�?[�	��%D�ӱ�e�צ�8tKfѠ��j�x�����i� �x�1X��8֌<B"��]6ō�,�qRa��^6��fi�Fi��ݤa���_Y�~5�~�a���K��e�0v[rI��]�OLcX|�tp�83kB*MLL��U]B���R��X���0^$m���G���P�fg���PG�WD�
*Mu�r�`3�b˟�j^K�U�t�欣5���T�n����e�<�*��,T�i�f���u��$���oN������DD1P��5����^�`j�0��+���k�S`Q||O�g���o^���+ T�����y�=���
DJ&�OB���͚������Vi%��a<֡�t7C����Zg�<;OΖ�~
�DY���^f��,3'��'����98?����D�$u��xY$7Y<sq~�AJG<�U��m�M���d��w������$����M/�20���x�jZ� *,b��Lӌ�GJw0�CB����p;���ٝk�y�1��p<6[���ݲ�6ޔ��Y]��Y}��ѡf�Ic��d(���
��7����K)q�6��QK�cC�h�V�7L<@�i�e�?�Ğw��+�n�k���a�0��p�D�F�?�"�} i�⭎�Ԝx��?5Π������̈́-�(K���DkU
%}�PV5����{9�m���b���,<6E��қ�!��~d35�(�ݲ��������b1��ao�<7�bm.].؇��hR��ĳ�.w�5�I�b�$�u�Gگɴ����S㍃E�j���ܥ#��8AN���K�4;*`Jj�4Y��Q��F1Mn�U��QΉ	9XW7�!��{a����Tg�ֲ�6�Y�
,�z�{l����3���F����r��)�	)+Aɲ��K>�'�u��q\GF�h�Q���fSԣ�/�-ޖ}��Ķ=G=��ǫ������OY�+_+H|]�>!�(7�?0���q�2r8f�=�\�!}��C�S$V�kj�j*�d-{Ù^H��b�{`U��W�x�dߓ0p��e&��98Ǻ^���-�Q�{2�m<�g���0Z��q�s!�)��.V�.�As2bu&�C��X�@:������(\��f� X�K�Q����WV&>�D�O)�
�2�a?�O`{Ջ���|}m�18o[�c��K3gD>�
Ԡ{����^�4@�B ����/�����DҌ!
N�S�#�X��G2�h��&��y6���[,�QJ9u��\p�W��3kY�YD3]�E�z���Ü,�t|*A=x����-�tnJB�[����o�;4���
�~�Ճ���`�0l��s��d�5�A�N?�NxP:���ת&/j�0�U&E�w�M�4��]7g�w�Y����S�v $^)A�5>_[T��U�e��6�Ȃ��ҽ0��J�m}���r�0�C��A�WC�Y��s��ꃝ�{'*��s�DEC�X���!4	��y>�����T����N��A4�Y������w�"��>Ђe����#m�3t.
~(?�`�Rٚ�/��**��7;��{������C�P�2֐�`�m�2]A��J��	����vV��]�T�n�tc|����������%��L�L�|}-.{�:W�S�2�<KG�sY*Pu���hK_�>�@Y�en^���[�hG�ǃ�WY;��$b��l�c�鞜������,��L�e�aY��[1�EXn��D��ƍ�Չ���h@����|�yp�h�x$���Ӷ�g͢'Y��D9<�u���,ǲ�m�Mh���z�9�o�\�i�:M��y��-��
ך��2�;Q/�UPjC�+7T��=\HI2��k��<Ђ�&�fo�S�L��4	g��(_��iD]���5,K���������Tȳ�Զ���0d�m�e�>_
��' 6��d{!=ɴ�%���x��TX�C��ޅ\7��83����k'�\����`w��7�=|sN̲���d�����5�uao���������EC:M4s+�0J�!Ҡ4l��|���B�W?*e5�J��g�ܟ�Q�bȨ��F�����P��T��>�U���[ʘ�wlj��W~�8�Hύ�ъ�&���q���� �u�Bt11��*����>a�2�r�� 8!b����0ǰU|v*�Y7��YT:_x�M�s⮉i��
m#I;�.�c�g�o��!�%���Ey!����V����P>q��Γ�mn��*Ij���	��fi��Ȟ|)_�>���V�w|���X�Z�#t=�6
c��
`��"�Ь���s}����j`���?g< �U��R���?O ��|�{i�}��S9����K
0h}�lܖIFCZ���|��gI|�O���p�AN��,��kkC��R�~����!P1�GZ�U��^�ա��W]�~JF����1����Sf�m+D�i7���\c�E��z�3��E�;��?b<�o��{a?<�h՛��)9\h.�E�H8Tm��4o��?t�ت����߰L��U?n�����L��,"DAlVz�|�9����Ō:�<1I���x8K�������!7�A�d8mڏ�r�b|���[M]��mo6t�����,��A�'�w\�GJ${w�$ M�����N`�P�y8��%:��ϖ�/�������
�Qb�XPt���l�N�����GL �� �Ș	?�r�:�Dk�Ȟ�[�
9���'Ơᮐ����@�)�~��-��-r�d��w�aه�_ee�C�'"�h����k��lD�i_�'I脩iG�q��j�TӤU��%���ȍo<�q��$�d�梷<�b�y���Y�Y�HR�>�p�%~��*طo1�0�B��z4��@?�I6 :[(>a�i}�#��u�����Tj4���-\�w�Q-zPwqR$v�I��F�]��9��2˽9�@ ���F��XE��%{;������<f�c������Nv6��&P����m��!��C���!�࠸��4�X��%n�����v!Qf����9�oq�VZXw��	o� t��������}��X[��-�O۾5�M8ZN<k��%�4���/f��3�*|-���ӑA��YT�*�K@�H�\������a��CG�ܯ���wm�U��eK��.ۗ�G�πz6x��+���AXD���f��=ѠMS��bu�W�4�蠙��i����Hi�?;N7,�,EI�mq�~�(�kE��?�����2<���^��QkQ|IΨ�"T��%�����>�ڿc��#�:��0t�����ǹ��ltc&_J�!Lٖ4r����ZT�isY�����U��4CvKu,�!��@��j��Jƒ|����ν��	t?�L}UϺ/�ew`�����0�!������ӻ�ٺ�$�SI���Z�w����g��D?��6 @���:�w�j`aS�i��o�\�	����v������{�����Œ?ҩ9zW����P�Hf�s��!�ɖKT�o�!�hu�o?n5��#�5E
��f��F3	b|i���~�[���{�Ն�
N+ke�`8�~��u%�8]EbWޭN��=��I9A��V$ �JH�/ �k��T�0]����9�Y�"{8������� {S�:#s�S��?������"&�d�h9�
�h���L�� �B����w�9�Y� ����m��CԾ7�wF��sc�;gƂL�)M&�P5�ﾾ��nh��W4��`ԧ�M�#��a��P��w1�� "p�Nm�2��)C�h ͗�i���I�=Y�IV��|�k�m�X����#?��bO4�{�㶿�W+�A�q��,��-	S˟���S�NQt-��a*A�ۇ��^��+��xT��o�A�(RPn�._�H�ܤ����!��+I��,�'��`���J��4�O�Gj߈��"���߬Csc��ڮP,	����b��r4�S�t����NIޔ���*�3�WT��0Q��e����zY�9��{�L�cs{��*�T�]N�d��&	F�>9�Ze��JRc�����p�Zϑ�u����4�b�+M�.����͈@�f�r-�E���9j)R,��(��;��J�i=E�[f	Ǳ��%��3���C4�)�w����ݺH�����$�<�^d�H�'�'���W_ё�c�]h�M�C@��t��<�.,
���%� �S�e����0
%�0u�&�f�W�^6���a��K���}�^�޷w���.ܟ�md<���U�#��c���E|��Q0=\��(0յ��O�i �W��>y~�F<���݆���t���QǏ>���ͿZ������{����݅ÿ��E�H��˱0&,=�]�E!2�5L�&d�(��o���(�&���VTud$�� |���̏L2� �x��x�N�a�&g��`3H7���
���עi?ܪ����ko ���@��sG�K���#*��L�����`�1�J����;Nd��,�,�by�+nU�[�l�����e���x����z��:w����)y�L7�>S�!R���k�R��H_<Z��pr@�<�H�E��	i#�=�$�Ƥ
|jS�E�*_����2c��Ɯ7���(�5A��P0�π�|+�҂{�U}���n)P��zT�]c��x�����#�-*@I6�eե���Xz`i���T��?�b���]yByϙ#�1�n	S7�V���Qwm�Fq�I[Wt���IL�;n��) �
��y�c��<�C  A��9jI�:8j��0n����j�"��ڭo�h�=�&X�)��̹D���+P-��	:ݖ)1z�]�j������ѱ�g�+ǔk�T�L����@��JP������X*{��hZ��`N�}����:о�mr�>��m�1�"�M^��u��:��M�X�T{S�<��aN���4�j^�a;*�yW�NÅ�*͇�\��cw;�Ez3�8%h��ꏒ��r%L� �'��Z�k*&49��;�y`,�Gk�E�.j*6�K�u�.��s�e2C�E�B���h�5��V��e�b�<����G�8�[���BK2+j����pU�\#��Q{���o�J@'��$�kS㊚6�Y�/��=T���󞡃4B���EU�A��b�"�{������,+EO�	8��1۴�"��œN'@�!Q,�{`.h8T�lk��r; �����}�x����R���=�U�t��:��:���$�ؽ�����^Kq9g��� �z���dG�-lx��[8�M 樤�M���9�	�	��:7�ks��2�<����,ʉ�{{{0�'�k�����K�����9^Sgj�q�e�מ��Z�z��$��r.��+��M;�{���=Uf��:�>�Ø."������n�0�ݝm�F���N\F��Uu.��g���[��hJ�ۇPk���6�xR��mt�� ���uE����3��wp�@y�h�xY尉[t�#-d�_%f��'�j.�q�\ug��q��ڒ|ۀ��T>*{����B[���pB~V=��?�5�\�gZ~�J��"�	2#g���h<�Q��t��C;b0��A��Y�ϒO|8c���q�!�|���X'� s��S�g!�∑/X�k2b@��Tgԯ�qN8 k�=P#�墑����NPu9��Zy�� ����������י)����� ���� kdx���Q��Y kĕ�ͦ�a?� ���9��(_��a_�|ק�o�ӌo��Gd����̫m�f���@i 48��$�'A���D$e��t�K:(�3�XmM���%�'���p��mlC���ٖفFR�����K�	K����P_��	����k�ौ�WcHB�  �e�b���(�KQ�H%�2E@�L��}�?d�f׽�GN���u�co5����wQ��:p�K`�eg��ZzX��;�	z�l�d����t0�@V�\̫�"Tf�]�2z#<�\�D'�X�>�q_о��\���!{Fa���%,�G0�0ۧ1��dƈx㋁%�	��\5�>Q� �Ԭ���K�u�W�`JT!�篝��Q�<E��Q�'�e�M h1�x��%,z�_�y�z��N�'��&BP�R��_I<e��.�)��>+�v��_Q|�F'�8iLi٧T��.{�(�z]鵥w�zˬ
e�\�n��_�Ԧ��E.�F������%�,��`�(w��$��<������	����L� ���^�����O�)K﵃Dm�Od�@uiV�fg�n��:h}s|�nLT�T������:B��{�� �f��i�|f3uI���+�) �ݤ�9_ږ����ut�v�� c4�}�/G�ʻ�+����s؜��Mݬ���R�^N_��:޵شno���ڧ$*�F�B}���>��D�%P���f��V]�r��S2	9���{��5yA��&��8Y�fW�"�6Ԧ�S��!��5��@Fk��=�_�s��Uz��P�Sh�vR�i�;=��6Np��'�۹�Պlh��h�t0z>�OUF昀Z�n>`��V�[���X�LmΚ@G{�f+;#|���m.*���Td8MY����kUsu~��T^����}��-��][�~��l@�#4a�^s���Ʀ���1K�C}������z��11�W�_�F�H�"77�����U'�yg݃O�$��h�0�`9]*&#\+��,␒��sC��1��gţ����l�4�^d���1��1Y? ��C�})����qÞw���R��`�)+O��3G�p��
i��4"�"R[ Q�wTyYB}ř^HwQ�"��"8��'�����;�����J��#���nڇ�������0��}:P�$�jm`�˂1�f)��=z�r��i�~3�q��b�mM��}B=��Z9�Nt�!1�=Ȳ��Lo��=@��*�Har����CUFf$[�ŵ�P���`���6R�)~��U�WQ+<�����J����S��u)`�!X4>���uI�ö����̬M��b��4�fʡ?�Ze��.�l�	��
��*e��!?�"F��(�J*�.�U�Lq��Ht7�U��{97�4����K�Y"�A����q7Y�왡ps���	�*dP,�� g�5�i�@e�{
���ـl���q@3��񉢸�I1!B����*��E��>�cG�i��%5O��� ��1��/t��ʱ_$��*��+l�0���]뢛�,�T��v<By ڸZv��0�����*�)m$�����Y�]i�4 l�!~5��������H����Dz�w�S�d.�2ȥm{A4C(���Y���6F� �����mD�J�������O���ud�R�����W��WcX1��3��1%�er�e��&���膩�j��\��6�^#��8]�}���!b�G~I>+ �6��nX��Ka� h~�S�ʩ!{
)�S�����		�;�q�Zz�b�a���-�^�F�|����}��l4�vsX�Eo���2	U�� �"w-�rpC�Y�<`����L9jZ%��W@��f��h',�rÒ7�����P��#��P��0JM-c�w�P���n�ޣ�LC�����/���T,��D�/%r���NݛwC���� M��~�&Y�q���o��}��گ�5�c��c�y\�� �,Jz���H��,��ժ}W�G)�`�k���O��Xݺ�Zߜ�/D���$M�C}p�,_������O:�0%�:�B����ehS�v��l��g�/�P��t+���"�# �HyX7���n"¤�,LrB�h�f�(�����B����H��4��,�	�-��yˌ�=J������L�( ��/�G��yL*@q0?�q�O2�dv+�֫��s��s����OH�*Z�t0h<]�)�-Q�����,!:{����ʖU���������Vآ�%�
� �/�	�Y���/�r�D��eu��d(��E,�n����(xd�d�JfT$�`?0�˟��.9H�:�NX�ye&�R��P�:�Ƅ�r �V�`�ؓ>	�8��b� U��%�KF�2��F����wpA�62�i%G�@�G����Db��z�>��0�ߟ�}s��@Lw�o`t<�k�b$�Rȁ�rF�@N9ݛ4�{�ju�-#Su�ځi���"|I�h�@��TT���%L���t1`뵞���]A�V�i�#W#,(.GP ��Gs� ��k�	��x���l�)Ew���C���"v&���p�����O����� ;*M��rw2��1_1Pً &����e����H��H[;���~r���� ��O��t`x1�?�R!.��v=K��w���" E���%��[<��/N�ΡW�k��KLY#%�zrCu�}�GM� �?�h�*��W��Xy���u�Ef'�%�/������ �l�O�װ�up%p�B��#=���jݣ7�����tfz�hN���4"�SG�R* @�&�8��~�\���z�vN��n����Y� ��Ԍ$��Q�32�c_@�2T���G`0iRf��'�I��i1-x" ��_ �TV�	L��#��	4�{�E�����9�g(�ǋOd|�{	x�H��Zq��у���@/�-�k<U���Oiq%)U��)��'%Q�3���ח�0�W��̄�p��1�8��2"l�xj83�����{�8��E1u����2OX��$��E2�!��<�n�i� ��y׷=� )���.��l�F t�L���g�����[Sk��RI@��ȥ��2Դ�+sW����O�� ��T�Un��wZ{�@���6}�����@.����*v
��2��]����V��R���]�����7V�|�Yv��=�*��ȵ��mO^qrE9'Y�ve�x\%��#)M���b&��������S���et�a,����H�([� *���H�)R>[hB�����D��P�Z�6[���`ˁ�ܭ=U�o��!X�ԡ79	x�0v �i.f"e�Y�&\�=�L��:�W@�;��v*$KT"a����`���7�ܣ$�9����O�|�[L(a�,>�N`��*'c��!�7\w����7��;��f��A�u?�R�瀓���Oz�r�5��m�2_�Kȷ�ԏ�@�Ҳ�\^��n�%x:3� �.���)V�ce�u�>�g>����ׯ�NLz~����)��o���d���>W[<[��*��R��*
���P������ɲx�?,�Z��sQz�>�iU�B.��Kc4w���b#��6�`�������
p����T�'�i%uÎo�����H��ֹa68'��'�ӂ1��$�$�����8��e/T�C��"�X\���l����T��ؚK��S���^HRP�A"�o�U���<s`�h��pk��۫�&dr~C��\��>�%��͖g$���gn�t[ti{���a`�� ��$����������@�M��>^�:�t��9�q^0�)�.P�Of�M~ت[1���{�<س �q��PDp石 ��l姇p�A�1�<�e��L���iԏo��F�e,U�*��7U��h��ؾA~[��T��l),��a�i��"�Rs�u�S���]e��>j�S�OH��A��_����,zq�̽{bN�o䁾����/�	�6��{/��y�V�(/f�c��o|�3�·Oc��Z��2�S�����&]�@�y��4�����k�A�0$h7�,�I�ڵ~d�wT{L[�|�L\�vg����u���%��?�д�Q�L]�5�=�䘣�Qs9ɢ�*!��&��O�!���'7��yJ�hMu9�Ğ��4"�#*�1Ԃ#���dJ�=���
��R� ��ݧ$!\ S�Ds]��8]�+�F� �R�]� C�4��|���-ۑ��^(��1�����nW�3���Le=!��t�e�o��r'��p+��&�n���OM��#A0BR0����_mTJ Xg̞gU�̨�~�m�	X�mu@�J�;oA�������_�Ӣm`N7j��b΄~a��*U�W�O	?��pԴt��I�;���^��I�� �������E��=W���Gk�y��Z����jU���:,���i��f�h��;�LU�qt/v�~�m�������^e�
sT
]`X���G�x9��(^�l�B��>��_d��c �i��h�C���l�Π�G昀{�,�����"���0�Jl/@6l�p1���L��Ĝ&��(샽�	��tX��~���6d����i���Wgb5�v�>�Сࡅ$%�������S<�[�!7��� �5BSpBqqP�5ᐈ���~h74� |��k���^��H]����JҺ�]���H�W	�t�X�S�Aɷ�q�����硃���R�VP�y����l4��Ѓ�%�����ٜ����h�\c��,���%N)`\P�	��avB3�ɂU�Ka�:�~�P�8����� �b5�s����,���o`ϰ�<�°���dwP�_���X"S.O�~��7o�R6��q\�����1�2������y�����8�����ICr��~���.����۸B��(�T]ݹd�W��(\:U�볲/`���RV^,O���7?�K�Y&���)�?��b��e���ցwf(��3i�u��{�m�ϕecc���������Cٱ=sV�[���r��٨�'��\}���ɰ��&&���n;��ˁ�(����p�&Q�t��
�+��ؾ���轢�+��B"����s��Z(�ϧxͩc�'e|��#�:$�e�2�"sZWb��DFJ�5��}������������A�����T��B��r����I��Y���	��n1���?�hAa������1S_�P�
�LaK0Q��������5�k���Aj�k�8��R�_�;1o�R@���i�c'�j=�(�V��WV�
�rsso,--�}�;W�����mt��whc9�Ⱦ*3������=����L_���ҳ�ݒ��"n��!��z+_����N:Բ2�9��V��ow?�L��_̺�|ִ������胂�B�6�Cx2�.85�[AYos\f�����yx�8��։+$�|�?�U,�8��2�����a��U��=�kT��g�j���b?��LOOow_K8p�]��=�ϯc��14��;����w ���Ӑ�ਚă�y����^K�7�&���ْ��p����V��-x�ߝ/�y���`i�C7+�F|�͕��i����1���������D�_~�k�������ۗ����sn�u\1�=H��m��8�i�C���")�4)�ߴ�"4I]���W�煱W���`硅�"��C}%�v�l�sϡ���ŋ��z�ī���I��q���3*�0l�I�����[z����smF,�r���χ��ҿ�o���i��k����]�������=�������ggeeS��q�ӏ3�),m���mфSL��OC�d�%dB������kzR�WS��#KIRM�g�W�T�NN���(�;bȤZ�DgE�E�5<��yoo��M��D|﷣�ӽG�NU�D��":h�"���@�`D𩆑�bT_�Yg�����V��������P����\�rJ�.9݀��1c�)���i��)��}�1�8{~�#ܺ�8�����_>K�� y��ζ����m�q���y_C�M�&�9b�&M��p��A�H���򒳣V�J�;�����\���_z�ĚSD��,s��oZ�I�q�b*����|��EK9�꾑kMw�{Jw:kB�)dX5w>x6v�;�Z���4�&uF�z�Z�tddK^�a���K�À����ybP:�.
U�?���u����5��Z~�D4fؕ3��v�;â{5�_m��s���{��$}b,'��ÍA����r�/�BaX7?�?�&�;�+_����D=�]��<�^LS�w��RgX���򓚆�t5";��A=�|5۩8��d�97�a6��F�{�a�����Z��7FNY�uw����
g$��Q�6#��:2�ߙ��G�I%�;^|�I>�Bc���]JJH��J>�QC)�%��J�ni+���m�8�PK��%	2���k��N��[s*S1��{=L���b���?��7�?:#-*7��r�l�t=#+#��nݐ�1��d��q�.�m��C�t?�>���G$r���w�W8
9^��_??�̉�ܷGKO�.�F��~�^�ו��gb�&�믘����-{n1;�o2q�y��r�ﺁ�0��;��m�ޝzz\[��R RZ3Y�g¬�·�|��b`q�������}W���"^�&���ގ�m~]ئ��_3�+g���}������,�>ݩ�vgT݅�<TO�S�5�:�k�-�,;p�]�s�2�UQS���v����3^�54����V?y3�>�����4���f�d���N�i0����﯐�#���ůZϋ�V؝���y��y�������S;m�t��)�'���uEL^ɒd�/�_c-��i}; �=^�� ��O����z����0�h��xjyx�dx�bf�R�p�QG�Ġ(y�0�6wϗ����z��+��|������7|��j���w�)N��<7��1\�Z�����{�?BŚ {;�ͮcE4��!��{��姍��[͈��'?�z+����.2�l~k��'����s�^�Z;�G�1�iIWuᴼ�	8i�����Ņ��B �=c]�7�	��}�J��#T^S�xFf��a��{�E��ʕ��q]�ּ���i���X���R�ڨ2�{���XԫcL}a9�h�n��x?����p뤅"��D㇉��ӊ��	�/V�^f?($��k\:�������o��k��P��s:G���Ӟ��vlk����X��}�>����=̖�o�#\��PI�ظ�p�V�������aLE�{�l����M�����bXd��y��y�W�|���(3��[
ߟSc���*���L�����9r�l�+�x���U��d����Z
��v���.��2��3�#|����O����d�MY��K�D��;݁'����ׁ+�F�Q����V�N���6���u8�e�����<�R����+R��5��O�:�},Y���'-����O�{���c�f�`�ɿp$CZ�tl�x���yʗ��'x1Q��6*�J����B[g3�T�>L<c�H�۞�wZ��`n��Ϋ�m��eJ||q� *#�s��)�faaф\/ev��硗�r��,7Y�R�&:>ؚ7(�S�>=�lj�Z��3ц]=�PY�����8{󸦮�_X�+C�ZEH}h����Q DEE���J�*U!�@��$*U�8�U�$CD� !DD��!L&�$�2�$$!�O�־}���{�O��䐳��k}��vN'��S;i��{5�'�'�A��97g�D�z�:�?/~FLG��h����x��S-��v���xcǪ�2/��j�7�#֑釂G���Nv�v8Q���y���IX�:3�@#��I���DD��dDz趘���	m�����O���w���s9I���7�9�!?��
y��&S���+��d�R��/M~388������)f����d�vֆ0�[q�ф}EJ9ݺ�1�f�/�7Z�Or���� ��'�߹p�T5�HNϩ������je��ܤ(^94�`��ի�k�&7n{�d^�Vѩ	I��Y|�&���r����E�SB����
h�土P������
�ք��(�#�I�W�ADcE��E�7L�Gg m�;��C ������7����D-������jI�Ẇ�������G&�o���o`` A)�Y���2�2��2�s
���S� ���Նr�/(^�Y��4�C�B=:4���s���-����u������g��?�<����d1��*b���.!���S�K����n�T]L����(w���� �eٟ���k�pM9����Z�Q'$������r�ר�ѿ��(g���qNO�� �6\q�d�Й��ER{/��Gޕ�`���;6�����9�� ����-͜8��K�ؖO����b����v�m�f�V��._Ҹ��Q�������]�HY��&Lv�]^6џ)yf��ǝ�r޺����?��<-<rq��Z��}�W0
�q�v��ܨ�:�YR�L܊z��x�V�jF��T{u�y�O���UnVā�]K�M$/�E�#���L~_��S�֥���#+y�
�����W���J�1���aک'���K6g�j=�g@H~����iQ=���
���!SY�ez�����'hs6C��]�p�#�q�a(�uc��I9�NC�q��ԛt�z�������cj'��5�>��kv�bdV%@(�
,b���|���?��Tų�gHs��� ����q�ܪz������������K�W��՗�q:��X��~=tsY�-}� |�f��'�T,`�M�ѝ�Ǉ��b���G�Kg��y<S�N��������o��<�C��%��|��*0 �2�/|������o���ǟ�,�K�/+Ʃ�K�C'�_��k�,D�!&����ω,V�s���p�����!%����!J���ՑB1O3g��^��bҒ����M�٣ߜW��=}��/��H����E�+�V�P�E �ې�r傡TT�`:���Tx��|d�U�n�¾���z�#�܅�0h`�n���iL���w8G�O(����bǟ8��OH_ƌ[�ua<����~T�G�����Ē^M�K�{�l�� +ij��͔�����c�v��k�d��Pu�K�Y]���V@��;�1^:�>W��B�=�E[)���\o��9�@Q��b:��!O�C�J_�л��q����\�	�m���H-ڇ=�6"�~��I�uF	�)m�����kI/b���"[V����V4��ea�Z��O�y��#��x�jZ�KP�Z3��׍�"͠��)�!��X���D��!ol��O�vgE�))�k������,�4�'��|Uwڲ�zq���y��KW�)'�HgR3S��x����(��Z6�H�"��j�w�?^�'���1����'
�lz��۱�Y�V�=!w��M>��-i��Pb7�Lv9**�|�̙`���T������:����JZz��	F�~��c�h��̧�5�q�{���9pG��\�T�2E���ֹ�~���ҤׯP�>V44��*	�6?h�|8ԧ|�S���:�so.}_MV^�X��,y�c�?5�/��3��IUǶL���v�^��%�eL�M�a��8�삡���N�ǷM$���Γo�k����M8ٲVL�
*�Bd��7���R�q�׃#�?��۔8���9S�}5�
���-��`$9.Rغ�ap��<��E�
��G�e����,��~���X�h���ͷG��q������G�������܀�|t��;r��#iE�E��S���a�GC���,bQ~��O����C�`M`ɺ]H3o��g�f ��xVk�J����g9=�j5����M7ڪo �J@w���<3鴀�Z�t}��b�eA��(�s��g�(�2YV�d���b�힖�M��+f��g�9���_������(u|�/o�嬬,�ŋS��1g���sz!RÉ͛�⪩۵����l�L��AJ���(/{�Vܿ/�[�&�8��pc.^-L�i/����M]�����&��j���$��@1v31{_�~7�~Ó1��ٝB��)�I�3�3�y�x���l�ҽ����n��:�?:p&��o�~5�կA������V���ɉ�{�E>�o-�7�N�4�N�n81�0ڽ����[��i�Ϭ)/��N^tvG�Mhe�W�#���5 ��g���#]qז�q�}�����Y1<Fu:J9���}���)�뗳i'}N�	�O�0Z��=�q~�#�mJ���?;�޷��}��w���r����=D�П�޶�e��Ô������Y�>�������'�c�������za�;i����O�������m������'� ���Ν;G�g�T��R#ؓGf�ǐ��ȵ��n�ٖ��R�Z\|'7տ)%)5lP�YT�l�aK������B�^'��+����-?�-�<�c�I����&G����޾o� &D*&��~��3B�9�L��C�d����萟q���2�e9�z�ѹ�ĵI�!O��S�X_=��M�������DN�Y>��of!�!~G�x��+*x���ҷ�B�X��'?�$�tglIE���#�]�>Ƶt��/�t�@L�i���r�Yٷ����(�y�Q����.g���E+�G\6Iw���%.�6���[���72��	
>�ʼ�t��w�C?<x"�!*8���;�vl,ڹ�t��e��ٯ{��S�,E��]qo^����y��{�D/,�;4�痳Ь���:���`�?}ǋ�]���;J�ᠤ�'q�V�6�5�+e�%-+���Z/m�b/D����w���U>/qWK�'�=
*�!'5���$f�:�}[��Z��8�f����۵�;����R� ʊ6:�m�Z����I����$��U ��W�f�����Pb3P�����W�( Nگ��W��ZI�V̗�3���4៞�vm�zΏm�*-Q^k�������GWݱ4������- �}~`��'���	���o���Г]�6d[X�������]�g��T+�/nO��<[�P��`��z�?�@N��߃�Č�&�νXF!��7b�(y|0=-��~}h[6k�nØ������&��xO��vm9���Z�tI$��l}�OV���������6g�UE�<t�qI8�����?\��~�XR0t�2�,䱱�l�SNL����.h���$�>x7f83DĎ?���6�(�_U���9�m�7��z�~۔+#�2&y��y�qќ��uD,rb~���f'�hID�|;K�����;�����/;o�$]�!n8I+�~���o��X��U����T?��$�|�^���?w�tݸ�5���>�~Nġl䠦g�h?�!āw�zB����Wϧ��m���HÞH^��8R\�6lؑ�B��ֹ8c��}�XjZ�I��3����(����9T�3��U�uy�[����g��N��,<b��x�2hgw7�yl�n���^껯ԯ 9�}E'���H�'�s�����p���_��߮owڵ�8���|�2�~b(!��s/�ɒ����pRr���M���2�;���-���Oҫ���d����r<����� ��L��mI��¶�MZ���p2/o��g3��߿���)� ��~��N,W=����/9�Fh��>��Ի2�l����c�2����*�y�� t��쉻#^�o"LJ'�ɐ3%�O�7_L��~��f��ǳ {�_���ߺ���u9��!ʛ��x5:R;Y<��A�o���C�˝���������0��	߆e��wU�s=�S����5A3t�0�2g�[�� X|Z���V� �;Pwz�����1�qm��y�^�瘲Ǐ�*����~��\���!v]���ا��˙��M�_����I�bd�?�L<�g�t, EQ�K������+pUv
�7˖��p'K�Z�{k�,�N�t�<8B��b}(NP�m� |�g�e����53'�ܖEDDLtn������<R����_c">�W�R�l���|7���z���!���,b�>ꤡݝ��O��:Spk�l�����E���-_�Q�gg�N��gW������9���?`WG���g�ִ�ɖ��j��ӰZ�)���d��h�	�n�g
�o^�RH�����`��]CɞN�vUu٣yR���m�	G٪�c�q�����9`d�[ȫ��1�Z; 箸�9�*��Ѵ���zX��ij9bz��!M$4���H�|lllY�p��T���a��'�`ے��mh��o]'l�TT�Ґ��̎��F���*<�F��Y�1�wu���E�/�Z2Y��&ny��������2:y�O�S���>{�}�L8�������̵w��dlu v�)�9�e1���Kb�x%lSO\���5�����V�2?j4)w�ϣ(;���=?)N��-Ӏ6����v���	k���H���|^�p������˚��3~\]�h���황(_�˺���$�#������&��x������۬gּA�Y�gI�qk���I�ez׹��lԙ�M��?{�z�,��VU�˒���R'���<W�������LYӝ(��wdpھo$�^K/Oz%���+.ﲵ�W�rK4G񿶃]���$��Y9�388���ԓ���V����[666_��Ԏ�c�����Mf~���
� ��O�d\/�y�yb�(������Ef�l�Ţ�#�v�$���+,Gr����c6�,:�p{@��9%\|�Z�9��F�ӧ�q��M���s_\�\����6�S�+�E�tև��fs�2�L5��a�9T�:��ãY�+�,~Z������mے��|yY�H��!���[�M�����[���o��*1z8bun+��w\&^�y.5.�O�[�Nh������w���_����9챌[Tzl�t��h��P��jGǗ��f��N	ڦ%��$�͘�����,�'�F3����6T�mj�,��\4~���������r��dڃb ?�W���]��=����%Os��!�1���;���������|y�DNx���e��wě���l%�(���[�8s�c�~�����/z�UJ�\;���]�c-�����ڶ��B������3�d���+ݼ}E�!�3�/9���S�(���i${l�X[l�T}9}Ɍ��	ė//Kݹ����iQ;���M�?�����~e�f~�x�Veiea8͓D�O����eI�)��lp�ԸI!����&���Z��+	�Q��}[���e���[��扽pfK�Ŷ<�� ��� cG9թ{�~V������ZL_1�͇}�!����s��H��������
R�@C�M���G9;�/���սd5}���o�ׯ���liB~RT�0��=�8�Y'�?D�k��G��b�u�2�t�`�w��h@�p�d6}�df����2_zB�ibҷo�(s]��prUG�^���UL�-/�#:��<v�ï�[>���AE��}S���yp�ҋ_�ɲ�yl�y�;�!$�#^����xk���3�:i1{<�c�U��4�e�k����?{���c�7�{��1)Yz�;;��q?�\K��-/o�1�.��p���C���K�ȇHK��h�I�{�@���zF98�aA��2R��w����]�=}X�W~vo,e,�I�yR��5��!�st�����m���!G�x�G޹Ǻ��Eq��kMn�o�(��k��w��c�_��D��S�	�ч�ׁE?���ot�����"��"�[��`x���Su�3}�Y��F��+�����+Hq�4���ю�,g������&�1\�)Ցϔ}�)g��2d?��s��?
=Z���_Y~��Y�3F@_��@������W����3�O����8ɰ�V��sC�)�6|�f���w�N��p��:�j����V���W�k?�����	�z��w�|3O{�O�4V��E:׹z�ן��"> �ٷ�oz�\��`�A5�����]�aKaci��J��Y}҇�R3��O��vͤ{�X�@�Yђ}�z�!�&P��z>8�ނV�B�A��_��r�n��'5�oZ;��W�
|����b���=�H���������/�H�����v��P1�����/��T��'�?�tA�����Z����͞ѣ0M��%�nȇ�;h̗�E����偍'�fM_0��[�mk�g5��:Xv3�|E�f�T{�C9]y���H��1 &�����ݓ�>����u?}g.�Gu8[ǎSs�5���o�L�nvDx��y�����K_2�f�z��79.���jm��k�xy��1�̷x�����f�洟��p\�\p`��H�<�K��N�@(W|]q���/���~�a�)s֨<�<뛐7�N�s�$#�ʙ>L<}�F���c�'%�m�;.0:���Hoo��v�S�~E�v�-
��<����'99�z�l��q�z5!=��oPh�y� �AӮy��Ԇ|�,Za8� ��?ʌr�uBmL3��J�~t��<��� q�m�G�F��Nn�R����[�W�#&aQ����A��<�B������ׯ6���ͮ��n.95��W3i&�8�����ֳfVz�7̚�����϶�����2��2U^>sǁ��{� +
��N%��=��i��Re����=����pj��ï���(+����d��n ��T��Z�;��I�tVi�3(Oz������K�fk�{e0�~+�T'�c�a�.�Vjk�$�
�Sn�U�iZ��wu�MX�$]�|}�[�߶QZ��2�ǘ��[�ν��z�<���ɂb���}RK�lu�3��K�ےǶ[ɿj�*˖'IG�����(�E�Z:�\�[ޑ��qu���,�o����C'$Z����9&�5����8��2�>AG�g�v���,C��;KZ)�"�{h�5����dM���ڧ{����GA���*�+�������x7#���T�M�-��
����l7���o�"�T��=Jv��(�7��t�#w�/]_4�1M�Eߎ�5�9?)�Ӹ~\�
G6�oeܑ$M��+��8s�2.�a���r^��������δ�y���EHv�u��U/�Sj퀟�A.���o�j��)��7�����xyE��}����B�i��z2���7���Y+ҕ��(�&�vƢd�h�������J&U�S�h�hO�@���j&Y�Qq��ɴS��1|I�k��*A`������d��@@	#�U�-T�D�Y��s�K�AY�2�4�x{J{�DqC�%j�Q�+B���¼��o��Ҷ��H�R�ւPFd*�a���?���i�mJ�O�s=�^&��(G�G*/�x�R����T���L��{�|�ς�R�8��$��@�}���D{���{�9���8M�^]�V�L����t�?Ki�������^�b��Ί��^�&���roz�Z�E�Ći9~���3�)�ÂK�g�M鲐�~�k�3��p�/lXD�x���"��*kC�^$��M�J�}f/���[]��1��vDa�R��Ky���s�C��)DC�O�<x��Ψ��	"R˫[E�A�\���(E�*��J��%"G.j �����2��2�iܡ�k�{wE	O�T�"O�$��:��K���{٩=��B��\�Cߠ&���4�$g���[s�Ĩz�/�mj�
��p_�%
.�lI�0a!+^_k�G�/d9�_�*|WS��K�X��ˆ��6h=�@��'�'�M��ˡ��lʟ�C&G伧���Ҙ�S��1�3R�P��H\[誯M�#���1��|����ɉ���Z��g�S;���d�&.� ���|���O���"s9���m��Ӝe@���c֯��$�rD�����6��{���AB�7J|	_+͵}�A�×>#��2�,����{_��=�e)����j�;=�X��5`�'kϒ�Jv�5�#�sֽ�Uvf�i�Ie���_-�K�d��a���	694�uZ�4�{RW�����}��=��\�����!_K%�6(�Nyc�E��P*��ӕ�R�����`2x:|,�=�4�>5ӓ!���x0l�s�d�)	�Kwp��e�
��4M][���h\�fW�K�S[и+����}�V�1d�F��8�{ ���&F�!��ĩ�0i����1�F�(�Nn�ɠy�����}�'Ô� ܈eqD}�vp��|�G'}�Ds��L	�^�\)�~�H�F�6�1����3տ�L�wU��'�>>�;���0@�F���u���x�>�Q\2��;}�5�A\`q@ƭ��T�s��5� �I�<!XU]�xbWE|GWF`���-������-�aJ�����\������>�,Ѻ��^^â�����4�<�͹(��\� ���J���Uh�D�iOz���m��=o|B��;��m��p��,U�tԍ�=��cEт%����3��,��� /Z3*��eW�A��]t�5՟2�	,�+=9���-�3����Q���g�D���y��s��Յ����	�>nI�6c�D��WQl,G�F��v�� Ń�@��I���4�!ʼ��-�T��3��HU�5�)n��2�ϡ)$�NK�A=�A~t+H$;HZO���#EYY�y�,�`��c>��N��${��n?ϑbu�Զ����6E��)ʐ#���c�t<T��P��L�Q���R�	G�%�ȶJ+6��]L�b��#��:��>���ʟz{���|�JN$��r�:@��8������)��)F���E�oQW����)��G���(u��ů�[�*�M},�Tkf�/ʔ�o����B�(���(5I$�)	��K�m�RWY?�ݢ�QH��U>ڽ��̱t��2����J �t��GŪ��Ag�.eBbJ���@�O�rA��r~��*����/
�K�"K��>��U�Q+���8ٖr����9�&�1twX��1�q��Ȇ^������_�=�>�<�]���E�錤�˲�W�H�P*��@�.���jz����<-��X����W���x� �0{��+��Z��N���+݊��5�!�3Ҡ����Ǳ���H�p��$mpޛz�&����S�Lz�+װu�!f�ڭ�ܧ�${����E����A�tU�(��˵����na��9ײ�UHާpo[-���
�#��� ��Z����)8; �:V�y.��~v)m�t�������� }�ݴJ������&��_:?
e�D����bf��ƅ��*#1���[i�e������rL�I��y��GP��֌5����Q���z�b.����A���6�
jn[��ׅ:(����:k��>�����eh�@1�$�;3V7�z�V�Ȫ�� ��A[;��㊀�H���K�Z��%��WWy3��(���#��F��T�����]_��G�QC��C!\�Y̍��tR�J@҅W�����O@һ�s]�� ��B���D#禹���L&G�d��Z����K+�:�=:�8���]���n�Jv��� ��z1��U�Xf]i`�ʳ�a��4L"nfNe*O���"������QxG�7HRj������x�Ǡu�����1�͏A�[��m� ԃ�W���'eh	�Z�Ń��]�Ŧp�y󽊉�ٮ�P���"� �����_;jԻ/JҒ����F�J֕�$HC97�<-A;Ql.ʈa�{�X�[\������U`�����ȁ$�� ���;��� �
I���vB�I,K1¤~��(dQL?&%o?%ߌ��f��.̂R�Ldr����!퇸h��Z�?y�ض�j�O{����*�㖥LB�,UE'�zj�^y]�6�5qR��l-x~ju�2e���L`P. !��mM4��mM�� I����&���W�*�����1��@������V����	T��g��Rh���xGD�1m��l �gZ����rP��A(1x�~T?����m2?T�����R:��zN����R]���k�pZ&��z*W;�Q�,?cʙ"�Q�H4h&� ��+�：h�Z�ScՖ飩����H^�N|�;�J@�H����s���@��`�в��ܥ�"<�?�D�٦��"=�d�g>�l��9P�l��*������u�q��&�$�u���<����s��ס���u"��X�!3XA)�
.>C�WYv��B������7敛��A��z-xЬ��T&�:��]a�v,lUU��Z*b�$�/�������q�
 �+�,��]�%#��2?P/�1r�X�	q�#�+S�!t�Y߅u�G��4bM�����_��-����[�I )�_,^E��4 p�D%���9�g:��M�q�A�uls�w$�V��f3{%���@��)�@�9]`�E�s��o�, �H\�2l�����S�Pj҆���n��?�P������- �k�Qg�1�~'Uί$@�����l�d?x�A9�鐱�����v�9��G����`m��$�L�ng�!]��K����Ns�Q�N��|'
&��u�IȂ/(�M�D��kt��冣+����1��|Ԇwt�0�${������k��ŧ��?EeD'����*�: �#�f_KA�2c	�R	b�;��j^J)Sw�װF�x(Md�N�T�p�(a�4��%`ӡV�D�Nl!P��~2G�m����QbJ��c�W��,R�;D�����EO�D�S��9���If<�����a��4���,m��X��s�2e����+?��8<�Nh]5K�t�.�V����@"�_>A�k�p�C��h4z�Z��^�nvv���1�&l\�y �NAWq�<�4xmZ�x�AɴH� 	l��v���
T{�4Ӻ�0�Xu/��E��'����eˏg�� Ww�xc:�^T/��h �[�lc��(�/��j�S�P��8�:���|�;Nv۟4�>�	<��(�*�$A��� �?�X�>Y���8Y�)ݜ?����@�%���oU��Xj���ue { +�C��.���)>�O�ɰ�v�b���,����]�g��b���g)ٵ=K��(}.Ǻ��#��`(( ��j�҄��R�2�p��%�5"K�+�	�x�>XP�Ƽ��N�Sl��M~���~4�R# 0�S^�+�X���y&���kI�D.�*k�T�A��H��+96h� ��L� ��MO��x;8�Kd�����u���ed���Y��$���B��4��хBYs����Ŭ��o�������"Ҧ�)��R"+S����#��?�;�AG<��*d��������I�+�����S�>h��4�D�ظݔ�̔��h<yh���'l�R�:4�2z��K�bWUy�K��{jё��鈢�	w �;U�ja���V���<����)
 �=�/ ��1Wa�.�2�LÑL��K��K5�<�Z��o����ɮ��6h!� nG0S�;u(�{1�Ǯ���0Z���F��ֿ�Q#�'�&�\�pPs���d<E�E�	�Ä���e)3����5��4��7�6�Y���F�e�Q!�BK$�Y��\�p��S��U�YP�=8uj�:#�]�bi>�#�&�7� ���%Km�Fh�4��C1H��WW����[��8��?b��M��4�C�-] <� =�O��w��T��i:�u�|\R����n��G���ͷ���G�JEP����($=F"�5�@����s��K�%y��0F�dZJ M_+�z������Gs�(s�ƵͻVC�{*V��32H�
B���wB�� %����T ���Np5��%K�$;W�A�q|���c��&R�A�5�����6=��ޚ�4�����
���g�z$lqq}��RJz�ƈ'����KVd�H�_�
�2�Q��0�A#|�|R���[s�#�e��Ė�6	�J�";y�v���:e��G��O:�*��Ӄ�/ ���y�հ2��]v�Ddc�È�b(6\6n�����T+i��N{����P�8�`и]j�_�0���i�I�%��� �-��[M�·�p)�r/�dYr	��!��JRcq��{e�$�l���$#/<4���&Ҥ�lu�ǠB�8�pguW�ؑ��#�)+#8,Ԃ���V��,���V�;��z���X�s�tY��X��V�'6�]�K�2�S��Ȁ2`�eג�&��Y�:	o�yD�y\��xE�r1��h�P�!2�jW��g�@��p��*�w��83>j"��>�T�ʎ����}QZlm� -��}2{�h%$�>�%�k1 =Virn�ٿ��HzN�r�����a��-@"e)�5��[�RV_f3_�W!zA���r�VBv;I�Mc��l5#��� <�E(EM8=�j���C��֔'�%.�W"j�؂����Q�_� �nBǩ�* ܦ���%< �<�-\e������v��g����P�#��^� C�L4��e�KyM��v���Mu�<b*�F�Ar�q���۝s'~�l�J�Ci<AAD�Ϭ���B�c�<ãsyB|���йۖ<���%��Ď"�;�4D_c��n�=��B00h���WQ7�Ƅ�#��痝�s�x�0-]�*g�k��'$	f���x�8Fp�{\��G���1ƃ� ܆�Z��e5�#�k�跑:�zdK�0%�U_t�XC3Ϡ���iÃ�t�A?����)�f;U��:��*�xr���Z����ϹE��q2�׌uD6u�\�S�zs�b�$H�~b����z��X^)�X�q�^ǰ�*˥��EC:#02���իb��r��'ak!�!2��T}��=�#�jD��)W���p���:��&+��k�(�\q��b,��$5�F�ݚ=��0;�
�	����\���)e)�m}D6s t͓�~c?�=f�;P��*.b�i����c�_  b�y����[��RUs�錤�@ďJ�k�4�o�����M�W�@�xЭ��>�y����)���w��x2Az�@@�4�p���	x�_�4.����
���,>e���˩π{�kސ���^xb�Z� ��H�Q�,����	�3<��RAш�@�#]�;���ҦA�3@�	�qD�>'ʓ�E?� ���Q�l� I0���Łκ����@tL�]���;�Y�H�T���Ɓ�PQ��q��K��/s>�I_t�_
�P>�� ���P|E�ɶ�<$�h1>����M��-��\�Ug��}���7�I�)���9:��>W\/>�sM-��tSܝH|�k�V_M#p�O;�t.dO˶����@��0������g;{��|��An
�'��O�D+�%<�{�3	�d�Z��qڱ������@)��]BJ���N��\&pr�#��׋jp�o�隣�tiP�� n��(E6��,{�=�Pk�H[<�S͕T�$D�OSb7?�O(�f���:�i,��T�x���W>H�8�x!@τ��V�7il�z��m����oP�${���"r4�&� �S�3čJ��Y��*{�آ�q�͵��rP�c-��tI�V�?����l�׆����a�4I�9�X�ǎ�4��%�0�.װ�<�aş�a1.��%�����U�U�lk�+m�ע��WRo7�[Vm,��Np}��(Nd�R���je�n�f��H�s���B�H��䅈�SU~�&�"}� ��a��rF�J�^��D�ׂ���Ds�����$	���-T�_�h�Vo
[�O��G�Dy����A(���%���H���\i�(~�$ju	��hV��H-,�o�+�6�Z�)79�:�:��?��n�NpZ +fcN���vS�����!���{�4����v��N��k�af�c�2�=�4N��zF�Sz�&^��ҫ'#s�!7}Qc��G�!�\��f��ҋl���X�-�v��SI�(h�?5���&N�� %�cؑt��P��=v��k�rD��T���(}�h��ʽ�]#�.gdW����/���3?�!���(����IX%����4y�lW��!���|;r͓!�&C���ܸ_ِ[�:|�����$��u�T*�E5T	R�  �
���&����}N���U+�q���M��2E�gⳤ�c� ���@|��q�h∙X��.��uSXQ<!8:I��Ndo!�+u����zU�r�~h�f����1�m&O�-\������(��Z}U[:�0_��٠���X���n-D�awh[�,�� ��Al�DA��N�N������ �^�"�2�[�:h�E��	��j���W���[�(HQ�M���&ac���U/�����1.�K��Dg�д���mBث.�7�RD��&������1JRo�5�>:9�;�!��˼�0�f���Gg$��B�@ �t��X�J�j6�TG�0�@�$}�8�`�2;n�幟�K�q�e��6�'b���n�ѡk� �j.,\��꘱��^@z��}�@��mcT�Nϴ��#��]�J㋲P[�Ӆ�ې��ɏ��*��x��w����J�C)d�������%i�X����s��B���uu��$ �nN;,���},����.���uS�v��tf-%�4|$z}`e���\���3[g�������@��0H�[)�h/� ��O*O���5������o�xv~��R�"g0�;M�B4�Iɫ) ��D.�S�QⰄ�Cu�h)__����\�Hͫ"��R����,�牞JGc�fxjV�gk�ż��~/�C�&ąH�#%���8�s(��٦�*��q���ȑ�O�l���A�4����C���\`/H�C�H4"FpeV�Z�w�ڡ����c��;��e��c�V�tiAY��^��k��D����q�������l�ߦ�m�s,��AZ�W�: f|"�XH:4�n��GTO���� A��q�����VѺ�P")��$�<�f���4��Rn���~;���spd����Jr���G�2!傘S��VR9"o�:�"�^�%K`��
0"�Y��ϭ��R�\�r�"�����1�%�) j]�o�uGģ�\��
�(p���Kj�� ,B;�!�U�?,�$��$K��U�AD�ҡ���wA�K�	�>�H��z�$ʢ@y����1�/�)R��?&_q&�5�w��<�P7�S��޸)g!XpN�^���B���!�z�����g�&�e� BE�9�a�AA΃W��	Vy�4ӽ�Kc@T�.D�Zr$�+Eݠ�� I�O�89c�*;ȸɚ���c@��tF13i�����p5�Ȍm{�jc���������Eܨɡ�@S�Ԡ���s0�ө<0{��R�闎���+�/^l�����[��$�WK�8��ɖ���X.V��м��_M�N�{�50!��\�՗R�a�g�|?j�{�L�=��c�WyD�M?�O�l7	�/�LSWcW�{-)p���Xw�A��n�~"�8Ӛg1�.��s�+�鮋(����̜#�<�>�D���,���d�;�'�ȧ��&l�U���f{6(���͜��W�:��S�g��=B�5mj`3�8���0`�)!@4"�ȵ���W�b�c{��#���42ҷ���jopDV9��6�
����bR��,#���+3���W��<�YsŖ�5y���g���E�E�	Y�����/�e^�I$p'm���}55�․9��ɨ���,cL�$,�B�DʀJ��x׋E��gr�/���8`����Cu2%�b���E�FeMs
��pK]�L
R��(�CP����)��,h��LQ�|����H�`�ŚZd��<B�1�\�����:U�Ð�ְ�rD(���Y����Ş����n�Ŧ2�[���
����&FD��v�5�o���{�*e��xȯo�_т�ߎ�di���U�=�!�Ե�Ҡ5e��?�j�Ho�9B@cJī(�(����9��眞m��H�׆*L���2F��Xy� +?�h�zv2�h� ��D�p2lrRC}A�I`)�0�L�I��`
��ixнA
�m+c��K�`�v���2t��X�݄�����[1��!'A��`	��KR��`�<���h����z����?�!��a��s����_����O��-^Eia��jD�����E=d���W��[
L���O���/�`u���rDu�u��:D��b���\�(� ?��D#d;<{�ǯj^��<�s��G��S\�o.J����A��~������K��Nm$!ngnq7� G���!qL��}.dMŷn������`8"
�g�_1�ȥ�d+��G��t+?-~��P�-�{�*�f�?ۖ�"���KL��p�;����B�|UYz�_ϔ"'[t��$0"0�je.�o����1��z������$ȐK�(g���nd�5=2���Gۆ�U�Ț�Q�;��>Fh��WF��J�7ur�	�r0H&�8�e��p��/��1Gs�X�s�z?��9I�ʲǝ.��f�(*I�����W�QE�U��kׇׅ�)�=d�!0���*�LE'��DHYO(��������r��� k�z�����?���.JwN�������_�=;��{>5��6��6��rV�b;�5�d9��׹���?N����\ı��`��;�a	"�~7J��.�:��Ǳv��y�1,X]�K[���.G�`Ս�v)�9�j�zOk��a�uk��t
����T�0}@0n{:�3��3�/a�C�-Q������!�D��W6�҆I{�kc򿭵6�s0��+��
T�_�B[�2O��k�A
�h��T�)/�|�@	pn����G��E���$��<�v	]��7][.����Gǅ"^C���>��B�P7���n����"�F�,U�	���1�%Գ�	;������6اO���Pl��V��؇�}\����3����Əg��Nذ�ʾR[19��PAl�T�5�]H/���l���I�	"��m��0���<�H_Mcu�Ra0a��w��!���4J��|!�w���mt�Kw2m"��]��+�
�|���ڠ]ev��i��MBa���+��+Nl���5e~��zy�'e�.�d8�a�@B���=������͏�
E�B��i��H2S��6�����Kf��2�v��� �n0���!,���]��%�����w�QM]�Kk�E�S�����.��ThE���Z�j[�S�j�}�� �@�+-Lˌ�EA��
*�G	撤@�"`�@ 	A@���%��ܛ�!%�>;o����R���޿�����ۯA�A�j�fB��W���c<��|nQލ��tW3ߤ��u|���)��oH��q�}p=ŚO(E���$�"(�IwE�ƻ4��,��ɓ~[b{h�P���C�U��;<;��-�
�D=��L�T��#8����[y�b-�sgK�-��!�H������=�s5_�ȸ��N�-=�Ʃ�$�����1��W�Vo��q��]�)1�M�8-����gp#��(������?Ŗ�?qr��J������5�[b]\�=g�b?6i,�ŊJ�4�^@x�LT7b��{�/x>��:]����O���wώ+�p�2m�ez�| ��"��SC�5=6�R\�x�߭�AA,�Ɯh4%`\�ɯ�e���!l��F��,�ǁNT��P�l�<QQ�N�xOOqͷ	�2�1�y������~�7Se�U�(�.�Oj4��O���k�������Z���s8H�?ڠ���0�3]�㞾��1�VAl�W�/#7��	X(���+N|cX�hǲH��}����'�5� lX�X���/c�V�Z��Zh����bl�[}j�1 ?-��ll���."�"1��E�������W�w>������
�%{�[���-jQ�-�kH/�c1�P	���⃳]�wI��0��M��#�e����ԙ�2�4��c64�g��S|N� �v�������x�ؙ�o*�~��ζ��0�����UT�Kβ�ǈ�B>���=Pg��eUʽȰe��D���zI��E�6�{� �3��U��Y{���<���l�S�^t�������Q����w�Հ�`����U��fuIXXpC�V�<oי0J�Jg$�D�S�������>�*�HL *��L{]?.JD[��66������L1�:q���"�N�ؾ���o�`��q�bfv��8+|\9¢��liآ�: 1�r��m��,���7���N�;(S���/ �9�4�y�5c�Jb~K��G�Zl��65���������I��K,�WmP���$���m�*[���*?U�i��~����Q��P��7s����:� eЌs���Ivb����}!����.�`�H&�=�Yl�,
9o��z��sXQ�ļ����s����zCq#�P��ͥ/U��K�����#c�����bg�0Z@J�ڪp�1��J�ed�5b�?KJ|��JP,_N���kc�b�w�%�h���I�~J�;�Q��`�%�"4@�=���3���U���%��AbW����i�N��m �R*���G�@�)|�������,P\q@���O�a#�So���J�(Ǝ�&J����i �����w�#A��$\�8���P�gٶm�Pܢ��u8.�����+�e.m\�����;���'n�`�f����F�\�]��[=��u`C!�)� � ��"�z{T �PR\`��Hθ]��c��C? ���T�)v������bӟ�.��2�2bE�7\�ZKH�aQ��)��U�v1�����h�/��_��?��Ȑ�����H$ୢ�dA'�������^2?��A
�
$�R��k`�j��q��* ��wUp�� 6�����X!�5\�2�f���S����	|��=�!�Ea��^\X���� {�>�^����2�G��!��`��}Ğ�ոr���%E�av��ު t|���^$��r��c~1�J�[�o��.�	��5�./��#���h�e �{B�-i��F���5\�<1&�G�p��t1�P�o�ܗ��H��J&��5�n�Ў�&4*�Cܞ�rԝ3X@�|]��vS��?σ�ӟ'���K�N�j�'���'18i�m��ӝE��W,y�G�3�P����T0Fc�O|�mG�Б`&j��'d.������ӆ�
;6�߽�i�:|U_Y�x3����Q��4�b���Ad���WiT��p'=g�]z��=�����b�#?:9C��G�G�\T���*"2����Q�y��y�Zş�ԧ)�K�\X���5��L�S��c���9�bu�MI���N��CI�{~R]��{�d3�3>�\�D���V����H����x���$*׹Y�]���u��G����=.�l� ���,n�">'�<lӔJf�������r��1��MW��].44��NN���S��k�e�{%T�j_f-0�X���0����ʄ����z�X���P���t��e1�X��+�A;W4�̖��.�����������R���7����ۅ����~І?��q�Г��s"Ȕ��7��*:��7���WV�d���.��E�<�_�������_�roffERi�W�OT���O��J{���T��%I�Q#�%<��V�o�W�n�\�8l܆_�'�V|���_l-�� ө���;�*��S�C�)�'-i���ڔdB΍�*�{��QXBo���--����ܫ5�@>����l������S��PGJ�j��_�O�+O�9�a9���"$߼M ����2;ZIo��2�D�"����)2U�9�q�n%Y��Z����
:�r�[ĵX=�����'^���d�9%޻JﺶV~�����E�st��u���=I�O�:Qj��'�ȍH���O����e����C�����X9e#2�XZ�|W��g����KS�P@7����飝��Y�-��`Ϧ��(��X�||�ⓕ��\���������y$�����s�T�mʞf��G"�a��]걿4z����A��e#��/�wo�<���\�1�	������b/�P*^��>�����wA �*��;�SG�o�N��CS�d��7����\�Z�� /���`����\���sfJbE@��ܑ�r�*��~�I����X���L3���M ���օ�'ُ����Q�Pt��	H��ԇ�����%�Z�%��tn��2|�;k7Zſl��3��D���[o,{�5Ms���h=v써r�m��s[�O)1�/g�Mb��c0�~��+�� r�<�9�v\���� ��7'1�F&R��.i�ZV���/m�:�p�D �9=�g�� iG� �C,_����N�3h<5;��i�V�g��&�.���u���G�w)�<�Zayv��z��,�G��ݗ��>�H�7�	�g�"�nca�W �oc7B��N{ˢ�׀����m>W���I|4[���]�9���y�����y�chxn���َ���@π��O��]H��]�]%u��-�g����[P�|�>��$z4*D���5��Ly�!�`���"MR'�=�%6��)��0��K������I�5�Gñ<X��� ��Vo�B�����V��Ҳ|l��N)�����>=W�vu/��l�����o�\|Ay�p���̄B��@�xz�w�ݵH�Y�35E�K:�|y𕁜׉�'Z7	p��v�M������+�����x�{A�&��L[኎��<�	ƻ��dq͈��X�S"�?�:��(�|�_}�x��R��,̲�=�׽��@�%� T��Q6"}���IEF�'4�g����)+�(��4����F�w����!���y�S�Q�g`�k��Q�{-A�l�B Z�Y�_1(�ݮ�Ҍ�� �>6��ᅊ �����-����SL<־Ḩ�~-۞=Q�9Nd��n��3oFN�i���Ybl�t���u%8���8�e���a�ϴ���3к-��{��A7�zG��x:$��gZ��vdٶه^ז�-�呭�(Z�aWi&����W��a�:`���?MPߙ�0��t��9h�d���h�Ry�;�"�BN���s4��F�i��b9�%?W|��M/J����IFk�a�!t��[b����/&ڲh�{�����}��XU�!�߂���y���R��7��s�m+A�cT��m���WL���ż�ʃ^�$Ḿdն
�u��B�_�@�t�3�<�d�]�sޭ=���I��7f�m� >��y�E�x[��4JK~3}̂���0^o<^�����St�3s*����.�����f�ōܙP$ڣ��D@��V{M���ȯ��t��b���2ɹ��@Tl�z�9l��Ķ�v�#�̥�#rw;���`�Y���:s�l�s.�RU&��>����	%��$j
�ۥm��b}v>��+�-�{Ԗ�*|:؜)v��.Zu�/��b��kc#��N*��/♱��_)��N_�� ���&����칅�A�V�m#n�l�P�Z��Q����eb�Mi�5��Y�N�=ei�/�����}�2cಝ��}�cSrݤ.��i�,�*Ev-�=�����Cܿ��2����4Li}ωhڿ��a҈��52stО�W����R]�H<�����&	jY݈R��Bn��[+��(�f���x�n�7���U��sǾ�?�}��ϱ>�>��PmE���n�)����)@B�.�vJ�6CҢգ1h�b[ͲIE'�BGWG��r9�z����$i�Sc�"|Mi���kN�0���Z�\w��4rNN��mG�T��T���Z�^A���bPY"�Idt%2F���c���H�T+�����ШF�hhXHA��� �Jjn��I�&����.���ϐ����LL����t���WǸ,tD�Q�þ$�%�Ԓ?�mȨ�=��4e.���0�,���W�>��
=�#)|gmK�r�ɖӥ���a�B�&� �<Tǿ��(�sGh�P��WtŔ�JZU)j���H��/��ۡCI#5y̜D�X5� ^k��R��g�\`]�=J�=W�:W�.���8�6�EG#���7D2|���������>9w�����'��ߥ�v(�?����\�W��خ�L���6�+җ���52kd�Ȭ�Y#�F�_9��S]��|����������������GW���9퇈����&�BK[��~�bnm�õ7W���˻uq��8	���t�z�����)�;/��w��{��z�.583k`����Y�f��50k�?m�� ��;~tq�C̓P�+7�Ĥy.fҶzQS6��[��&w[Tul��$֍7���*{��dnuT+0�㎷�<yܕG���s��~-,v��	�goy04����������!ǎ�+�mbҾs��|�f����*���uu�Ĺ&&c+�_��}��H����Q��ê�AW~��1P嘲$�00�.i��q�V�Є�-r}Ш������奻�!��9\��h4���p8�N[�4<N:��pG�=S*hѭ�y
�jA�.4�* �J-���Zm��<"�!�9lN�Rt������ܘ5�l�*�ۏ
��PM��	�κ��	4��u������ޯ��Β[�d3���6{m�ywߩ�PK   ��X��x  7�  /   images/865a90cd-818d-4d70-9e9e-0a073e8e8390.pngL[TT]�>C�� �� ]����
R��t+����R�!#��JH�H��CJ��0���/�k���g�}v>ϹwB55��()  T*�
� ��?Br�N��a�����)z`���Bs�. 0���]��	�d权�����E��Hv��d4�M!���p�w��)�C�������iE����r������2_�|�T3����=�I\�����,-C.��y�
��I�Ck�+��I�.�^J���+)-Uo7���+�^�`]�^��=K$����o���eK�9ߴ/�K�b]΃>�v5F��Ku��dk��Wk*}	2�[>����HI�NǮd�z��鹇��N�TܿA��*tGG��]w�j�w��C�p�B��Ua�d��M�,�����U$.ُ����냐��Ҍ}n@j���,<�9)s�Λ�t�y�n4�sv�V�-�菥�9�����}s6��z�J\�Z���X���e��e7[OM��d��/���xb�և�4��_״�$�<��s��^�0�T���{��8/h����2�ICE�v�Kkkk���Z��mï�9�v�?M�9��gW����*�����R4.�gK�4d�VY����
L����,J�A�W�x%'zg�~}q�������B{M|l���wr�$�?��2�}�EǊ ��M�'�N��22?]Ck�M%F_G/�������1��`�J�����rZ�9@_MǄ��H�g��P��	HY��dJ��n�O@u�J�7jy�$j��דc&�(�]�����@F����e~��u�ظ�fa8���.e��Hc��.ݓ�O�S��7��kW���z�������l�"��%�Z��g+�V�>[`��2�	U����nq�YoK;{�A+eR����ԝ�����yD�t��"�֊�J��{�����`�UR�5_҉���l���{��Nw��/^]���V|ǰ��o�}3x<��@&�e|Lv�yes~ЎR͆����'�b?�f���;U��?�[S��7=!ltm`���e����=�X�������.��T�����(j>' ��j�$m�W�8�sz�d��4*�&��UٷV}�������}�=F����+������e\���<�9Kc��19��[�_�~v�m��(p/.`{[���u�.^�J�,B���(�o�kGu]1���'P0����NXX�"�q����f� po���A�#><ͯ7YB���̒�׺��U�Ȥ<�[#����$LQ�z�?�B�z�Z-�mIq�C�{�����@�C�K�N����c�$��r����3�"�b0�z��r��q����i���;~循e�ګ�t��T�j�;��J�+&Ne�P�`�W���H'������5(y|�nU�j�2�C�&/��%~x�`�!��1H�����]��>��t]�Ȗ�ϔ�_=��K���X�_�]=�� K옇��=��	�{��MZ�]��̢Tl���)'�{ڏ�A�vm�*���"�2��\~)!����2-ղp�����繀�q�%��˧����T����%���M�N|A��Jap+ъ	�ܿ�c������Y�����N&���IK^�O��\E�7������cϜ�?�S]l�(�;���m~k��Q�g>9KN��̃ؙ�.�����r-�J"S�}����X'�o�����k4�VK��	��v7"_���y0�_#"K��Ɋ%�Xvȿ
2�ebe~$��!�j���ɜ������M<����󼛎K�rѸ�]4�'�,n�f���t-�jH�����W�+�=���E�'�j�j�%�m�6sڎ.���)WRvm�0���Sk��"���C>{ǃ�^<H���_z�_-�9�5ا?�Z1��mE��m��b��e㜲�ʚ��_��~�3+�
|��Gq"0����/K�$��u���yU�5\�Vq�e>&"�˼l3z�*A�З�=��TL�p5�ӎ�`ձ���|63��i��k�B!5߬ �! ����	�.z�4��y�1[�����l(�@Y�}̓��ݛ�Vn�.&�Q���ޫ�W��Z��*�jO��<.���,������?����k3f�n
a��	T�P�Q|)�Cs�6�����g+��/딤DF�1�e���2�P�1j�[Pq�^���V��3��2�~{0�G'#bj��3Ry��
��vfN��8Fy�^���C$C!!��m$�eN�~ֈ��j�=970�Dʶ�n��X�?T��D5�O���@c��iF�)���t'����K��Y�w�"�1�^FJuO"U����zЍ�}%�����ת?�G�߉GH[�-���^���T���,>�b�q������*��k?��3�1p�S�,w�jU�ں�Ǡ~?!������!���G��f�t\)vǧ٧�m��xoo��@�޽�?5���~[҄Zv�-�OA`�l��乣oc�Ҧvxp[���AA�Z�z�g���{)l� �`)i��k�#ڡ��j,|�����,K�
tok@|g�m.>�w�lXH�ۣӞ
<��4��Ы���V��d[U�5��w\I'ؤ~K9��i�?��~�h�K@N|z�{�D���1~�pеI�-Z���r���p��4(�x��WX��1�m#���+�%x5��4��f��??�b	�E\�M'(���l�+ߨ:����2&����fG�,F%i��|�Jg8s�^�v�p8> cϼ�e)��8����.��Ztz��R��3��-��bj��ns��,�E�3/�7��	�G�R�S��g�rO&B>Ӂa��TC��U[�%��5�B��A���o��������J7o�nU|ԦSγE�L躜M��-����b�·��<��H�C�Ć��jx��g�ۯZ�܌>�'ݎNL�K�)������}A�{��AKn��+0��s0�_�~���n%��)�}4?��������X�4H_�/��qq.Z��Č^+Q��{�߹���g�Ӏ����7f}�Aǅ.E�<<Y�s>H���)�٨ӡ��ܫYJ�ڠV�mXL��3#yM7�@�Mc'�#�90����5�t5�w��촠4߫��N���w ..���m|;u��2���;;*g�Q�I�B}{tկE=^���`�V���\+#d�ԹAk�� (���9O Rf�
})E����ׁ�O>��Ojz[
�4k��Nf���wB���>kO;?��[>����)�����
���CgP��7$������ܑ���Ǐ#ҥ��r�ﳴ�.M[�������;_���u��	��z�=���3�y��c��'k��{�LzO4�C���l���ôpĺh>~����=�V���@�y.�~��%(�wVa�̏�;8&FF#��K��"�w��!϶}$,�@������{���}�Ị�N���0r�N�
$���->T������5fW8��t�#�(7�.�h~K-S*9�,���w�MC��`Tjo4δt�>��mK'�\��z��67�u�$~f���|[�#e��Gm*	,<g�JP@^4a%-��������j5���v��IW''�Bj7A�춴�+�Xs'�/�GpTabR���g�b'x�I��=9�FJy�g�L�������MSqnA�i �>3�x�i�J��]������<��!��c��xa�3����f �V�A���Ì�7p��7�4*<���g�{1���:̸+ᦒL���`�Ơ����Q�1�K�D��"�Z3E	���Az��hs���LY�--��HZ�^��ocn��FGhBҬ���e�r�&�;��kN��:�C���s;�_����������E&l_-۸��gy���
5F��Q��)"`G�߿�^��HϞ�u[&��?������D���8���9$��WZ�ə�{�Â[���Qj~XG���W�*K�o_ ^��	�TE����5�O�|�a�������Fڃ�s&����or�Mr��	���3�cm{_8�W4�����%ܤ���>>\�����ĞNGJ�sq��.	�бO:Q�&{��j>[Q��`�Y$��1�h+�U���<�������<Rq_��6��b�QE�%�Ij�s�<G��\�)�B-�Հw�������q��pk<��>c�b��5R�l�
*x�L3���-/�f�M1��3Һ4�v e������݁�hIi��U-*�͒�D������9@O�ૣ�*H�=��_�h����F�ֱnN��������$b������_����A�J;���� ���k����>S�rZ`К^T���e`��]:�_�S+��0���`���]|>�}8w�JO0����5|6��5���er��f�������c+�azm♸|=Ma�"�lMhs�e[���x�;n��a����%�S����B�~z�Ak�����x�\���W� ����/$+���ˉ%�m���"���0��8����N��������õ��6����1tvZ�<�L�V1�Ph��O	%<\X}�?I�}����n�rG3خ��e�̅A�Fv�|��]{�hU�ā�H$��9�Q�.��u��<�����[m�ᐊ��/lz�����.��x��\��H��ƈ��}ɽ/�_[qR�iR����9\)�D��Fin���IL�V��,�e���T���V��]��2�K
J���u����m��`��=!�{g�k����^!<ZȖ����U<�j��d2p+<���պj�f=�v����7�n�=��V`�K��UQ�9#=H��T��+x����6J�����=֝N���#~�{���_������av��{b�LYrH,��R!g?��3����t��{e��s�z堿%�U�C3�~ +z��$��ů�����9�|ӎ����Ҋ��iQ��3�ފ�P���M1­	ګV"�ڟYF#�k_U�~��p�������(�9lc��	h�-�,=��m� [�]Y-U�m���nm�bi��lt)T��ܙ���S���{�C��o
B�Y#gE���3zj���KMф�fo����vz��܍�r�I 6{k������ }˩��<��dHȀD^�����ӂ�Bs��F�N�+�����Sg4	x��y�`���������-^��������Y�_���:��Z���,{�L!{ޯR.��w��G�٥>n�'�Q?�(���z��V@'��Ʒ<�% ���P0x�܌�z�V��ǉ�u���
�Ζ�}�1Ƿ�)��C*em��a��U;��8�G������K1`I�ǋ8:v�'��T-�x��� �54�_�	
1����~�:�m���7���O����;|�`XSE���N{=�eS�J�e��3�۞�d��x?�������b���%g�R��7,�&���{�9��h4yϲ+Y�l�a����\7c|��9�2P�B4�qs�9��7��Ìwj��Аw3��_?�\wđ��E���{Z��CN�9
�� �2
�i;�F�Q}O�;Y�NSU�`d��*$���+��f<�*ॢ�~{ڡ��'ܳ��M��?R���� /az�!��}�f̙�~iW5**
S겓��}%�fo�D���l�9�W�N��&q��ɯBg���8p���S��/�S��#����T�j���ZE
��a�f���Hc�-���ˊk��j7m) Ʉ�yy�fP��(��􀌓0=��X?��JQ=��	T�?�}Cͤ����2�^��\�	T1vB�v���p43�Ia3q�qf�?�plt����������w|�3q��=�a�S�ptu���]��ʺM���g������������ (�d�B8Y���??`>��wM_WU�{2���2n���7��w�~��j:J���q�;Kش��w׿�S#"����g}3��j��wR#�#h��X�މ�1B)GPC�G.G���A�[y�}���� q�=o�f���P�+�J�خ���Ɩ�L.Fz#S��蒒�ڣ�{S�������9�
�%�TYޯ��~���ʾt�rcW���2[�5�Ve|�-h*�o��w��^�݋\��Hg�s*��]D=�/R>cM$_����rŬ����t��?B����=�ӳ��.����$o�Ax�� ̵':R@��m��wށ�P�g��W�ĵ��M��+7_Z7�zꔙ\g��<Z
�_SmI_z)[䎈�^��{�r6��֧�f>:�N�+e������+1K�6�������ɭ�
ٷF��w�=�I+�fz��X�2��vO��x�"%FtrѼ@�5�.h�����׎+L����z�	�M�c}�XR����_
���1ߌ3�h#�S�a�!f���OQQa�.����iF}(��YDWo>GG7y�\�?6�ͭqr~�ǿ��@򳹄8u��H�������>XRsQ,J�:�ފ�<���^�����g
�#����F�ō殢C��*���7BD�tx�H�E�H)�h�3HgpG��t�oY|����/��1&a��FO"�N�Lc�X�:ڲ��C<�;A�}��B�MO͂6K��2v"(A$a��Z�yA��pT��팿a%�?Q?�G��jw"ܧ�c�٫8���;����IZ����l��s2
F[WM �7_�A��Ɯ(�g*���;y�(��s�6M�J���u�=6� Y��?�A������#�{Y�3c�޻�ƣ�����(�%��q��O�Lt����٬�<>QA���h�Z��y� ����&�ʎ�\� +횿�}�%��kj�^K|_����,�y�Qӗ��E)���o�&I�ow��.Y�1'��}#gqUB��E|��5���i�:��h7#}$cZ�f��~���18�( @w�G�'Y�TT85�C; K��O���0FЩ0Ȗ�j�^@*w�4���\�;�1�{Ł�֧:r�SU��ӧ�IUU3�-r���L��u|O��	l&ߑ$"�=�4b�:�.-�enO`��N٦,b�f*���r-�OU�g<��VҦ�o���t�Ώ�\,�,��~=@
:;o�Ο ۰�؃��X1����xA"���z���K��z�J��:�9䳈�,��Q�:���,D��9�r �f�S9�{�~�ZBv��i8�/㶡���|f��8йp�!fK=�N|�D���L���SO�ԭ��EXd�N�S��Ѯ���ᯙ4y����;�d���
^�nV��e�[���_����JGk��S�@�3���ۼ�aRP6'����z=�:K۵������Ne_��@ע(D�x���Bx�qaaE%Go@����������a��v�wYJze�E����ּ׋�����.�~���|���y�7���tzR��{;��ϲ�!}���~̆0�*is�S<^����S�v���U�:4G�q��|�Q��,H�c�Q�E��>G�#Г)6^��['��:	ٙ�嚚��S���q�<�͞ξ=������/?B"5���>����4���x�]I�(�!����<��|��#�����_�WWR#e�5X�P��vC�:��O��}NJ�u��qtW����F�#\H�An�ML5>����S�.c�O/���vg����ͭ����~�a�z�m�H�W?1쩨E�>?ɔ�x(���3�h��)��~�g,,��6:����]�D�,_!=�he@�n'N�m:(Y �e,�l�83���U"}�K�_,���ER�s����%g�d��h����x����M'���%5ciF��t�WYhs���VU	#����q���o��+����	�2�v���dh�R���\v��?z̛�a�ezǷM�Q2������O��+�!=�JQ���-߂[+��#���~�·+7�{���c��#���U�knOF)"���n~� �W-<����[�G�{�V����i�ؿ�1�c�ʣOx����J�<1��Y6��a��5�Ν��2��L��1ik8��d�KNi
��T���U�n;����E\p�~3l���q,`;F�VӾ�,M�Y\�D!�Ş�GO��ir]X�0QμvA��+/�a-�]���4c�ӥU���Nep�p�������W'�	��Q�5���b�*��'�e��\��������ؓKw>�wH��1DM�b���z����=��awۊ��G�������X籛��s$�Cqt	�p��'f��{A�T�3Kf��a��%u�����Ȃ.�w.���_|����S$`��Qm����5Is\I��0�����ȷ�$e�`�������>� �6�É�|S�7l|�ӓ7��a�2���Ca�4aVJ��Ķm�p�����"�����V1�됗m*��_�KO�ڔ��aJɴ�E�5��ケS*�
O�:vMг�V�}����X-.��=���N�*sd��u�	��j@�- 1/����͝.�W���fP�{ԩb�Z��7��j:T{� ���ڈ�Bb?;7�FC������<�l�z�I��h5W$�HY�,�������?jQ�����d�#<����=��* R_>�f�e<��YM���2��������u���	���mw~H�Ľs������~_�՝��fZG�W�۠_���YR�/9�﹩�R�4Rv��Ε;�#bb�Y�9#-�K���|����o���c�j�zk��ͽ��^��QV�=yz�;k�ӳ�(hĄ��d~^Q����c؏R��8���/D���el�<�5+�s9���ɸ�[�������j��Cq��r���0t�gf~s�~4^v��i[�-5���q�>rJ�Sr#��t��$[�HG�7����[�"�Դ<�)��0���W����}�]Q����SwE�b���ʇa���y���	۪7��
���������^Z��ؼZ�')�!ŭ��k�
$ņ�o�)�}uU�*�/�K�܁|^M5M`����k�G�\ozC�v��"m뙽�f�	bߡX�2p���#�*�i���?MR��;*;ZU='�g|�SIX�B�Svs�q�K�ʋ)�CJ�%yXyd��6-+w�K>/�}+Q*����67?j 	=P���:n]Z�J��qU�K:Wa��ǭDL�.7.�JNL�no���$���E&D�~Bv�����l��9��������h���w{����,g�t�v�?�M�f�J�m�;�^#`Y��JF��8Ѯ����uڜ���LZ���s}�d�x���g{y���,H�$s}D���h�N�vu���uE-����`�U﨣� �o>,Z��3��ś��_�G]�)�ݼ}w)oј�͜p2�Yd1��_[�Ug�w�Ϋ���m!�%T�U�4��rG�Y3y.���&�*=�?���/�ޟ�>�XՍ���A�ig��i߂"�f��������k��Oʊ2@d�4!|�Ahn	G��7 U𛏶:bNnF����������ȝ"M��b OF�K�X��F�aR|y��6��V�Е ��A9��UX�<��u{ט����ߎ��bf�Έ��a���2����BZ�~r*'����4�\ħ������00}&����h��w���Ơ���o�4}�:�`U��N���K!��ZG�x����ˍ���ě
��|)ߵ�Qz��3tǨĸ�?y��'�;�x]z�'�ȟ�:���ᗌ {Jx[4���X2?>���X�Q���og'��b�&��Tے����E͏�S�I`�q�Y�W�?z-)����a��)q,\����������d������M
���A����A��Y�0L�J�����O�u/�{�::@ͩ��l�`v�F����EǍ��/'�k��tw�7(2'�h���|���Þ S�#Ğ�߳�z�%�1��1ۅ�k������b��m�����*�>��R��X�6r��qr��bbՌ���H�I FE��JԛzdoKc����T;���l���.�{V�)̯B)i���6�fӎծ��R�� �jsq�'��C�b�z���_O�ᢽ�jvѓ���`8wɉte?����l|�UX��B�����y����&��N��Z��}���UQ���l�ˤ",mӕ�����ZQ"�\�e��ܟ��G�Y�l��������'%ؕ��]	���e.v]fujU�>�Z�74lm�
�l��S벦L8�6j@�B�*�~T~-�5��9t���W1��a�'bJZ�$��{�;���E�E��94�i�0������g��t��C9��n�\�:)�rS�9B �QEH<B8nV(WW���Կ��~{Q��Y�:�F����ѕ���%l����1���!�M�2;�3$2��.<-��U���	\#?!+:�0���&���.%�F^�e�����C��Ԓ[K\Ic?n�W�$��|�x.Ϟ"[H|��զ�@U���a~[W74�5�@jU��W�_� a�W�ly�"�-�%�z���9��M�R�|r7��*ܳ[
0�I��5ƃ\���S'$��F?�deU�"��U��c��Y�|t�x�v]�Ǔ��6�s�]"�o�U�\�Lcd�����*6�QB82�q�$�u6k{v��:D�� �+���'u�ҡ�<�t~�,�C6.�ŧ�s�#'����z>I�z�&��L ���/G�x�E�{ܜl���#t��'Z����EВ��fK���o��O��$���#�Ç��D5�^�ǿ����&<�۳,�x�jxi��K03��]�U��QU�DN^���Q>LT�8w���v$�$\֘_��q�Q�����k����HӬ�L�؝�>����%ʚu^�J�߅P�A}���z�~�Gy鄆�cJ}�K����.H�Q���Mu)M��o�I@�YG����&wQ^����>�3�"du���.	~>y���	�X�
��7D�焝�D7���HF�E]]]˞B�&�巒*JDcS�&,A�cÒ�Ru��%X·z�aoCuI`˵9�R�<4��K`We�E&ѣ�:���`de��O�$�q�;ps��jz�OB�_���~��b��w�Z����P>�%���~q~#�0/�^z�)W��a��u�r͟#�E�� ��lV��%�u�W{�н�P���{P��&�\^�s߭6��+��C��U�n��ߞ�>���= ������i�.,&�
89S
�F<�����;�Ki��]�{���]q��閤7+�+��pY��9v�>���I�|�n�!��}6�1ߜO*o�;�a���ȍ����֝?h߳���������Cj�'N�&���[k0�R�A`|�����o6� �p��Ғ���֛/����^l8&����$NQ�s��SH۹��y��~�M%gܸ[7�%w�-1����f���	q���+���[����
��4�6eޓt��	\�=��qU�
Ƈ��2�,��8����g3r���!�L�G�7ا��e�`i=ԝ̇��B��o�|L}f�(������^�����/�~Ҥ�;���)B2:��&)�9�`o�u�;���ihr�Lú9��#�m�{ɼ�#i���
��o|�/�Q���а�Q�*� )�I{��*0���R?�]g-x�
��^�fm2�~2,��,��;=TO��S�`裩���`l�@�1�ec�l��diL8�W�;������m5�.H��Zw��PϤ���S�T�~�!X������jWZ)Rl�k4�
�zI��J�����_:�i��  �m��j]�h/���^Db:�VjJƮ�z��pe�� l\��d�Т�ݛj�/hL<Y�ƴ=�&3Eb��!����ǧ�6�p�˙���^9��2� {8��'��,�y��
����&���������̈́�X�S���;�4+�*�����Q�|��B��]�"揦�P&�Z��B�Ý=����囑�u�x�6�r7�	��sxpKm�1��ml��˳���J�R�;��+�6w��l�tp���x�M`�%�[�%���
�K���͟	��oO��\���;�w�����?��b'Q��j��S��O��Ć�a/�R�ӶKu/[|���,�Sg��}�����+#����$'�ߙ�U��g蘕�9�=����5iT��w�rZR"-iF�1�ï��d�kѯW|�Pݕ��ɺI�NsDc��F���y���+����{��d�ܮK'�E�;�;��aG?<����e	�K{�#Q���r�#fr�]��?`��=����~���
Ԅ���a��O��}b`?<��Al���[�������5q�.�Ki\[����C��	G�+�h��vP �V�Kώ�C�u��}�K��]M|�Dd]���}`@�T����-{ub�a�B��.�\[>p���;F����,�4A�*�Ղe�
��IF��a6��K��B���V[�?�>� ��n��6;T��USb�NL��*UY[��`��m�l�{^ES��D�ڛ�wiw�"rr6��#n�@_�e�	U����_Y<�[e�ő���i��HZ,�X#nR�>xr�Yz��!'3��D��1�n��	@ho���g���ª��L��M���p���P�P�u��#ߢ��q���0<�P��0�B�{��D:�˺ɉt�&9�X��# �͹���4H��B:�-`*�>�XD\P�����!�qC�Ǐ��.�N�-2<c�s��!_n.���T��OA9l����jO:W�l[�V%�Մ?�tk��b]��-՟�bʆ^dF�7���p�}�.
��7�%b��UP�YDa>3������:�)���΅�6xPiћ���E+���e����2.�q�3���D�|A����ډ��kJy�f~�~Qpݗ�7�W[�ƨ
��3�}Y����w���/��H�Y�n84�L}�i��U�_x�f`�f�޴���SM�Q��I�`�*^Y��z;�ۆG}��ڈ��UA˶t�ds�Fۜ��u��'���A�<�n���/.������nf�Z��g[tCM1eo��x3��^�����������R�V��n�x���m/S�&~/'/ʔ_�s�jKɪ �p��<��i8� *�4�q��6���Z��j���7`�YJ�Uu�E}g��w+����s
�W��Wz;Z�\�V�m���S�#[��_�s����7�[�rz��)�KbAi�� rno]�0�K�NJ�a�Z0�!3�:f�-�ң]���֠��£͘���UŬ�>B�AaG�{���K�	`n?�����;�lu�څ;3H�n_��ߕc�I%t�������D�T\[��wM�����֯�?TBKe���,���G��R��T̅Wk�w��������p���ێ�$�	\g�6;���?w��[�z/>�ui-�>��7�^��1;z�<���&x�[lr=ċ*cN�8���+�Y[���[��������Ce:3�I>]�yd�a�q�ᬞ�I�58Ԉ�|�{�(�ci�����b�>Pu��Ew�S��v��{>d���E�����rRX�65s�t??L�CB��Q02��÷�hG����AE�l��訒䔘d����Qx�Z��:gm�T�+�R�,�$R���3	�� ��i�*�β���ܰ���X�o+KL��,�0qƟ%��6ʣK����;�"��� ��,���I�4:��
��j�1g����*��c�l�o�L��6������8�N�נ��V�����g/	%0��s�����k���pU "*Q�{����`ޑb��
����߯�o�E��A��Q���PR��ޏ<LU���&w���Q�U��>�FO�Ғ�h��W��p��ǖ�n>Hz�S�e"��3�6����Z����mk�����2f3�r��O"�o��4v�z:�	Ȍ�p�Կ^'�u5�>i���W��+�u3~�LKX~:,�{��^��_��N�����i�~" ���]0��l��Z�}گܤ~iW��������1)<R����eo�!����L���o��%���DM�]y%��X�o�������"[�|C���ܒ����!.��U�	s��5���ި��Z&�.T^Ye����l���KνBq�w�����K;�!����E��s0���M�q"˓uG���-��A#|)��б�YB�ے�x`|B�`�2/�����V��ʙl ���5X�ԙ��2�~{������H<�R_4\������������4˵:��t�]�G�e��q��-䳠4������M�ൗv��4��x��W�So9V�2`;BK/w;��s�_W��x���Q/Bs4�b'.*���v�Z�� �jd){��C�V\V(���]T�޾6�EÍ�,.U�=�w2]�!�$�`��r�o�{ǲz嶸����xR�$�LF�%�����x�ЙM�������¾�<�=g�i`/�(����"�����$ǭTl����mߥ���1l���/o$�� �)��`Q�-U)ܷ?���h��ʩ&�O+�?k�^��lo3�ǎ��F�a�+�UG��M�::Ɠ_��7��F��OK�Yp1�%9�4��O&�~h}���A�!#+9S��k�P�ں\��h%���׉�M��� B�Ӳ�ڦVꙹ����T���<K1%��#j���@W��<����B�v��\0<sb)@Ǜ��>�@��0}VkS�7�������|�����+7��1��.-���B���u���h
�DWkv�8]Z�?J�®�o{����z&�ʼaKjh���v艍z7b)#���iߋ����o0l���!�g1���~��I��R]�טy.�\^�X$���J�R.����nO��ROx>��>��1&X�d�g�,��+���2dU�AMrbq�B�^�D`�����h��`�[)e�Q�W���+@ot�G�*���m��0����v�Eh�c��؞����� L��}f��"䑐��I?Mn���Z���� ��_ɟ����o��A��V��k�"�P�4��o�K�ޅ}�
�u�۝4M�~����}-��Kf/�m����!����!����螽�X{4�p/Jv_����/y��E���X|����[ьwE�����!����#<Z��
��c>1UM}c���g������|�+#��\�̙�7����s
�Vb?��@��ER�T|'���ӗ��X�M�I��%rv�US��D��Itgj՗������[dJ�!~���M�"H:�*����zu��-������d��f>��?��A�n6�\�5Z��ka�"dEm�ޱ_F�0}g��8��52��x�6N*/�X�*vK�~��Lx��Q������Mx�-�]Xo�ѹ��r`En��~��|,��!�6V�glJ8̯�%�WG�qս��>Sp�J�U�݄Il%�rB�Q��
��弇j�ġ��Ԯ��zz�@�J� �j�^����9��Y:H�}Q�g%��`VB?�ӖPC�^>���[�+�J�kUV��=�9ym3K�=5Q1���l��_�V>08�<��8�˜ߴ4����W���~{K�`j&s.Ty���e��zs}{��!�}�F��Τ쉕�a,	��������k-�1!�y����(~K�wq�MUnR1��n��9/�!R;\:�5Qtw��-�A����<�Kr3|Ͱx�`UݕxV�hc^9s�<��-��v���ӌ�<�a�ӓ+�L�RT	��Bw���)Vھ�ٯ��2n�����g����+���| �)��f�O�-��]!���Ϲ���p؟a=P�9�ᄾ�RuS�Q >�����{ur��]b���� �p�ʊxi���P��bE1��+ŏ�a�K�T���r	��.Q��|:zHh��-������a8��a*Y.B}v=���)d��q��-�y����U����h��9��
\�D񡢔]�F����^lS2�<\�ڪ�\�w�g���CL?���cW볳�wx�x��"�����p�Uoj5V)�͙5DaP�D��EmC��	��1���-��-b���;9���M:Z5�0u�ѭgbrxr$�ڀ����ӻ4�f�����C"�5b�"3籶��URU��䄛JR��"�V��N�n߄��Gs?�tB�{��f��:� �/��K���.����
O�0�"E�u�K"o�DY<�G�\����tS02��KW ~�	�!V��F/����w_c�R2P�0���U�����9�`-v�&e��߃��l�����;:��P��̧�����G/��i���������<'�f���ₘ@�~����@.n ����"	��._dw΁$�!���[;��<԰���|r7;�'_�=:�T;퇓�O�ْ�qxwAFYj��HR^3pe~���Y�\Û��u�?�P�b ������B�7�,��IL^�N��<��)J�E}�:=�ФCإ�l�y*����%?g��H���$�A1�N�άo~��������EDU�����j������۶*A�*u+�Nl����@5I�b�gg��}"=z���=DQ����=l�R�`v)��o�y����2C�9MS�9�G�.�5�q��- (�ݔ>Oe'��$YM��=�����2 o��L�ϋ�/.P�r�����k�6�|�Y�]Vͻ@&qܗ�*,�8��h�&�,�@�Q�<�R����-y"��W��6G��'�ϔ�Y�TIU�V��<	��(��c�g^|��P�������
��jQ��$љ�M����S�A9r���e���uAv���u�,�(n����ꀦ����	?")  ���t7���0醉����Hwwc�JLB`t�������|�gn���=������^O�7�q��&e��<sj=1�7��M65y���_5��.��j[����=�,H�p����5��nw��E�<|��K�Mo�2y:��w;'�ϘtA��|h�y}��g��H��l��E���F�J)~.��?Ғ��������)J$|6�����:�%��6M�q@`�澜��])/;-�دd�O�P���'�K��3@�h� >\5��(Թ�_>2��׌U��v��}�V�	��!��I
�6�{�M!��L�� ��:��{�p��o^/����Q�	�?$��E�Z�lnw�#��(�.�ju��HX ���`	iPO>
?<>azKA�Dy;X�p(���LR6&�~�G@�cB���5�o�>�\�l���Gɉ=ݿg�#UН�2�*�n�!�>2p仰`9'y�&�i�Q�9��_�t��s�L�^t%�W���S�0%����w�ЗR����߻ֻ�w+ �9��� ��s�O��F㽢@|�%�IY���h~�q�u��h�4������G��<��@I�^�A��m>R� 2�Np|vC A{B�|���ב�Z�2۩�Įгge_�G4�����՟C�夆h�w�>�#�n�u�N��q�+��>B��pS9�al���*���L�<L�**��VGD�����>X���JM3����a�
& ��G�0?h�Җ�&��,��Y��ov���o��w��ikW���\3�Gy\���ߚ��L�E��%����G�Z�.#D� �H���^s��CG`�bDe��1g��/xD�\	>~'B������o�B�-�$V^�9dij��yJ�z��_[�Q��M&:�qC."oq|���&f+�rS6$s�	^֕� �G}�uL}���V�H㷊��I���%H�y���m�t$8�2�wTC2��M����U|x�-Z�T[�eD�E�]-�����(\ ����.'u�;��~t?P�9	��vvNv��`ZڳW�8��1?�r��Wn�F��6��7���?=�
��_K��D�͊)�|�R�}-�|��#�w�6��-Թ�����z:��l��=qn��8v-g���D�����w0+����.ɐ��5(�g� ��ZBAr�ﵻT��}Hؽ�X�;o�ж�P������-��"byY ��!��::�Vo��A�̃�vю�l B¨�ڐ�ߧɽ��q�KT�~4.21��4dq����d���zVxחk�ߍ(�o��K�;<n8��㞱C���7"���J�y��Z�ڴ��x���u1�W/!]�����?��� �`�bғ��F��Q��^��k��l��d���j�#,fG�M�=�0~�w90���+o{���������El�eUD;� ��8aA�
�I=�	t��2�8_�Ɵ���*8/B��S5�K���=�Ù��:+x{ 9���_7��dHa �	֐��:c�~�ixvBoV����U��0�# t���䙮���ëE����a��oSr>�<��{v�q�N5���m���xm��"U6n�����h���=�D�g��pW�>�݇�0���3�CD�Ej��
��t�3��TU��"�=�}F�7��E���a*P0�~��gM��8Y�呃J������?9����
����R�m�G�^T�4�-��ղS,�;u;"_l}��1ӫ�p"�O|�d��c�3���9��f����pj�*��z{&%�*�1�Ld!�WqL;,3���;��N��A���C��8���>�1|�jV�o<�!�8����,�����TKEy^���xڻ��y�ӽgH��}�b6k����I�h��o�W#�?6�s2��	�v��@s��vg�L��f�S�;���XA�ϡ�SLJ$��0m.���Ҝj���tn�Pb�m�V�N�F�L�}$̤����kޛU��{}�j�`��Ɍ�,�DL9h����.PMI����awf]���e�n\���F| ���� ����Ǩ(P�;�Y/ϝ�3��ꖩ�gPe���ƕ��b!"�ZԷ�z膺���2�<��_Z:�r�Ή��rC�@�	�cϖuM5l��?c� [�Ю!�@�:��?����]�g��=�
t�6�1���ͧ@��`�y(B�PEܼd�]D�� &�a��Eƴ����pe�\]&��]�!Ã��x)��PVX�r���^Ή�/��Fw��*�>�6�L�Ͷ�捷J��~e;b�&�b��g���}��FL�� Pj�������m�%��y�y?z������% ��x	��L�Lj�������T���W�S�/J�_�����#�Rֈ��2�����^t�J�!�Q=j��[0:�� V��fj�:Z���V�j���^���M4�tR����e���w�d}�5B��4��^��,z�C�1�}���y(8�Gf6WV�@�wf�KL��������}��]��ׂW�@�4x���'��8W�,��5�"�L�8&p3���h� ���	;w"ocȘ�M���ѿ��}Ҟ����f�����ܴ|�I�g��	0YK�(��J�U��,�} Z��FI�E���Q�1���9����Y�eڷ�-E߾u��R�|fX۽̗��kzT@�jj���Ȱ�\�y�K�HuS���{�.b�~��I�0�6y����}�����S����� κ�4}C��AWG��C������C��x�EU��X��C�����cO����	�z����hM�_��x��Bc�RF{��?.��]^G;r���xv��܇5P��-CɵЬ��U�Q�cR�'� EX|p~�7��/���۵D�o`�����]z�!k�RS��D-mӫ�ch��v���J����3�g2��t45�c��6#SUPK�%�~�s8��g�z2t�;�q(�Me�Lz~Ż�_�o��'}��{Ҫ��N˭/U���
���\�N}�n<�LX.Q�*6�^�l��:U�Ctq������;r���Ot��]�|��L�����.}��`Eٲ���̊��L�=��_#�5� &�y�]�`l�h�'�W�[�-۫��_���Ȼ��.8Zv��$�X6��>1���;4�v����_5�AQs�O��a3u闼��B����������@��6.0IL-a;XZvif��YB�D?υ�,.çX?˷� ��P�"Տo�3r�2�bٔ�>�i�g���N�%�<'n�\� ϧ�_]e���5����1Z-�%������>P}�}=�/ٻ��}@��U��j����[���|�;:��7�\���'�VqD�!�߲���ǎ�g}ªX���p��gA��ͻ�����\]��[�l�a[��U�c*�������y�.V�?�;"���]N���Ŗg_��Dn�1ɠU��g���mvR��_�P��ŏ�Y3'�;5�٭�#�֩��t�9&t4J�A�>�D���4�­H�2㽐������W�_⻚����?�T��u3����֚�=���&��/*��WGi\s�E�)k���3�����1U�[6���;=�R�i远c=Z��{�I�L������0I��� |�W�����*�|�c�mLF�5�U#FC�-n��.� ����[�zp�r�}�=��3�G�`�l��N؃���|��;3���\�=���?'c��&b�M�HN�|�/ǟ|1C���x7`h�vV�F(�z=���fr��>��s�}�Ɲ��/(�0;A�q��X��!�Vꑼ�$��]N�\X��+=�D�B�8>J����T3�]i�E��U����	ӘȾ�Vy���PT5����t���ms/ ���;zQ�δ���膲��836}6�J�J����jc�^_R����x�wf(]�fodq�)�;�/�Vz�^���!�J�|�`��+���k��;]�B8�6!\�`�R6��f$GZ\��	\"=���fu�}-��BXq�Ca7����0�/�_����wt�/��\�W���72|S����5��O�ٱ����z�����3�s�rHҫ���V�'�#�}��m������|�Y�;��4��,��F?��k>�'3J�]�a��,��善��\�jF3�3Kc��Po(z�}��3�e����B�紤�o��/��&��!ip�8C���-�6��Zk4�\B\4Q�9��j	�]ܱF"r������V�Ԃ�fs����dF��}3� ����r�i{0(�1�>�O1����M�fb�o��n�9��d�� ���?b~'���C�b�n��|ti����;�?�4-4r$1�N�;S\�5�P{kDS���*U����E�VV�!��:r���p��j�D��,נ��|����-��j�^�0�U3}��m�o>G������pcw��K��q��l>7y/��`W�\��Q=��s19Z��s���M����d��X��~��^5��;>7竬!ˁ�Ej)'<~M���;�"ǉ ���O����qb3�2�{o�5&����S(�-��Q�Qe��fcdãrg̙�#[�n��Y�L�?�]�!��^S�Sg+~˄���2���f�\e��Ը��M�υGm4�O���{���8����չKfa �^:�a��v�
�ӛ�X`]�r��Q%���,x�[|7x��W`�U�/��¬s��:b�ڜ����z�G̟��R� ��G��������[���[��YH�Hl�ξU�=����?#p~q��f��B�X��5�o��7��Uv���	�*'��Y�u�OFĿ[&�Z�"�WYX��7l9}hz��P����;�M�@���N7��r�9�B~X�C��m-&)u��E��k �ư<nENa3�٨}��FE��J�.w�ۊ�)6�B�Y�m�ˇҏ9? K�]�'Dc%0c:���j��6�&�J����Gmg2}7b7Z�"̇H���&l����
�=e�~km!�!Q�bD�mӏf�؍I��Y�U��g�'t��7�a�d7�����U�3�w0��G5��_��c���Ӹ�+|�_�9�𡾔S:5+��_�+s^�z9e>|��Ԑ/#M�	�{�ޠ��uh���OH?���Tt�N-Ox*��:>��MAz�Jצ..���좔c,�~YЁ�+=��k[;���	 ���]��z��M�z{�u�r�^r�D�#�Dl���E�$�0B|&�yŮ/\5�U�?FҬ���~��o��X��-�)m�FE}Y5�W��ˢ��ul+�c�9�R���1�����޳)���;EJ�b���Y�c&9]:*�`�#�:����5��b�H7H����JFJ�&)^
���\��׺�lk�CT
w->���"Uz�|D�3e`�g�rJC1�l�VT���t�S���PH{���e�����?٣�m�3K�56��"v�o�#� �yO<B�7{=⩕��D:�Ⅲ&)R�iH�gi����:�������H��2A71rcu�)�Q��P�b�e����^=��[�{�.���&���h�%�X����]�qk�ݱg���!jJ9Y#w-���},��n���g�yx��0�m��������%�&���U�����Ӷ�;T���`���=m�]�֝biYN İ�h�b�V�:�0/��Ꭽ�3��!�V�4�J�<���۞�T��4|��o�hd������7��CO;,����5ؖ%?by��>�����sNv�Jֱց�((\#�6�����x�X�e�Jf��x��
����N�I��$�Ժ[��~�����Ю;�(���~s��0Z��g�,�/x��_�;E
���(YDg�y#��5�B��S�!�܂��kqx�1��O%7*�-���eN��W�Y�I��X�IE66��q.n��`�9����fܐ�x�9��Z˺\��A����o+�� �D���{k���2�k�{賮�̫�� ��0�|��M ƘǼ�EwƷ���H0څ��0���B�݃�ꧧz���t�������vѶ��Pu�*6cS���FZ)�	$���7�U^� ��qH)��e�:��#��E`I*��V!�M fA�:�_����#*���e���
�����k��VU�)o�ņ����g��Yb|���Zы�Zjg��ǧ�w?\�o���=Z��9��|��4��'�#Dz�M�n�>��F�@!���_��w6�vpQq%f�\����ޢ���s��uՒ&.�x�jF�Eϊډ�����:8�u�*'|�.vS�����q��:��?FD����O��4Apy��#��8u	��X��]�ʀ��~Y^�/O�h������ǙG�c_�v�fi�g�9��6�я���<�6_Fǩ�?ә@Z��]����x�{���Ԃm�咩���(�y6�����k}������r����H
4+/�4�fN�c7h�W�]����Jf���z�W���M��S	ͱ��P���y����o��:�"�N3�� �s�f�E폛`�52�4�zy}7?�Key��vv75��m�e���]�eK����ϡy��h��m*g�N�ی`�@��0v3�*�!;h�`|8��I��,�f�	�����+5}� ��ʨ�E���d�U�}qp����
/��'�Q�xnF��=� ��L�|48U�����_~jo���]|$o���>L�ۄh��>������������n��C�8�!�+*�E+��+1?�j��l~�qǻ��g���hc�\�����t$�9[bڋ�׶׏�,�,�<�]�j΀��$*y�2�Ct�G�^NL�f3z��M ����*S2��m��;VՖ	.�`��ܨJik����a��$�p����K%�"��[�6?�3�^a�R6v��DW����z��fd���@fҥ���R9��l�$D���<,C���wU�p�����cI�H4�s������V�GG2����_��ӗϖI��4�t~*����i�� �J��9Eي)��k�4�F���-��f�?5q��͸PF�i�x/f��s>.ݲu�$���!�6
W����G�%�6����ƿ^QR����u8\�I_lۖs}SJ����V�ͥU�.��ȟ����CO�n픜�R2����v5��j5�P"H0�Q��G���)�����2X����.���sz����v��+�}�Ǹ�Y��{�!���S�Yf�5`��rwB�)z?+����֋���^�/��%*�U;�?r�-�a�>3b�MY##�:��}�k[��F>v�߽�}��Ϸi�Y���P���yu���1�<1��k
���F���:r"@�zf�g#r��m�TB5*�$^�f��!�9����#���{�2tt�k��-S9��h	�;�*�@޺i�m�*+T �cTm�}d	;��P,u����XN����Z���[�t�R��>�>�4�Ԓ^������0�L�&��U�
�e<P�������xy=���=��2�H���#R���*�����\�,|�_?mX��B���r�DS��y��@����� �m�@����&�����D�����W�ر�
�"PΥ�Y�������jD VYN�R4&f2�z�r�����V�K�s��Ԍ��07��r�����:���$����~س.Bx�����ޛk��§�a�Qy�u&�mRȺ�"�Ӵ2��?2&| "��йG]רf�%������ʅ�+k4}���� -�����<��HUJP3���x���牦�
e���L}������Z�޹�G����(�����v�;b\x�S�>����[��Tr�[���,o�zDJz�`���N>�;���\�ӽ���h�wV����')u������@��"꯮߳.S�4u�e��D������.���\O�������,�t�r9��=�
�u^V{������F�CF��ޕ����}Lg���%	�a,e�ۭy�_���Z���?�#�����OE�"��l���c�x�A�J��[�2�(G�F��4S�ΖS�
X@Ĳ����^<��h�LIO�A�0 �Q�����S�3�cI&  *�
v,r�3ߥЇ����:p����׽�*OO�{�@�V�x�scZ'i9@y[����*#hG5~W����Z�9�2;���Gq�|��<76�~Zw鋐�О���2Z�޺�)q?���=J^'ڒ7���$F��w�������.r�|R�R�����Q���욬��::hO3E��O��������Cm��I0f�5�O��{U�r����d����9�������RU4�������Y}��|����J��yr�D�E5��\��\h��z]�T�7�(�q�k�y@k_���4Bp��K�O��!���1B/���$9a�qo��k�"������P�K_��e�b|�}R��X �$Ե�I��o�N�?�h��y���t���0�dN��l$���k?M�I��3?���u�i˓Ⅸ���cNEJ�]����'#�sL���b��΁_�j������=��KX[ݸ)��G���២�5?�B "d�0���&)�f؄Of;R���ԅ�*b҆��\�������M��5�7]�;���0�"C���^y�ہY��7�(���N�ѷ��Y@�����B41��l�숾�3����!��g90Q��w�]�v8�Ɲ'��]j�h�w2���N&�i��wX��!kp�/�Cz�&��In��r����n͒=�Y�h����"�n"0�����ʯ����ƫL��Ʉ��,�����H�p3���aD )���:d7_$��h����*����4�G<�t���f�W���٨ ��`�'�E2w����
/h)8{*�:�b(|0e<@�̪���*Gq59��� �\9ۏ���#�NQ�[=� 1��kVI]T����[�靧�Ѵ�DK�h#]���O+Ir�jK3;l��P��x�|h �=�d�����E����*�:��C��t�(��%D����?�_F��TVF{�{�ZF���7�i�$�Z	z�X���j�d�\j	�C�V�A�N�G�����V�|�?�++�̧��pF�`��� gq��#���4:�+I�Ұܞ�Nz��~)DG/n���:]�S�<��r�f��-$7~��jR�#��~3a��L����Z,}�0s"O[�����!Zq��A�H�ZZ����@v?}07G�g�3)��(5�g�����phE��gm
�#��p��A��uF7o�v�D�ư�P������65UUf��RpNr)�T'������PX�S����N��hj��˶�t��<�Aa���7~x	�7�K*%��-j�!�ſ�[�R�G� hUۉ��X�t�V�"͋Ӗ��"L����C.'�A[��~H��<Iu(	�JMM��.([
T�Ƒ�[{� Mq��g�-�ᡎlM��$f�O��`|.iҶ�1�F��Ierv��$y���Q���m9f5�#X�1��Q�T1�'� �'^ �7�!U���i±s#Cf�u��M.:QϬ���d@��7R���e�q�a�	b�J�����ŏ��]'T�D�l�V ]6�O��i>��Vo}u�^=�^)�T�&�� Y"��X����f��6=~p�%;�o\J�/�(c;H�������8-�Y�j�	��x��.���6�6S-�[c��.�×B/Q��`�\�w	��W�����{��u�{})�}9�g�;�k�ݎ�10�:����ȉ��3�e|#��,�$��G;�!�'��Q��[9�����<�a4$���~��t�eك� �2~�������h�N�	:� ��&�м����l��.(^�ш�6�r��Is��e(C�7�y�`v�a���{��^�19=�mZ�6W ����A�UH,^Dld��\�+����6�Q0�m���_>���UU2yW��D`Â�h6������6 �;^��T�/ݣ���(��8�&��-5iK].���@��3㦏Ao�8��i����/�oDfߖ�-��u�k1]�M|Z���(-��	Y��|�TyiN�7����KRo]���r��4u�D���1��B��2��ȝ����r��)��՛��ac���,��%�l�7!�
���YO{&~*"�����5O�5bKD���]���`���+"@�wxE�k�`��ܠ���.H��VI���ҝeG1��O��s���-	��4�Ѱ���O�����]9.��iei���d[������h'�d���G��_�m�R�ZN����ߥ������~F��߈T�W���ߟ-4�6�@
X�������_oa�0��T���� ��$U�R��0������J�M��d@�;Z��C2�K#1�=Y�r�&T��T���;�V/���ɡ10�ĄL�o��\�d�v��D�P1
?� �?_F�P�[L�G���?FmGg�������n�ݳ6���g�o>�R���w��A�U�:�^�2#������P��]���ڀ���_��ꚏ�2d|G�$�O�|�vw+t��(��rE���N���2���O���y�e������<C�o��"4��p|J�a���ϭ�Xg�D�Sd���!�i~����ID�g�J[�c�e�6�ip(~$��G��ƆL'������g�k��͈7�_���T��� ifO�~��_�-�C�~/p������M=�,O�ث�!`�-Qk>��jp�����P�1�s�"���7��A(�V�nI�t��@��h܉�5(�V8AD�3E+���y&���?�����`+4]8���*{]��8����"�D�g����,T��M����$bUU�S$5�1�(�,�T"p��ok�+�zˆ�䢿��C�{��|'ɳ(r<��v��R�PF�g��ʒso�B�&���me��
v@��툹r�7/L�E���1vV�Јy����9ɂ����v�� �y��MA~�i24glLf7\83#����^M_��i�Y�`1(O~})/^q��uHhH@��jNs�C�R�f l[zsqk�HOf��u>�O[}��y���*�H_�
t�|ux���q�g�\��Sc�%�T��>��Ƨug_�w(�U����cQ��.�Io��"�ۍ��@� �.��2H3�ƞ�)�G���*���Fᅉ��_���9��VNv�A�M$\�Έ����˛9���M{��/)(�S�pY��7�?��X��K�6&cczO���S�Q��B�=`���j/Z��W����Гs���q�kBM}�.n���k"�=Xn�R��4등�4��i�x@F7K9�/�d^�{�*���5(�b���}>rd'��ˡȜ5�Ň��:u[ʝ:��)�������Na��U�C@��:<�C�I��_���ŕ�Z-Y���?O!0>5�TX�J�y���0Ϫ:-�y�9L�#~C�k+��C6�/���Y�c��G9/��<1�m��``PN����n�Ƴ*?#�S��J^��P�y+��%��c�6FS�I��Y[I&W���A�n��rb��c�Rm2tO�ZK���@iO�0�A,�w&m�-�h8U,半N#<���Q�{4������iF�'�bpۓ%�<4��Z��u������C�ڟ�N�E���k �������L=]F)����!n]�c���e��AOK{���Nq4Ɔ�N��dF\w��1I��p$�=D�u��G4K˦����`�q�;�G>b���:ˊ�Y���V����n�0���@n �r��\������1B� �ؽ �A�ِ�a\cQ�IqE�pNt��.�@��3�"�1�Mz�8�ުSW�յ��/�bet�}�~��\�p�/&��[0�����-ݽ�&���W�S[S�L�����U�N�!ߋ?�B�ubJCH�b�Ҁ�-�F��h�qi�w����Z�(N����ӡ��K�=qU��g�����u�]���J��o���OɡSe�F���r&`O��zXo������5��q���:�?�9��SJA
�W�6�v��\�ށ��VNw���d�:�!=�x�n�U4u�O(�	'�b��a�3پpz�v�ɛ�&<޶�@�����(	~�Y'��%�M�4�����vϥ�!�5)�.�h�����FA�G��Ɯ�����:�+;l:5����ڵh�1��jh�}e�;� �)S.WU��o,����w��Bc��n*����I%���0M���ڽ���K�)LZ��M��0��VV���L���[�$�8�YĕS4��8@d���Ƙs@%��R�
�^�p��)э�=�Y���@�*D�{O&䗌��ي���T{�4�q�n���K����]�MV���9�-�@�>�}��#Z���X�Ax�Bw^����n��n�R:8��F��@0��Y��_3��׍���<�ӻ��ވ�~ٟ��x���P�;�G�9rʕʷ�������j��<ʹ��7�㎊�?��窚��g�āV>�u�$)�#	h�ns��=� �W�s��N	U�WO�x��{;���6&=3ѕ��>#K���XZp�Ҹ���[��+|�������i������#'�e��ODqEm%���X,���9�2��)���<��M�*������m�;U3��f��y��^$��n&q�d�u��"�t��s����c�;4�����kw�mka��G�� ,��=�z��љ��[+��Iص�ga�-E�Ԝ�ȜrT7�p���t���P��0�^f6�U�������l���/_�DA.&*��B\V���{=��������܍�^o��}�s��xNDD���%����	 �}&��T�\�]��x�K��N�����∧���7�JEk�;IU��a[��vP��%�O�J�]��+k*�ג�}\��bk����eŪrm�����%�j������;�=���x��ڪ�$��FU�J@���0�wQ���Mt��F�|�������.z��v���(Y��z��U`�fE߳l�sK٠����Rd�	�|�:K�1�X�Pmޱ��Ф�d7Q�M�E����R��&���J�+�rw�0�o1���Sʠ��EK>)�6�s<��X͒���pڍ�|��BoTMބ��(P�i �b�
h�%���ؠQ��,�,
K¯�μ���~'#���>�8���-ޅ|$���G����Ԫ�Icy�O�$�
��,�/�w�˒�����l�ȣʵ�u�6f��|�:��4�O�ʿv6��U���\�۰��KW�p��>���n�2I�u��n4z��.�SA��)�KO/�O9I-/$�ݿc�}�J��e��?�,㘨��&�r�;`0a��E�����y��c�J]���T�@Z���ɖ�Q��.H���E����&�S�VԴ�9%��8*��a�SN6F�u�ꒁ�݉
��Q���"ջ#�x�tϟ���W/����{��<R�R�Q~a�M�k�� -���᪙����,	���)���N�1��(^3HJ�'�l�jl2A'��?��[mhSw�?n�;S.� '퓛�4�z閉�JI9�`��&��Қ}`NAU�u����Rf��2��U�.u�&��k��4�ZM�ZQX-\�Gat����H��Q��Ξ8R+l�n���-��~���ʣ�jox�֎>�Ss�Ï��C��@�h�P"�9��ɯZg'�������[q�U�jT���N������K0�)=u�>��O!j��K�V�Xr�u'}a��},���4�����s�p��O�.oM/���EyK��,(MCV�������{]s~�k\� ?f�B�+�M�Ɠ��+�]J�3@A��w��e�0�;���ɥs��#�8Z8�^YA�~�]ˠ�PK   ���X8Ȋܸ� �� /   images/88c2329a-9b4b-47e1-bc90-005d0a7e43bc.png��S]M�6���-x��qظ�������;�`�݂�ƃ��y�伟�U}]�jUMͬ��>���U3�
r(��(R��J����a�7b�gD������3����S*=*!�Ǉ����GΟ�3MU����ݷ�ao	q�D,�$HH)�R���5���:եS��e��󪪃��RSz��:U����QQX�)c9B��� �$gqQ���/�K���Liߣ��������#�K��\E��dH@�R�?y�L��o���(&����R
�7���?��g'��,���p,u8��g�'.'�Uj�Γhx��������d�-�g������cn���T0����M����dءho	���� U>�2����6��邿�c�}O>�_�=���J�7���zG��}\_ /,� �ǡz�/���@1����_� ���Y�{���;Y���;�������0ɠ�}��-y�_�yV���Iڜ�Jj���!�J���z�8V8w�[�m�����o7�|�����?ud	�/#�3�O���ց�5���]ni���"Y&+>a1�&V�����X�z[l*hS��0���no<���	��h�<��a������,��!*���&�Z>w���D��vȔI�'���
�E|	�7ĸ�D��bH*i-���W�_Lqb�7_���_J��_7﨣"�'���������q����4.M�+��(�:MI#���q�S��{R����ʥ�5�S-^����°T񡌟��\�}\�)������y���Z~����ϸE�`���>�k�������h�y�A�LH�-5nBS���00�#�R����JqɗZ�Yz>��?݃ZJv����M��������Z O끣Y/�����Q��e"N�/_zmn�͗�R�]��*h�zrB�bfI�j�d)��ڇ�j�9��S�GU9J��<��0˄^��*����W8�[Oa�����Q�~-������{�oC����D�'��� '	�:Ɗ���IE%UL|X��C��L��*��45�j��ܴ�ʫ��K�,Zh[#�Բ�H�*���G� ��m�8,���)����?���������b�#�t�G(|91�$������Ӳ�Odva�
C��"l##���#�f2�`���P�'�N2��W�,r�ڙ올s�������IN9���������������"��?T@�����޺����p���y�!%�"��X� v��m����|
5�M�E��E�	�5(�g���BR���ny��
���N0T���9x[,]�|�\���Iv&��\���@�������"�=�WS��][Fyx��k�M��"��� p����o��Sv�]c�Y�ʫ���������C/�	��7��@}����3~�����<�m��/�G�?���R�����T��R6"֣�-Ӿ�_-X��h�ީE�`�|IFQG�*aF_�tj�],�è��w����j�򁕂[ܞ;�����������S�g~�w���´�x�0���r�.��""e���Ȋzs:j���8n� �n�<��%�����&���c8٤U�J`|\�O��!��BJ��&��F\�[�ے�t�����6��������b����ʶnڏ�t	uͿL.��آ��K��Qc§G*���I*7�U
AP��������Z�����ױ'>d�U��N�)j��.�[G��od4P�'��pf�;*���CNS�%��2g�T�k���X�o�m����|/��_�vezo���.�$��n��e�O���M擕���11���6^��Cg�!v�9qW���NC9c�����ސH8΋�
:�8��E��vB���%�����E2�>��<LGdݾ��J]�l��ݤ��w��� Z/���L�k����_�\�a��j>�
~����
x  _r���D��4�vf7%mm|`A�k�`4�?!���bW�%2��F���$(�*���A=[a��5�Ӌy(��ą"�j/wA�<2��~�BJPE6m���������a�=�]e���~�W�v���:�qQ��`�?GA����y�/��� M��⡢����`JW�s;��kX�����n��'��j�\wWuRIO��h��"���Q����3,�͇�ԏ��j/!dC���Y<yY�c���nԿg����e��^������|�q��f�}����`����B�S@�:Ψ�X:��Y��b:�?�P�D����`�xH�yU��d݂b:�d�
�h,粛�q�l��Z^�F7q����\Oq�����d��H��>Z�&Te��sø6�����VhR�?_���>(�N��ʇ��s�ƤX��=�,$����V:���ؾ<3�Q�^.������y�������"&�FM�������"W������Dn���XG�mT�?8�������?����}��%���%DD0C�l������q~������N.���
�������#��'-)�L�=����� N�Ŵ����D.�b�f�4/���֦T��E��fz<0��JU�]\ו�ݘ����Y�ʃ�����߆NV����^2��$��㴊��Q���9*�����K�{ƀ��*��D.պ
�m�X�dD�m��>�j�� x�Bva�3$mI"�9*�S4�D��I1�E�h��'hxgE3Ϛ2�c\%���}�iCD����~4���S�A6v�k��"�pTN��K�i��H��X�/Q��d���15��/���Ki�C��}���CD�Y?-����;�V��a�p0��X�n� �_x\f��BJ訛�,�=H�	�V騷Ru$�6���|h���s�)Bƺ�\�j�h/�,����::��0�[4
�0��ۏ��h�]��TWM^�N��}Ύ��]��>��	~�9� )�����)��W��Ft@���a�!�W�� }s����4��B�8H�i�l5:��B�`��"�Oh�zH{���J;��о�% �4��E\:R��DM9"���DX��]*���; �,Teu���B��M<xյ���TZA0�>񑆋c{=��S�9T�k���8u��}o�a~�C��J��1�՞7[m�%���]��FC�%��EM�#!-ܲϴytj@�P�.�Y-?&VKz���_�2��A�3A�mT�C6�=]�V
�rj��(��DE���B��"���'Q��Ɓ$�v�G�U�œ �k^����_̉����/7^;H^�����u����7���6�_�}e����|+�~F���ˍ����-]����4/n�INd9���a��N��g-*3h�����`U�f��]�U���Ru|XwW(y'�[�,�ӏ�0���ƣ��`�B�=<���L�R^CN�G�(���)ih5�	0"�ן����^���J=w��_ڶ_V�<��J�u�Þ��Y��9��6CC������z�w�kC-��.i!�JSX�����v�r�Ӏ�ہ�[v��׈��;��4ûiI�.=+����¬�"B:����H�6���-pR��E��Y�A?��}��tJ�M�`�FB�L��R���U}'y'�|�{^���H.xE��_9���<������C�}��B��bϛ��k����a��ԓ	g�L��t�ۀI�OIQ@Y&�OQKM�G"\G���WF���,�i�=�r�a����<�a49��·q�`X�ǣ"BW˄�}�GGX�X�O��s�8u��u��3�)�VGUo��s����srv���̥$sס�k%M��I�>��0<�G���n�o�8�:�߈$Ux����O��0�٥���Y��}��\cg� ����*�{���+�����Q׉+��Qu�jL̴ �)b<��hod�d�왪�ݭ���<�4_��~�4��Ru�2*dGX4��Z�I{�:0~)��cN�K��Bl,0���nb���j}�-p���"���"#蒮�}5rPY��w>\���;��g|r�������-�UK6�����,9��?3a�E1����Aw�&��1��\�CDm�;�v�<i�ER�PX�5�B�d����W!D5T^t��Ej�����y���r*)b���kdbsZ�*�Z�5�WfE�߂T %�o؀�O^e�l�BMw�ݶ���������l<j=����	gw=xO�o�w+�����x��d+m��Z���NMI�m+7�����u��Ie��r�hj궴�d�,����x�M�MR-�t	9t��r��j?Y�V+�Z�ذ	�m7
�V�X��֫q������6�2�ߺl<VQi�a:rp�n��3J$	{3�6*����;�s/��ٶu�n�����@�����gu�7��_�n��_�-f���ñ���Ρ)ş`dg��<�d$#
2�d �*���I>$�&��~F�Q�p��22T.�˺�h��x������YΫϘ�ƈ^�Q�	�xH>�Vc90��SUT� �]�p�:�z>�_r4��ٝXѤ�*/�6�t�mҠ��E^��4X��^ B(���,��r�u6�U�兔��/��[�>���O���O���j���`���I���_�|��H.�o�VG[Z�z(L{��}�-'�,5K�k�B/��y����c^��ԩ�t�FVԵ)��pϵ�'2l�(���ӫU��2��%�A���ް�k L���w)�s��I�L��z��Q�ލPVYǋ���t'j���W���ax:{�䡋�hM' �
���$QX��KK:Y�	N޷�~=M~���i�[r]�OG{%!?бwU�z_��j�����ߟ*
��>�E/8��Ѭng��O��ĀVb�>�1�.���.���k�0M]X��O�=�: �P:��K����3��z��VWM�F��"uǴ�y`���L~SU������-��Ȼv�ef��x|N3E��ι���Q�?�A���!�,�k�<��g�,��8��9U`��pNj�ݪ�@�6a���|�|2�t8�]���Y��y�وy�b4�í��$�w�I�?صL;��w;����1��	0d�7U���=�g��f�W�HvzJ�����f
@��3�'�9��G����k�������/�z-f��Zq�e��WE������������0N���q�*�+;yd[�!�I��?�v!5�2=첔��zYD���O�WAU���I(K�*�9�i�����ޭ���g�a�Rՙ
KΥ�b�~~����T�L;�����>�.s���1U=h���3-A������]����T�J4MW~����v�Ě�|7z�I��w:�q�M�:+�ݒS�%w�0q\%��P��l_��?4�)b���D������]9���<iB0��|���!&QJ����EY�����B$��*���{��Ϳ�&A�K6�{����@m�V�5�~ l�AuoR�a�ɣ�T�D��^:۴��h�4z^��o��N�{/��ʷ)�����x~�����M�m�����gՍ��m�QTX�=9�R��_⮖8~�QJ���Z-�_��Լa�]��V�X{��N@�'PO��X�i���[�p5�M��)���GL�y�Q(��+pgIjU}�X�Q��@f�U%@�e,��J^�#��77�h���y�������5o7
�<tN&U�d���
i��}x��n �����	T�d�V�Pvp5��=��*A��_ar��Ԉ��O�#y_�Ĵ�J�V�M�Jj��$F2cm ~�mN��L˯A˯!��kaǟ���l�����Ⱥ&���F��[`��:�]j�WgϞb"_mlt���R��9P��%&�̣�AKE��+k��H��$^-��X�F�*�g�
�yT�b��㖪���f'�$	�T�`�{G�77u��=��`��҆/=͋���:�Tǟ?�z�4ww3��x��r����6�3kά�o�4.�^*<q��aݿ/�z��c9t.�K�|z��F��=�5�6��˄�GX1N�^Wr��0�t}����e��������^�V�C���;�w����=�P4��������x߻��RvH�����_��.
�ݳR�7GPp���~��T��"�&l���{�m��15��8�w��:��	_��[s�:/�����ɱ C$5r!���H��]I�Q4��/�p��C��6��+NΛ��=\�$��Xj�*ʹ�P4���a��`�X�i�9:�ߒ�1�Y0�%�`�I��'�D��+�mZ�t��'!7}YV�>	�t�S]�ԔU�?����E����a�qTY$n�a�����䆡a>eh@��<̘�� p����T�+�jԃ��մ��ORN�~K	f����pb?��7�_0�:�7�>%��K�ٹ�K-�2��lr��3����"'��ղR�����FP(�(�݉]�&�o��&��Ż�Zo&)��j�!@�Z&�K"��g���_b�ڬz2]��`og��rtl�� ���Ӷg�3�l2yB|F�E�@���Q�!;yA���������a���=��
A��!5�
y��Ux K(��e|�>j�[��3 �~�H`��?����Q"�{��9�zB�r|�񹸩�`�h�l��=�-��T���g�����$�7R2��� ����O��kn�s��kTbȐ�\��Gik���"u2��t~z\=��`&��;=M��wn_�,�x�3��c�ێ����o�vY�a���^�����R�`�R� B�}>�{u�3�3�����t��wFFF���\tLTk���7�+�4�$�q%s�K'-n)Tf�z�b\2�!HoSS@���P� ��[��d��N 7��e��K��h���\Fǎ�|*�<�~R��KI笩�'���
��~��nJ1^�[�u�CtI����&g'���ù���&��y� .oo�2����!�R����|2��.iŃs+"ի7	��1��7�ݸ�]J�qR�
�G�-c)w+����i�@G)���-�u���K��,쇮��gƬ���������fCHucz3e-3H�3��>���m��ٜ�q�2a�H8kj1F�:��r�ڤH���`o���@��^�4<���ƭ�Z�G�?-����Kg(6��/�.��;�r�7>�(�b�/�p�*�hL��!��Lg�����5�g��St��c��@O��܆{����R
{�����_����e�����@j��'�I�P��|����	g��W\��4�V��T��3�
��[���9�۾z�q�o��Vt���c�y�q3 ah�!N���v����������x�c�������	�)Wt��f�߬��X�Q	ڇˀ�oK�����nǋ������N+c2%�?�r�=��6=�E�$�6�0��M��J�i�(`�]��;�r4��������HJ(�4���q*��/�~��88��~���e�\����+�T#:q��d�a���G������`":nIU)�.�1OJ��<<�T�j��w�M����F���'�dG�<a�l�j��:i��Y>})]��LͽL�0�-G��a��0R�B��@<����4A2�vNJc�3�X=7�qv �t;Ű���6J�>x�	8�Sƴ�T��Z��Y����v�%'}G�ޗ��q�b{C��p��R��EE��&�$����b�	^�np�����ݠ_��I龈�6��j�fog2��PW�?���y@�0�P�A` ���[�� �Rvye�3s`�1����������k�T�)�z�Y!�1�kh&��6�"����y*y�@�Y��#Sk����H8�v_u'-��SG��f���l�_�)~~2��Ym�9�'GX���ƞ�7�3�첾11B6���G��>��R�s��ҥh�������6�B��y�P~nR斧g�/��6?>����:�D˱�Mx1��z�d]S�'$�+�&����r�E���'�h�j1q#P�/�"+*��ަ�I�_'6���Y ͯޅPe&?D#7&{�i��JB/`_f��=`c���a�w� �خ�\�OW��`��3�_+>gi�͘��Í$���(9k{�XE��6\���N䍴��v����L�5��	�Sw@�Q� ��̕��ũ��x����^�(9����N/�Z=t�Ҵd9�$p�(x�Y�r�(;�W1��l]Z�V�=LY��F�{ox� ����lB[�b������Yh����m	���R_��2�6͛��8�b�ޙ��m^�%������g��iQ!�<����Pk�w�'����wζЈ�P�Gn�Z�ݭ�����Ө��hz?�Nr>k�o:z���jt-�0�p	�p�۸��v3Wl�}̰��Dv�^�CߐC��Ո�?�g!\��XO�<y\g�$�<����z�	�@�+���G<M�y(��m�h9�=���]9b6O�7kё����N�곹c'jZb� %��قHII]:gje1i*��F�@g���D���g��%���Yt w봽g���"0�����n@XF�t���ˢ
��%���.�M^��J�u��Q鍙��^�$QX>h�p�ܩŴ|�F��@��o�'�ݽ�I|���@a�8�)ᖆ�c���"#�Ɇ�ꙋ���B�]�$�n��>QWX��tp�)�	M����5���F(���7�;}#��=q�3�\�
;���ʐ���8a���I:}���[�N/����ي��-�-7ȁ�KNR����Q�*��*�=4��,�TB���[c���Hz�	��0&2�g��o��"WK]v�)����nQ���q`O��|4���jfQ��X��*�v��p0������^�iBm�]3�	>�u���a��[e��ǧ`��S^Mo~̅�����p�n��D3HTФ�v�˨�GD\��̀�Q[�%5�KR&ɤ�AS[Q����(C�'���H��,��3��G޾?g!�����֦��=�R�O	H�i�#ڢ	��>��G��J���G'k����5
ȑv����P�Ye�mK���+2E���'�m��!]k�a����!1co�#R��X������@2�d5$�=�"75���<�ߒ���ao�V��V�m������������ڃ�<�ۺ ���xr7h��#�|"̎�=�ύ�s�b��htE�md��v��Ki�@�O�ː�8x���(0)<V��C�1�7h�a���4��/����@�mu���v&�T)b�c@h�0\�ФE=�,�~��_Y�	tdE�$��=p�����LT�rB����0�K�O{i�Khm���a�'^@�坁�+�����dH2.4��Y�N,���$f42�o�e��8*MT�!��%܊]F�)��N�^6hu�nŏ�\�� ��8�B����ez���cۅh���Q��^��E�:�8n��uQ�Ĩ��!b�43������I{t��3}D���]�D~�*'���5h��`��k�`�7�t�s�-������9ݻ�
C����L�z��=�a�e�}C�������c���h0��*����/����g$.k��03��4B�:a3?~�l�OƇ�B#��&<�LL����\{5`��.�l�i	���;�M�j�?c���{�2z8%W�d�����Z�=��n�D"?�^ D+ї�X�­Na/�E[͢�F'':g#��'��;��G�J��8���,ꇒՇ�J��&���J%���Y�O��� �=�En���[zx#��
y׳x��epч���f���W��&aŅ(����j�B*_���~�R�W1.�f���h#�D���a
+�m��3�N1�h�h:����FF�.K��9Q�X����Wr����&��z �DQ�4�Ƣ-B�2�Rv�'Ē:mYy�#c	��#��Ur�!�ޜT3��u��@ێ�����4�$��؄6�6���ܡ{��_�~��=��fN�6�F����Z��>��Y%�M��pL�9Y*-�4%��P�(�t~�O���t�I������N�Y���ٻ5�(m	�U�3����o��<�}JH�������wv�6����9Xࡥ�QZ�x+�e����={�1~���jz���sp(�r���QuA����^�끎!�'��$)E(u|����	�	
:On�厓�(����
�<Fo���>f����5�U��.�d�s�U��^�_s=��{ٹ����5���rm;8G֍;s�qt�q�e��h̃<V#'*�obt�������WCn�ڌ���)qq�
��7%oմ[p���m	�	�^t�1gn7�'�[&�#�_��B���+A�*%Ž���4�EĪT�����%��@3�Zb8�7�H� ����o�F�@��G��1XG3t��KCZDO��A!2N����>zE��xUE����B��Yx��<.��W��X�y"�'xf���@�F+��,�{�躝��-�S�Jr�g\H@�7�@%�	�a����**1!*{Tx�7��g+�9b"gA���ZE�y�&-s��mg�� ���D@�|�G��A�+mˍ�6`� ��p���e����ά��c�Ё�&� �U&����&�-��_9O�)َ��=�М���7�`��3��LdXR-gC�����������#����5�%r!R�ZlG�	C2ɒw��\��z�ԹΌ���P9w����O^R
Z�"��h&hW�D%���2�w��s�9��:���E�E�IW�Y�:�e�kߥTt�r�l����$��iJr�=7��3]"V7&���By�� �����':�>0�-�ƒ��������̖_2��t{-�pk1�z-��N�1ڃ�^z�Bْ��x%��mx�3i��r�K�1��s�ݰR��N������)�e(�;�b�x~��aX�C`��z=Ѷ�8���i��U,��r�������I隟�=�(��Z�hSy�������^Ip���77�jQ)v�q�h���7l��V"&;�+��)�S��U:G@m ^�I�<��>m@4 ����r��J��9>ʱ�]�|���2yED������<�[�X'˃��M�b��%��7H�@N���e
'}v<�w6kL$��L^���s�ɏ�� ���#�i%_�{`�%ڝ�In�6�x�C�Jf�����Y˓I����1�7%ķ�c�>��'�>��S�|}�\��y�R	�g�W�
�.8$P��qC@��0 ,b�7VW�(3W��e�p=�67].(|�z�*�LP�B��#��m	��B\�q�58mz��E��3�4AA�0y�k:�ƜYk��6o�O8�H[?�lƪB.�5e��\/���!kM$v�I����� ����*�K��/Y�cn�F�*1[-c\d�3Z��,ڑ9L��b��[����7�vδ�[t��/�%D�K�:?��v��ՙ*�C�����/�YV1����&�~-���j�=[��g#˪=h麇?fz��;Hć�q��g����<��[��+K�6��P ������]����é�!V~�����%w6pU��=�wP��W�����4�GFr������`A��h�n�G��q�;kkws$�΅�s� ?'2\a�O>�/��B�o�����襘��G�����Z7qjb�� �掠�G'���ɼöybFB����E�Č5���6�%��,4	�/2l���ez����N~֙A�㸣2@f�zM�P�lyǃ	p���q��8���}��m�\E��7�*���gX�i4Ĉ�s��>�7"R{	v��$C����̮��@��<| ��զ�K�0A�"mgi� a�S���3�NT�����_�1����x�_�/��a�����< e�ɋѧddO9�"�!:9o*J�e�1ho�x�WO� Bn�^'v.�t`&�Ug��\K5dG��}��굌�fc�x��>G��`e O��Ѕ�Qo�wP?��`�+��_J�h��#�Y��ț*wp�] 1a��4�`G��r��'L�^T�(�/�E2���U��B(�\���sm"��0��T5��&���5�W:mBҲj���=�Ӕg�8& {�e�u_
����h̲]f��	g��=�>�h�j-~�,<���b�w�Oؠ�C���í��
��l9�W��ޱD��K�F!]ԣ���L�ˆ���s�[R)��]ϊ��J�ZHK���rI5���J(�͕nxB���_P� ��=�^6ʍ�T�����\�1�7�����g��$�c���Va��-�.�#9~us+)�U
_t*~������ܱ�Qh.w�������RC���æ4ʮZ�	�hQ��)$�i���G(}�c�e@�~�ǳ�VQRВ�󳋎p�z�5L/�s-^��n�� �'��M});5:n]�g{�P�M��l䕂��l��A�R�wޯl�P�����S�����RUb���OU�tŞM��R���y~<���LY��T��N�J65��h����'Ҥ�M�.�[��^�~����;_F�k��0����/���R�j;I47<N_6	nĵ}ҨӬ�2�o���L����i�'�+^r�er=�Z���f��4;�{�f�m�\ �bA�[�������S�dO��kУ�/Z�6�f�u�Հ�;?��9�%�s�]	���'�o�N8��y�ιw�, ʾ��T��%�M�������EsΓ�m_�ؙ���̭���M�S��A�<̷��_���Iμلg-n��*�HA�poa��gXbf���t�%ª{;��L�D Sޤ�xQ��'DD���L����K�#���T�#ƃ7_Iɶ�{�hM��\��8�b@e��͵mĮ�=8V�6����T���9x{ƣ�b��OH��⏲su�x�)u�b,� h<�׶�<��" ��㵺�د*��'Z��^WGwIXs��L�A�$?҉NaI����u��Q]��JHJ�~����!a���^�j��g��:��v�P��|Nux����8��H��Q���c��~�+=�̰x"@�|\�?��|H�H�Z�R�9����YS�*�w`�R�ߡ�t��2�ޠm���w'�?1�eD ��ˢ}ц�iAϖ򿊄jB&ݛİZ���ґ�ͳ�y�~M2������<Z��z����KT눟��"e7[@�^���2�i*����S�6c���q�е+i��&i��$n3%&�<���cn�4��;u�G��(��Cۣo���pv�^�.���Oz�A���ov�39v�J���Al	�+�R��!��=_�^)}���<�V?k�@��{��~�	՗��]�>��=S��7u�Ÿ��[��Bq������h�1��\G��f�uu�$��ش�00�o�a�Y�1N�b^��s3��0[��u�"$O���[w/��4˜T�@L͡`z�ca��r�
�"�4%�ak��#�ã1�q����7��V�'7�p9������t�I�S��4�|�R�E�����gf#�?HEzBj�	Z⩧zN!�nܤ��0��]%6���O	���aD�}���8n)-$�rNm�Ya}0B��b'i`Q�� �Rk�g �P�H�g�5Ps:�8�7�����V���z�E��VJF�u�����ۛ�<��_��)�ˏ�	Rћ
��@mc����/M����1
��]O���I����(�x�9�a��>�|����M�� ��W�r=��c����)ՔG܍]ɖ\�f��>�D��%B���� �������6Q�*���$�^)��*��c*�gC�T�����d`��-�c������'�%R���ٹ���E�>"� z�YYf�X2�S���UGR���6_�aT5�/3X��j$�\R�&V��'Y^�ŋ�I.�f��A��6��W��6e>��*�U��2S�R���Ù�C�_�EiNR]�R���l�����2�_4�%�k��.L��*�é.�Nת�I��:�G�BC�\g��=�(f��Hj�FO:Mq��4��u�W��Jgo
���(��]YsT����>�F9k�0k�Ӭ�?�o"d`!�G�A�RG�.+N5%�p��~G8i��*0�kKMS$��ۉKF�g �C'̢{e�v ��梸���>j��b���y�v���}
./m��ʫp��Sh/*��)Ӷ���@[���
����Z�Q��B8�AAI�� �nU�ch7tѱ6�ե��5��T�h6��k�(*W�OV|� �j��C`�ކn$Ó���P����� 3���b�=HM��=�Sx�-���qe����VAK�l����¸�|�˾�B�FR�:omq����{�Z�=\R��t^����\��x7������ΎR-��]���z\�٦���9��i�5�?[��ћڒC�It��*Y#�Z�I�݋t��3�A3b6���Z)�z4������]'<&J���xG�����mA�	�s����t]%�n�V!�D�`c߲��~6�\��Y��&=\�,����*#S���
�	�����Ƣ����Rԟ�N�{T{�@�+�{寮?�356\x��a|���u^��5Y�n3�(pw�����/W#�����h�T܅s��>��Qȕ���-�3y�ծp:��¬mt&�U�8��0E,���#R!7���J�lʖ�%���>��f|���1>v�q_a�t&m! �t^����#��&I���sWFt����;>&��z��^,Z�{�dx�7�!%�9^)���_�G�xKv�x�ѥ�4gIcp9��G3��_�B��;2�%�rA$}�c�{0n��3�#Hd�2�5"{�줭�Fї��pq !I�/���L$X��Ȋ�����N�t}+HM���s �XS��eBvv@�M���2'�����i�(0G�s2��m��R��64�*#7F�"i�C����|�A����g�'�������&��/PM�Ή.u��'ND���H�S�����ts�
z#�#���O��� ����ٜ�.�v�����~��T�mb`��U��Y�1<���'v��Ή�5G3�$礰$��7�6-�l�V���֢�V�Ūp�|�>��U��o9c�v��{���h����� �怪�J?FE��Q�������%���p�'EZa��,��G�d���A  �IԹ��Dt���H8��L�T�c����񵺮���?�Bg�(�%��8}>�)�AT�١�v���9�+��E���9����|��w* �Z�Z��)
�hP'���;�B���r�Py���m!<jA��]�]gI�����tDn#7��h<�R�b����Jj�� 4��5�q�TUrꘔ%���-(���)Ӡ�%5\X���+@���C����{�����?#Qfle[�\�M���F bUޭ~�4�$��4��@�P�&�I�ֳ�C֞8��E���Mk|������l5J�0�]Aq�0���
�x�XIOV���f&��?%��G�O�(ь�+���>%iz_�d~��1
�j=��a�]����g�v_,�6QZnZ�(�� ��f�/C����-�����Pb��h�#jy�
��8)*P�����2P�
>�Pv��0�܊�4��(�,��s�Ť�t"1):Vj
ŋO�DeKɔ�`�Qv�T1��x7�+�++�P���15�Z�*͑��,�%R��Q��a��� �HbG������ܡό��n�n)"��.��XM��=���J%�ؘNXV �S���&5��؈����y��E�B�I���z%a��'0�gy����~�e6/��SkRX���¸�q_UR��G��=�D&�T��&�$��}�p GX��<�ϒ���I&���w+��&l��wl�W�4Z�I�Z2��Ek���R��#if�M��ΐ��r�,h���ځ	��j�8b����&�`ԥN�u����DŅ�s�@��!)�e�QS-f��=� RD�O�R����?RBV[��`�y��[���I�+T�47�I�o���Wѧt��X�$ַ��
�@�#��a�%�iH�#hNl<�$��IޤѶ�\;�A4��$�c�jǱ��o����|��@���bqz�֋��4̋k�ÖOn�/�kƇ�ﴔ��f��׀<e�'9�?�c�S�r#�=�;�֐� ��Gj�K��2�n%�'�@$i\�L Z�

�UIg�b�c���ԉHI�}C��hfK����9�y�`ͨ�5�����k�,�*gF�7I�@EmT�`d�9+�b�+ ����+6���J�24$՜q���Q�f��ɈR���$�ɢ�`E�ݎ �\�N=�t�*K�ꞣ��S�&y�W�)�o!M́@��{�p��������1W~p����b�bK̈́(����O�ËRc+i41$���/�_��k¦!�4�*	��RB�uj���XE� �k�?���\b��`;���lt�ر�Jl�<D��"q߰D����MbaE'����,Xd�JS�l�)�l����X��h7~KF���qP�<�{&���c۶m[۶m�v�ض�db�6'v���w�?T�[�Oww������aU_3�԰�B���y�2�m·��DA�ʵ���v_U�3�%�KB�L��3j�"�����qܐ�LԂQU	܀q���ٙ#��+䉴�"�7�}��6=�i~f��AA�&�1�Y�
=���j�����6Iޠ����)ad��9�CΕ*G�.�
q%2�?���c!�5��uEx���r������x���ܨ��r��ˊN'��}r�������@�	<2�N�{�`W� #���*f�n�Zd�F�� �~.=��vQ9q���z�k�j���vW+�ʍ[-���I�Z���"�0h�T�vJ�����"�oK8T(Y�:�ʉ��6�}�t��.�h$oc�_K���>g'�֐�H͋��$��^�}pT�p�`S��b�������bd�d�Ls��P���84Tsk8�e㶜��]��k˨�[ܐu���X	C�*̬.�	&��n�"7�t�|�yR�uΗ꣥dp�Օ�F;jڇ~�(B������ �"P�Jjgvڲ&s% >� |f����ӗ�6V-b�Fؗ�����%�����8+{��E���M
�����1��B�&�B���|s]6i���*=;�N9M�٧��m�[�ݹ�Y7E��M���nkt�:�eQwml2W�aڋ<]Z1�)޻��`P5���s��  ���U���e�T�ra>ҟ���Ѹ�~�� ʅ���/R?�{a�v
�θS���V���A�f�d�v� ��md�]Qm�o����]����A,�"��3������x�r:r�3���z
s.˕aT���\��X�M�|�ơ���H�ߠ[�|� qR��uv��H�?O�Ӟo����l:��(���=�\��e�U:�,��)_2�r�e6]skǀ=����C�[�,�:Ƕ�Xe�]�}m����`~�����s���(-�r4����x�9�d�K�Of� |���ρ���KJ�BNɌ��s�P����qo�|]��&c��x�9�J;O��HN&�LŠu�[FF�6=R0����:���k\؍���%ބ��;�	���4D��0$�"����.�+:�y�y���e��W�p_dt�X��9�~�D,�z�1G���ٓq�]�n�[a�Z|����x�IM�ũC��0�)!qKO�E"J�9p�6it�:�=z�8R
�:M�S	G�p9:�O��C1���đ���L�w2��]m[�dvb��XQ<�0�����b���w��m���Gd|����*�6Eץv���7��qr�$Ԩ1ҒK��d��Y����#�2���q�c+�YK�?,��������0M`���fr�+%�-5��ޘ�u��� m�e�Zt:2j8��r�E���	q���P>�Bznu~k#��_����	����:VwFb��>t5;�k��W�g(b�i*���ږV�V��p�Zz�f��ʛ�;�
qm^���V�L�o?i�F����"��|�<'�r0�ׁ˩�ȓ�"2�#����g$��9?%DbD��
����>��V�oG+1J�F|��׽�~4}~߷H��q��[�$5�e�i���DlMW�?�q�����\�0��>���S��f} L�`q}wI�O�$0q]4��w#��в���8t����?�(4��0��aIjш<���K�����^��X�K��8����s�=����=�z�$�M�>��D������bO��X�h���>dȭ��Z
8���N��KYԐ_�B�~�����i�dX����B,9[�R�-ܚ��Ã@�TL��OÁ��f�V+�=��"}�̿�]y��n�Ȉ����tr��ο�V��s^3��<%�鋯�+q�˼���y�(-%�`&����W��{l�-�Wr0�ڼ�(�&4�7ߓg{�_���e7��ǋ ��й��<��{�,����z�W�fO�>I{bh�W$b�ׇz0�s������+I���?�)�۵鸷yQ0 �q"�uD�r�lT6��sa���l��Z���ue��Z����ۯ*t1⼍�PR�wP|V�dT.SfhNx�Wt=;8�+�K����0��ORs��C$o����NpQ^��%�6H&�m��Yv˓n�D�Α�y�ɓK��G�8�KB��rV{mH1�<D�5:��F6'�(\4�͞��5�I)]h`<3�Bn��UWW��7�(sN�3aRm_@c�0�X6̐B".���[��.N��?�ULZsw���J��[�"��"�g�A���`c��"qS�"����<�m�2yfߐn�$�H8./ ���Q����:�'�n[�y_:㠈أf=��_�v鐻��Ӄ�KWr��I��]��T����X.��/Zry5�w���r�V[ni�[�Fn�fdzmvq�`�!��#�(��N���	-ӎ��̍E���Ҩ3�شI��$G��O(>�<�X ��b	X=8Q�>-��:�_����"B="��C�v��޻�w9}Q�(�d�Q�]%����	I~sSms�w|��'d�-[����S���w��c:�Xt%��1�L@��SL&j�r?G�tF%�m6Z�R�W���`�,ߖ�ź������!=�=W��Jh�)I���D"��;8�X)'xGQH9�O��#l���[Ξ|�g+�:ZOs���?�!�}#O&�z�y����{O��%�5��K�89���]�.ۂ!$�9ɟ[%�x���h{�:�1���J��q���L�	�	Y������/�ҵ~�,�Ћ����̶Z�(kA�	ۄ>i���P��iP����D̐���U<S�>�x��V<D 24�㓈hj�A��Rd2�Y���y���uud�Eb��GE"1��%���t���-�욦 ��ׯ���`��}`���ʎ��m+m���l!�,H�R�D:f(�R�g����~��0�&^���@K{H=a��Z������U�Gy(0Ռ/#&�6xI��S��t}Ov�tp��L�{Y��wƢ�9>��1a��c.�2b#�6YB}��z�_��ɥ��2Y��H�j�\;��U}�hoN����,�obx{_�R=�3�o4|l�$�2k���(�Qk
�C��Z!�񬎎�uћZ�h�Zą��P4g6�7\juz��)ez)���A%��Q��}{�t��T]�N�n�^Ŋ����]��F(��
t�������)V�,n�<��-e )>D�%TI%���!
�����W���Z���
ee��+LdϮ>���n��<{�)ߝ�U�Z>����կ��n|��dB��,(�=��PJ>�]a��Pks)dQ��ɦ-BW�ȓ��s<�W�C����"aW.Zym|�Ax���W&�c "Π�P��}����TCtS���,G����e�͊�i�dR�ǔL���^��l�}�:=	���z�BQ��WHn;���T��J������{�f�e��LwQ:$,Ϧ�0 �6��&�H�:�m�'ʎ�x�\�H�J�s��t�D�Z,
}�$�E�W�?��U��(�;����@ϊ��ḑ	�#�j<%i�^�i�~��_���BEFov�kR��!z݂��w7��?H��H�D2�[�eϷy�$@�v'i�z�q��5��h6�w�S`�Y+$ki�Ґ�y���k��P�|��7�ePy-��[���s����*qn�神��Bw��@mTrȰ��A��]a~.��vo捰i���d��揳E�g�S(��VM��?��hh��s5D�ӴgY/9�"1F,�Ff�K���HCRPA/v��
�̈��(���Pa�6p�3�w)0�h�D|m�f|�S8��c��YI}������I+�o��/�s�n��Fn*4���^�Q��C����"\$��@\�D������	�_���W���eߘ��6i������L�ʃ$+�9K�md�C��D�@"r5 ��uv��`�ǫGIS����� ��P$�)��QM^���M�+�����ü	��V�&)��R6b�=��&�eEB�l�=�>�Һ
N���:�ѡ�4���]�#RMOko� �LZ�h��6����'���aa�_A���%X�?�W�ш$�jo��`�X8^w��͍�e����1� !����4a9�٦a%�ϋBg�I'��˪�>;�ھ�Ro�mn-���3��FC�qb���7�2e�e���%��NWFy��mT�������.�	[�G��m����C�B01"19*˩�'�~X�g��MQ��PH��y�C$��&��'�-j��,�\K.L�#@�d�V�X��=�e_Îu��6��°�6%w���p&Tcӊ�7;����dw͆u�r�r����
�A0W�5�u�qk�bu����4�|/���ڇ�9q�:��f���Gi�(�F�9b��]�B��G�2�� ���G!��z�ŒY#��N��|��5����&#�#2��)��X�|����p�Ct2�8X|���CT]���~U��x�\t�n��K��ǳ9��;NN2���t4c �HA5$˸����k�u���"��6�K�F�D��t`���DhA�S�ʜ�=���ml��g�d"�JIS��Z��RU2+��&GM���'�C_hd�fp���^{<ǀX���H��qO��]��]�l�ڥ��*MJxz�i)�w�ʭ�W6��`yyJb�Qxs�՜8TW�f^�TIZ��@m�H�)W8�q����%���/��/j_m�Ϡ��g�.�\�[��ws�o|��v�c�H�J�S��r���,�
'��Rr���Ą��s��U8|Vz[���L������>C1��d�Z���q�xC�q��]�m���E�֘�ZI����=X�;{^$�*~��zi�b�8��1}�>�2O��n�i��B������TՕ����7Ap7�)����2�$�,� �Q4��W��['U�mK�X6��4����4�Z8oQ>bH��4����W�>||>�ĭ,��O*��*����S@<Ć�SҞ����$�[!�X�x��6Ƌz�ݡ��XY]E��+�z�6C`��,�U5
Y�6��\b�����H(Zxȗ�]#��q��Gro�`�y�Qe ��S�=��ZZ��#KV��,G���`h-
S-�%'wROV長�^K�<�Z+=�;:<B�1i���;(6��m�	��pq;�<SWYUU<�✂n~�ߤ��<}X(��(i���LPk{]L��`lx41)�r��}���%�� �K�O<�\Y��6�.)�ˬ�)�G� �� 4,5[}��/NxI�W���+W��׍�eZM$Nt��lnƀ�wM���;9���7H���Ϻ��:C���ؽX�hA�F�g���eɫ�4�+9����ֿd��uOK�'�S�)WE,�P6|�J?�����Q��m_�Ivb�H�G�n6|�u �{٘�t��b61�$��k��j��������`��\��Q[����q�z�*y�'��T۰aWo�k��`u�Tc���;� ,��P���q�?���P,��7����
#�"�{��raʽ�$�$n�ğq3���.Q�lh8
+J�����l "��J���J��q8�����Y^�����k��ڞ�_Nq^�s�h�aU'j��"�	�u�IUYR�}VìT���Ps�)O[�0����i�@G��G"iN��r�ľ���D�L�d%Z���HU��(��
��"�z�r���K�-�G�7�y�@�����yۮp�ПZ�c1�����Ppq��E=���6�0 ��^�tsٖ��U)�>ң!Ӷ[S\���ǲ�Wjb���0���;�)CWb8;_�i��lndM�<1|� �p����T�S��q��n�Ą���ý������D`�y1�Ʃ����_2��;r����ʐ�2w@�h�K�赃�>��8��Y�y���8]���:fK����v�3q����ź�$�|cYRG�/�vT���>
��[����x\�-�J7
����D�L�Xo�����V�2���^�_
�>L٪�'�/f�*�[ tzd����IͩM��� �(�������˫3�Um �|�^K�uj�����Dj[���^ڔ�<JDXt��,�"q�iZ�̓�za�|9b/?cC� zq���\���_�fߘ�P� ���,��G�~��@�°~��
>�a7J۠���H��#�#ڱp���6J�S��熰�6��L���vF�.su�F'���w��*ظ6��u1tᗹ�j j��Fs9�@�M$�����7ISEY ~EK�;�)[��fjb�	N�4�2~���Z�އ���H��dІ�.U���<�uL��b<͖��H�Y��I�q_Q?�J�vg.����_|�sn��-3]ڟ؇kfd���:cq�qir�#*������|��L�8� QE�}]�ZIM;Tu����t[E����2����p����(����[�4{���ue-̭D�cDX��.��X�Z�xw��V�Y�^*�D--631�&�:R�fl,E�2���ڶ��!Ų�4�Q�2��qQ
�J��K6�K{��/�୨e��F�e�3�5w�� �r9B��%��q5j�����9��nBUI���`BU��d��zl�l�u %�Vܺy�F�O��B��Â�PG��GaiC7��j����[I�M��ŉ��bj2��Ԃ}h͝�AC�"��$�J�ȠD,�Hkd�ڤ��{��"��*j����/ѷ�;CN-2�򏷾�ZC�QL��ٰ^Z��q��{���j��������X
>�Q ]w�!8��������p��T���S�NGa�Ŏ:���.��-��j��T�W]h��h7��ؖ�؋X�D����.�$|\�������N��@0���y
�}�f[��/�{z�x��R`�'�
T�&4������Se��0���%y �ݜ%�����>�~LY�M�o[@"�<R9�3�ҫGD2vvL��nԬ�-�����Vp�#�R��:�O������~K�mM/G�$_��-�"���3�b���/5.����M�s��1ϓ�h�S���B��z���#\׊2�N�'M�N/��Y��A$�b9}��B̉&� ^)���.��p0��q�RR��+��)�&-��8ڔԿ�[�����y�0\R{��4���=O���ц~���X)��g�O)��T�'
0"�fy�o�dZ*_�z����sN�ː�Tu<��D�I�D\�ھLz���5�j�3����?�sJ��7��uD@E3��Z-��dM�/Apu@��^ϝ��L�i� <i���!D`N�pu�j�] S/ޝ�����P�����[(�ټ��L���E{%oԻ����q��R��D �\���ڢj��j���R�Dj��=0d@�/)0�3OI��~(����T��T�DD�LGXxxԗM���9�l��&�&n$#F:�j�%Fg7DANy����}�ӗ�Y�م
��C���=~����e�q�4�J׋�����S��3C0N��f��b�H�A4�=���a��D7�d��D��@X@�U2n�tn���b*��a̧�����)��O�Oe|rӡ��sV��u�+=e%J���3!?�$;梵)..���o��X&��c2#�����ǟ]��j�����y�ơ.��	�F�3��C���r��;�8W�g�@��j��)�9x��g�S`&f��$�]�����\랲�@���+:�p�[x>+=�qk~��9l'��E��Q,�&p��+��@��R�Q]�4�+��o����ޕW��wȲ-Ұ�e��ӝJ�; ��A��م�Y�o�؍;e37˄���G���_�x�s������tɰ?g�D�u@�o���b��}�Bs�?�R8n�������aX@�l����M�O�|A�4kovz�_dy����9i�cGa�{�'��Q�c�]e@�	W��e6�@@eҌ��)2�c��E��zc�<�aX����tR��/����$Դ���z��b�� �ё�uL�t�.ެd�/ �YB�&����NZ��w I��]���n&�a�ߕ�������g?#��{�������/�5��}� �>�nm��<^�H�~�t�>~��0��� ?��2��|?&�溲����P컐S�/��G�Sg���ݮ�������΅�t)��y��D�kˉ@������5��9?�`�C�0�-�,^��0\Q���O��(�;�ܟ�v�\�$Nu ��@���� �smL�5Z}��brˡ�����+��r��s�y��-7���X\#�qYޟ���AX�����L<4��.�=M�����F�e,m8	۞!:��
�-���H-�t�gq+х3��:nޓ��G���\�~��散����]1�G�����7XˆM�{vjN&��E>]�G� �C�8�l�6;��oB���r�q5؏H���Y_������'ʿ|48^��nI�&���Vn[���@�a������-�[�!��3��c�+*�I�+����� ��d���\
$��Pvg𹄦�~1����a>���B��7ČO�Ы{a清t�?^�g,iN��>�Mm���q�z��s��SeG�Mn<#��?�t����TYN��d� d�2��jmA�{��"�ӈ��� �揈PN?K(�}bϤV�$�=o~9-6ٰ�m�,�Ҧ��.6��!B!3��^�"�ȸE$������C�\g�5�`��
�K���~��50�䄬F5ߋ��8=r%f��3OG=�M�Jڿ�������1�g����ASm@~�U�
�\�	���d�C����w��$f�����չ_r�K�%��d�&_��\�n�%��N�s�7p��3��%fP�qKg�=;Ү�ᔓ[�A,�qA尾����5T��yI�ƒ*\��,z���_���~8��� h� ���+G�����𶚞����`o�>���C@D�w�@����u�����+)j������'����ȟ������w�n7�_������L
�@;��o��7����{�M]�κ� �P�ǝW�95���I�4B���3?��sl_��-��㈗��ͯ�2�܆�i ��w�O��	TC�@�g�8���a9d����Z��Ƣ�of��5���~Tn5Э8��5}�(D�J7�+o���g���w�h�&l��S*|�_�V#E3ZD#{��iS�4[�A�?�\^ћ�0�z��[ad,��d^�W�h��4��5�F��&��k-�0�9k��l�0r����?ѽh!����ÔRf���=ڥ4-��iMF*Ai�s6�Q�[��~�Q;�[;�rt6���UtI�e�}��TYY�n��.E�g�5&�SeY)<�Z�bY1����+<����uMV�y/#DO�T��4���ߑ�僝��;E�k5�>F�"�}�3���s7���׿�����
�_�Sb
���ã��i��Lq����;x�=k�Շ�4d�8��3����#!EG"k��YF�8�'mAw��m
��Y,���D�ښxTt�0�pr�܁�z{7]� ���Zy�4�V��̙V�[G���#^܏c��e�~��^���|�տ�h��<�U�F4G8Ty�%C	�0�H���T�(�}P=�$
�&F�MXGc�|q�����۴�ړ1IZ����-īQ���h�P���H�o.|{���m�V�I�`5If������ۿ
�2�$��6Z�{�$�i��o�Ο����<181�Hk�@5@�ie�Au0���v���w_��up1����S�j*�Z�X��S����\�p|/08�R�JX�,��������~2���x2�vWR݄�SPLM+��w����pe'-])���c��(��n�$Z����M�A<��L�4����5�1��v]y��&'ө�ڧ�Q�0m��?���R�d���l�&Mo��̙�;�3z'ϗc�4�_�l0@��7�")"��֜�|�I���?���|�����qg� `dў=��ξ��z?_]�  f�34�*B�����V[?���0�"����J��)#�c�ۊ�kXk��ا���a�:�s�k��ö���7e��3s��jo�y^�6�cs���05e[���oZ�N7c�)��#.�]���NG+���D$�2�畷�	�b��y�Gcv�2_��|���r�rpd4XX�d�#Vc�u�pk����	3҉�`�	��漍e<(�~�=E�ϊ��;8�m9�7�ڴ������\��OK�t2��P7���S�ƿ4���d=�����<q,��ۏ�2^��a7^���亙}�АV���0��C�d��-^O�~�+�_�g�?�Ȼ+��5��L�D)�Gn0�?�����;paP�p�W)�h��)��Ly���z�*��̝n��Bv}�����+Ӵ0��u^��ـL�H�XعL�#��+�_����{�*<˔І����g��w<�9'��Y �-�j��f�4V�7������+5�eh �&�BWg�R�4Q�߉�U<��O��}�z,�8��WG��0���>�n������f�ub�>�d�6�YE���:'ґLؼ��<9��ge�K�.ͯ<`��|�� ��N����ޘӄ�c����=<|����O'0�i&�;y>�5.�ܲ\��N��ޤ�y�qa-�Һ�.Z�uh���=r���X3��	~�/M{{4<�gw���N�S�jԓ��k�VQV�76�+��\3�@"�C���$�]Xp���t�/Ҍr��{=`�Rؖ�IV� �Dm��=�П�G��W`|D&a���M�?��{���13�-*�����L����A՚��Z�JQJ�⳺�8S�Ʀ�P�?����od��<�UWt�!1e[�Ԃ�*߄��_����}�2�u&ck���ߟ�q��0��M�2�����/�!��HO�.y�S'�2/�*��7{HZz���i8�F޻�೔��:v��ˬ?ł�^ϙ~��W˲�c^l�0�4r��-tX�}*��&J5>�@�Z8ԕ��f �y>aG"=Pl�Vp��^���B�k��Q<'m@�����0��������^zu��~��U!pw�t�2�zT��p��kҩs9�6p�G���Ԏv<������Zf� �^���/5O��Αw���7�g8��o\Յ���.ո����a|��R &H#�n����b���	�Qu���RYu���E�->i�s���Z���u�i�Gnz�{3���v��a���*��y���O�����!@�Y�����2^��J���5�9^��!�^ѹ+�.o�ǟ����a�x��
��YX��qG6n��v;F �D�(�1�=-,���Ş	���Ƥژ���f�	�x�j�{�/up濳�ڴ+9�!��c{��z�X��.��{)}@�E�IY1�<R �=l��e;k���:y��.�����]�KП�S�m�[��3�����IR��o�YA�J��8����롷��S���{�`ꁳ�Q��'��I��?�eɅ��tPCشomT��;v�5	7�7Q#�T�vm����d�
K�(3��l�����69�Y��7�5��
i��v,��u�1��:R .T��<g<]v�6j�xZ�I�=�y�ҿ�בj���n�����?�
M��oIjA\�cZ��^L)�_�/���ҳ���f���w<��n�qR ��hq�d����%UJ5���d��i6Gѐ9#?�a�ΓKU�z�'�3$6Y�L�$�]�aNc�|3-����b7�="�+1b!��Dz�hq�>��y�r�Yn$壻Fh�3L����#;��F����8�4����X5� ���()����+
(Rt.Q��I���𰯳�̳�IƮ&�+e��&�zb:�el��,bq|hU��[��S����6&����r������b����y����iP�فQ�n�	`C+�Ӑ�O�����B���$�p�M����q�}����r�q�A�G�J�*1!&`#v�$�4b[-
	����0[���>D09#ߗ��g�n�!#@��d��M�Mx�w��������?]�pG��C�~�C �{]'F�Ah}>OZGH�~m�#,��;3U��vJ)Rg�j�-Կ���ʾ�tʿO~�s�=��������l�OCNŇ�,g��l��5�KoM�v:-��1o�#��������a&?�m7�9B3���ٞ� C��3�$�E༚#�q��I�pb[��|����4�;8�"���@?�6T{2������e�h�7���3o�Mr��/�Y���-��-���M���u[;�,�K�( �5���-X��9�l�ݎB�-�	�ڄ��g��'.&� ��uz�@�[���~���G��u�|-�A%���ܪ�����g~{7��H2eM�j�;�����~sU�i_�	$�A��]g���b#*�[���>ph������Z�J܉�j��"h	���׆N�E��Đv�}aH�[s�r+��g�@:֤!׍�Fg�튋�]}�	<��ԍX�1���S�����Bk��VbN�F�I��D����l�W�T�
`��kD/�y�I��#�Ř��y��*pi�y���?0�B�h���ri����Ovs� ���Ӗ���yͭ`m5��ƹ�m ���U�� �ߖF0"}%�'���|W��\��e<�8�w��t�+���T��]�Դ-��Cۗ����;�Όf�kw��'X�nY��A�=goԽ�5�2�}6�(�ǣ�䚜�x�G�ZK{K�"����6m	$4��i�$� 9��hua>��q��or�cě3Z��_������Ȉ̩�5��p�"M�L ��yN����9�@���f����?�䝛���[�l� �����
&��N�e�d43O+� yD[��}�p88��rG�A��$���rY�n����Y#�&��K
�_��#�k�6D"��������9�1�W��xy�}����B+㳛=����P���4�������7�AO��%WVs��������Д�N�]W�=�6�b����>��؈T�\"mi���ūck���I�Q,$i�
�D�oS�6!�7����rޜ�����Nz��xz���I�t�o$i\�b	]����ψ��$Y�c�i8ײ�Čeg��1���D�9*���M[2��K��;�B-�D��{����cwW:AJK�uwf���8��Z~$�i��a�ᖐ{=�'.���Mo�����9w�4�E=,b5i�ʜQ9�聐]@��;�]��$s5�p���l�F�����S���o���][c��Y+TWZ�<���q$g�Y(�Ɗ*U���y���!�X4>�/b�IŔ��~�fxalZ�_��ҩ�̍�˕2��\q��<d�Nj�1 �[�w<vw�����aMt�w٦b�y�+���w�K1^����1�+��u���f��V�A���O8�_ǜ3��<ڸ(K:��`u�3�+<�����(W���v�h&F�����3��#���`�c�l��Q�g@B�a��}+Q,����W"k���01>��a�tϭ�������K�*���4A	Z���&���6M�v�6��J\�|>�_�¦��9�Z9aB���h�)�;����V��	��>�T�x���^�H�Og	d��Ya�:���������7�ʊ���*�c�����z���]ܗ�2�9�ė�frF#���-L垥O�\x��;)=U�蓲e�7˛�ӏ��^��<�����+��|7�҂� N���F��¯�=�H�	~	a�͕�,n᢮]ޭ���i.���3�
A(�N�y|�m�/)�AHX���Y��+���cg�\�N��P��쥟
�Fxh��rsZڻd�'���Y���������1aʶN�N9��F �u����b!v��[����I�F�e�O�����ȋjE��+ �DBJz�'�u���]�SD�׿f[�1O��va�h�����T����F�$
l�w��1�B��i˷���k�(�*�km����cTF��7���]u���αY;wR�7O����wӐ��V�i��t�(��\+��]⥫��M�zcx�\*7A��k���[9*(�p���/�7����b��y�=}� rB�2�mD��B�k8�{a���g�/�S�i«'f�r4a��:>ύ⫗��>����c!��K)y��
��q��������R@���/Z]�<�G�x�<O|Ud�|`��Rz�������C�=��"v���;)�c���h�.���pݼ8j���-D�l�4Z�q�����d�Ǔ�,��@z�JlQI#�}�>3��s�
��g9��T��\ �c1��@��o�G�<�0���c8�8�u	�E���I FM��;o>�IvC�Ӵ bcI�%�L�j�x/�i��	������ʛ̝.���'�ɞ����U�ݸ�K��Th��8
%��ʌ�������^'ڽ/�bLx%�^�+
��m��9�6~^���q�Ժ2˷�djh
��D1f�P��1������ݜ�p؁�{>&ݺ���E��g ����DXL ��ͨ���!��Y�昸�U�����A,Μ!��	���jd݈�X.��w\�w��y��^eg��7o�D��S�g�ͳL?��z�?�>��g�L��N��� \`�A��h	�,�\�Go��w[�l�� %�BT�����XbQ�XS	;w����UH6����G��&.z�<N&g��M-��zT
ˆF��wy�L�2��kV��'����LMK�^�'���nY�J��p�!��q ���΁D��j�_�n?���t;`��"��"	��40��]���N�e1��2.����T����]5�?B9�aJ�+�MXr���A�it;fr���ƨB�+e<{ފ쳐 EҀ[	�I�����w�5�y��㚊�����b�����{�xy���{�-K�ϋ*a�dGm��vc��Xx!u�5QT1��d�'0]M�&Y.,,ve�gp?B�t�f�Sa6���i��9#�" �z�siV��1*�Z�t�2�e�w������~+�{wJ?�}�����g�T��u��k6�s��g�o�
��
B`צ:;H��#A�ˮ��kj1�rU%��M�1Y�ZE�z�嬯�1I��w�������j>&��&�����)<��f[J
kZ2�n͙�0���J��f	�)�\���vO#�񮻣�dc@������mʆI]JE��ɹyy�(��-�1W�7�~��T u���}�ލ�4?M�Bt�ܥ��o�"� �3[�8|��I�쾼?���q�볘�:|�ć�q@���8�M����C �I�]��L��`.�	���W�;sw�xO�1~���5��ɴWҟCVM���A���/F5:�{d�qz�l��\�0`����Cr�ˬ��7�)
t�̱��ț���#�g�`��CŨ�փ��2��6z%ڣ蚑8}�-�0`2z�K컅��Aԯ�śyCk0�b��'�`/^�@�C�؅Tqb�VE��zJ'���Օ�Ȑ�<E0��A��N�s.z^�6���-��!�'�H͘䭾Xy�#���E�*�}s<n����s( �I���i2G�2�̨わ�Q�j@�������?�o�K��I�R٭P*O�]�����0	� )�X�F���.tN;�\z/���~t
��M�f��$J�K4Ք*�|~U�G�6��z��|1>?����G���ٹ��-iH��3sw7x�������c�y8�B��1�0�Å��C�=Dd����k�t���w��2����מ3�����Ĺ�4#��"�V�;@�a%4F��\3����d#��a>�?���Hk���e���dR��a ٗ`�=+�!f|�y���zԓ(��U���qǷ[���)�8�e+�H'�/ؕ%�+]�mq���,<䧄1|7�7:���*�h�n�ѩUw�f�(��L��bH�J^�2'N��S�T��)����/@�Ĥ��<R����/�+n^�!N���K��u�s�ƕ-�"��l/#PoK6���~�ߌ���.�KI`�`���;(��f�����6���ܛ'�y��p
�0��:��ɗ�E�����L���Rũ;#�� �F�*B�6� ��Oj�3M����K�l9�R��
,/ )�`�8�A�q�$&k��*O�Yt�v.
�^6��i�I�m{
3����nQ��*��ة[���T��s�0���O�RЂu�D�`�Nf���e�#�)�l�;�g� ���8�:�o˟X'j��l��Fc7>щm������ƶm6�Olk���ܙ���y?{������p��}�O[����J���R����]!�nZ�� <��y�ˣ���B]���w?H��[����*,�k�?�hw�I�5+��Z#��n�dED��5�����v�OU��8� ���d���f�IPα�@h�L��~B׶��um�~��}<�sK��if�~�T»��f���\��.���!��w\L)�s}iX..�
J��p	��)<_	��;-�~����.'���K�!@��1n	�Ɔ���Qf�� >���&�\�I��q��>�W���/�a/��ݮ�qr|�}�hL��0��(�D��S9�b�?��9B�㙜��R���E������81�zd$��Ѧ]AL��������c��Z9�����;Q�c�Y��)m�7�T8�v��Z�DA���J���C�^�}������s�JpLj❬w(dg���.X2�x��D;��$X�EL�v����D����. �W�Gט��t���"�^7�����:�߷䳂I8B�"�aZP'��E뛲�	�c�g)������*}���z�ܢ�[o
�X�n�n?����*p ��)Nl?��%�J�h��uN�;�t:^.�ө��j���֚t�j!G|�3:c��/�b�|��TX��4��� �]��s��I����:�*7��8/:�
���S��Y�y�SR����H��b�؜�$�W�����B"%�!����KP���ul��~ڋk�\��<W�}��Iq��	����oCs�swؖ��tqP	=�A0�9�jt[.��bC;�?B-�7���q����7�����^��D�'`�icf`���pW�O`0�a0c��������p4�
�q��{�{�b.~`��q��.�Q?݅O'��jw&"����2�5��֒�����r׺:�ZPg���-#s14R��H?71Ӝ���͠����6.�)��j�{�E(��ف���}�榅���)�rZ�l�3g�:"PJ#�Zs{qn�Ѩ�T 
N����/�q�l"�3e,4�|'T�++�_����^o�N��$״O���Õt!�Y��Ǌ=���x\Sob�+񟇍:+�^Lg�e�\��
����T�-�AH��͕8�鵔'r�������~��M�?��)xN�(��II��z)��9#77P��4����Qŝ�a�`7ee�+{�Ic��R��s�9�b�nJ���{����y3��������%�$�|����"�� �N��W�;]�w��T��V/�Ρ���aM�};N���6\���Tܦ<|��|?����nwGz��Ί��Z�ot4��/ G�����{��JΣ*i��A\�X���Op�'S� ����n��M�������#��UIJ�e����QBF�`�U|/�M1������y��O�^Q �����$�(����D���.GV/�`�M�uPb*��.T/�Ҳ,�t��X�ʹhZV:�t-ҕ��" Z���!o��X�N�\��`��	i&R-�VǁO�+��+�o7.*�y�A�^��J�F �����3w�8�l7υ����o��KhJ�|{�����]V�`(�>_��TC��w�/�k��,�z��
��'�j|DMe��a	&��3;V��$�㋩����u8f5�$9���ݳu�}f�/ӨE!g�g��uG���$�+�Id�߶�Jg���یTƘ�s)eg�	�]^e�ݖ��|s�L,�����/OU���Ϫ]�ם�ˡ̇��i����)�@g��� ��0Ũ�v>�[�������b���$�LF�ʬ�������;xI���O	ϥ�,�o$�ā@A<��.��<��@�<~Gq��sx�&>$�[�N#��@y�z�H_�����F�|�w����wà�Î��w� �YFv�ACz���&ޏ��R(g��x�	�Gqr�y�VV'��5�6�T���v/��/��V�O��6����W4��_�%"��:��F?�u����s�9Yo'�Øfr���P�Y1�h���pi�P�G�'��CF
�A9�ɺ2.�ƛ\�}�+�;a���F��}�K���p��MlQn�j7u��|����AN�q����(:s�*�(yr���n�ڠ�
��)Z�m�Ȇz�L-S\�YS�\�\�l�q��)݋��P�9�A�a�mN4L/�GQ�v(�d9������(�=L9��W$��Q~ȭ���:�6a��S��i>p֕��r�02.]ќt24��s�ӎn}�:������;�M"բh��(o������Ә��fF��y�K} �5��>ɨ�~"���u	1�2�߶������cz�gf�2�=��>�<4W���
��L�ǚ�����~�\J������_�*p��2�Vq\`r�q.	��}h��ȇ���8|-��˴�SO��M�d����6:��o��(��Jno��>��6l�w;;��,O,xK=g3l��M/,��e�i9�%��j�~�nO7z��N��޷%����t��^�ׯ��n�aHf%�
o�"�����0A@�8��Q���)Y	 �k����#��@)#�
��Tޙ����C1,b�K����هϗM�ȡ5��"32�b���X(�<Z􌾪0rO"\��U<��5���@ŉ��ݨw��'yZ��w�5�\4yC/?������S��-��mp �aF�g���^�����1���=��e�gR*�^��c��zyQ�w��Q\Q�!�{G4�D2n;�����
���h�yD�F���j�}H��s
�1�����C?���#"�I.W��N�@�\� A�1���չ�Y�0��ϵ
�6�h���9��^�|�d٨�t!��d�}=n�f�+��={?%�Ϗ�Q�[�n%]8^s䆻[�%�Y �����K����<����șפ�K_Mc����eW]V5"J��`-\[�*�f��(���I�McOr����V*�kO�S��Yԙ�.3� wu��;D��pHX�ϩ_i���G������)$����?��b�|ue��J��% ϙ��[�w*�jp �8�� 3 :ܜ�rX���\ۆCm���2�����2�ZJ�.sr���
yS�F�}c�B�U�O�j�)ם� ��1����|��YLE:[#z6P�?Ya@���-*,�/B:�_ӎ��|��Op�S��Y�B�3����$~�<MHKRV���%�o�� ����v�Px?H0Ak���W��e�����3�s]}�
��z�~I7<��na�8���p�3����Ɠ��+̡f?Lބ�"PV�aR���ı[�v6�zGC�]��|�g ���*��9 �N��P������OG��0���Sj��/2k��5|�����*SE"�y��'KPdZ訙�6&0���	z��EP�q���Ù���\���-�'�RK��O���F�X]�R�-���̋���G�g�?�P���Ӷ�$��_8�GEσ����;����v�Z�N��`��T���oZ�y~����\����ͫ=;��)ťx��z:�`j�l�B������q�V7�Q�2���;{�S@7��)�~rn�P��l)d�/_Ӵ����x!��YݩV1*�z��NB>c�VS)tfNF΢DkG���}��p��H$4X(���4�7H�ٳk��p�g���_a�e;é�D�K�ph�-P�qB���'X0#�Tp}g��K�bq�����A��7Y��luأU=��{W��`~ų"$a���c����2<1�.�=�RS�&���!�����%*-?�a2�wy�RKFv�]_/ J_���?U�B�]�,�Y�E�	ۣ��0ޗ����e|7�>�ShA:[v�V��x&w4���k���u�d�oO��xY&�6��i;}3E��<y�_�]��� F#�v~T�m7޿�U����n��?B����͝D:H�_�X�3��Ga�`������N��c�L,}H_�^�>���)�8kz��|8e�_����c�Wf��)��ߓ�S�����.���!~���7�+�qc��;l�8�N�0(��S�O�b�ر_h��D�j�����Rf6Z�����
�j޿��n�=&���%-D[�S3�U(��莌�����ϊ��#9�F;~�!��c�¬�%�Jф�N��j�Z�E���XT F|���׍]0D~_o��$��^^.F5�cE7�g�mz�QS��{��(�_̅�-
�ų�Fa#=��hM��w�D^��p���:��G�@��$p.��_�I��{��=�y0�{�����ɋ��k�D�ɖ�܄^z��M �5(�ċ��w��r�ci�k��-s<��;5A$k˚�]�ݧV��9<u�ܣ<j��b�������ͭ���0��ҕ�>fl�ņv�M��@L7��1
��ahҭ�NfuDXtT%�hC$�`?�s$�R�1ϒKa�����H�����;��8ӄlg���-�g�w�>�Qb��i��Z+�����t�O����ך\���1[�Sl�s��rm2&��rE����p�m��O�y����u��YD}�h߿�	mlu�՜�q`5�v��R��$E��$5�K�{Eqg;��%��	�u�[&��Xw���ġ]V�t�T��-�o�����I���rf����:v�L�|��kT�+e�! N���Nu9�7t�u�D
OHS�SS;�O � ����f6�K�b�e�0�_4�z1��+Z�gT̂7(�(�[�t5kמp6,@k+�Ҕ=&�#Z�Eo�/�ã}��م	�;|M�U�����{�ʇ�i���t�c�`o3�5���]Dٵ+���8����VCj�ŧ%������*���#&�^�ů�-
?29�m��8S���r�F�:�V	3�^-9����k���Y�eq�^b$��I����tl�$d'��8ro(Dbh���lZ����O�e���:ϰ����(��{D�È%�e�9p�u��"q���쾖��&_���"/Z�L=-��H^�[Q���N�0�r�d������"�F[����M��[nut�5���`oM�ۺ0^U�L��,=+o�e��u�nn��T_����Lݛv�lݝ������7�t1;:(ߌY�S��#G���]l���%���8}���H����!>�Rݦ��a��+�����8T�h���G) y�@.��r+S�4d[d�0�ѝ���[�)jPόO4^&Ʊ�֮dړ"����_���D_����'�Q�?eH�]�4���z;�j����"7o�.�PS��7r���?P9�:�$��i4�;��3��~�Ž�.��N��a�O�(��>p⿧��8C	�vs��0�͔�G?ܭ��m��;9#u�z��8"�3�-x_����a�9��J9ęEb�"��y.��m��DO'w{XG,��>.;�		(�uI��Ť}>��l3|(8��%[�O�	F]z�J&�j�|e^J�F�|υN��Qp�7���|ͤ%!�F��8�_9b;g�v������i�s|�3��h����ߚ�^�?�C0qB���)f*w%#��ޗs��H���؁X%=��P�r��˦�W.��2�x��fr5�wD�n�w?�h�`q�4d����FFZT;�h�U\[(��O�3�үF4&e A�\���(��|�2>;�-��g3���E��Y�'�	���li+�&X���q5�}v4�ц���lP$	�r�~�|�"��؀�-.M>GY��������q��XT�Aԍe���*�������!�,�p�"�eX��Ȣῡ;�R1�>�.��l2K���U7*
��Gâ1�*x��*D^>���p�CR�ґ�#�'��F��U��lG��W���8����ž��a����=�_�e�@���U��%��I�yh����t��_��3�΁���̑s�>�*M?+¸��A��5�{8!|.+��c�`�E��� B���Wo�M\�M�"�.���+��z| G/?��#)uvEpw�`2��s*7�ݟE� �]Ν��#�a>���0��K�	�h��jR�
3ok�����T~ �� ��Zo�|?������j���#کf�t���	���kؗ��p�o _�R�F������)alV���F7fs1���o<�آ%GM��7E�ˬ���(��i��1Y(�s�q�˓<��_��JG o�Ak���8ҥ�a�&?��=�و��!�	2���,	����F�[ri����m�v��AC���%ʦb�6��~�p� R�� ��#''��J�J+�ʍ����f�Aך���U�"��u!�����5��^��&���~an�����q!�yQ������܁�_LB7�X��U�����VJV2yL�����ǌ
��Xװk8gC�ީ��&*�ݝ��&�<zZ�� G0�����:����&�����]<��U!��}nm$d*"���/6>�yK��Ǻ���Q�tr��_g�k���\ʒT^���қ^���ºO�݅�턚1�הz�)�n�2o�m�
��j/i;�^�%3"�� m�YٞK2�1c㽾�Q3��+	��	��,Х��ы��`>|J��6k�ϡz�;��t1�0��W77�!Dg��d��S�͛�j�	eG~���o�r��$�F�j�����d"�%���Ѡ��_0x�Om�rLй�:}e���I���=�k����.S�vx/r7��0��_>��,���=�5�*�sDM!GZûAS�a�_�:@���byE��#��m]��]��VrG�ɘ���4s��"q���a�te6��3��;8f?C�pE�|�n��I�*��D|�l�$�aӌI�ē:����W�������ɼ��MlzR�\P��<�6���[5M��н� K��T��.G�C������hQ ���k�t-&	��(���c��i�:��!�`�H����: +b�p/3�B�j2���)u ��n��8�!��]�2�kf�;*s�G��E �KN�F�.�̐ރ=1�[M�83zŷ��޶�b}� {���I���ԧ�ڎZ ��xs=8�v��}_v��Cߠ`1��G�"�E=����A[����O���B�n@F,vj�Ir�{y'W}y0X~��O�$�ךw�~2y���9êf#'��f��llcQJ�K�pn���7�FTt�_�4��D׾�
�I�~��W{C�_��C���Z�����%C(	k�'�H 噯��g�i ��~}k�r��>+*�ѣ6{��
���祌^�Oq|+�:��˻��� ���P�K��T��Z�v�Ak��N>�=��;�FA�rز�-�G${��ݨ7U�2��gpƉ
鎕yC��gpU��(�bQ�vh�)��]S�Q�q�q��^�g����$�Б\�����ʹ�/6�,(L��Gk�I�8�ފ���)������y!�/�@}��(O���QO�X��	����q�yf).�{���"P�G���>��$7�6%NND'GH��\D!^��rJ;2�nn~/~_�R.�TVx_b懙���/zH���B��==�H�띙ڶ)�`_jQ-�w�hz������UU�����_THz#hXw��=�d^�2�?�oх+�O��=�1��P%���:<N������zzVk>�y�Z�^V�����a!6�Y>vwl�գ�;*�i��o�V�'?Uw>��+*�9�7�^6�-� ���ΜUN)>b�Z���ہ��7}��m�R�+<�6�1~���_��������t��'i�\���VFCm�-&�A�@���%��6_G��c�!F�s�9^��eU�!-w���������dn��S�R�����B~���!����4��y�B��C�x���|�#R�ݔ��J�A�� �}��A��yMn�Ħ!����`%F��Xǡ=�'�W_�A'B�"����P�N�*k�J���:Y�@���X�w��Nl����zw��]"���~���ӘnR�5���������Zɉ�q�ŀ���͂fƍ��n�����K��k�+_�e���������Ds r����`Q��{N;g5�ϐz�-UK��i�iKJIj�XA&$])~!i; ����-�[���}ۇ�����,�$��u��+�� |@n�x��r:�4N�S���>��Ʌgu}��]p��XL���C_h�H�?T+��7��2x��d�l`��I���=����z��غp�v?�������b����B�Wp'S̟���ch�m�#���Ѝ$՝��I�{L�M>�������T�Y�ۢ�v�T�Q4lg= :���Y�U�E��A��7�،�C����ݴ�o0+�M��r���A9&=��nw��H��Q��G<�7R��2w*��$g���{�|MK��f���l����<M�-�>���T���%�]�Zu�F������EH� +`8�U�'��E8��G����#ȍ���+�E��0`�"@��H�1^���"|MȖ����w3���z�J�_��&���PQ���YE}iED�����"T��̎��
J�"�tKV�j�b9QSq�uO���G
�΁�5�U{���j�{�	�zآm�a`�m��#�

�r��������]&;���@Q� (����~e�4��Kc�S�f����a�?s�O��ڲ� �f�	�)p3���v�ƫX�$W�W����ռ��6�A]%.�h�X�v��8��-�s����7y-�y���k�G��J�S@�j���l���,�@0�8_n
Bg�إ���ӛz���\�ECnH��5l;�<!'��V�+�Uwlo~�@���p�υ"����E�l�;��0�E D@[x�AΗ��IC���D8?Bz� J,����1�4�^�"	3�S-Jf���$��<����.���=����)p��μl�E��9���|k��Z�d��� q�X;�����F��/�O��*��36f�5�Ї��h|������x�����B4��hb�F�
_�p�52�B��'��m��U��7�����Ǐ��(6d�_>I?�5ړqa%�+��64��wQF<��.&2?^�Π�(1F�Ӯ��7m�X*����!�<J��i����kzg	IHRNQ�O�z	+���$?-���֑�\2զ���\B��A!��C7i�x���ɘh���?NZ0����#�vh@��8�Zwdn�un�n��m�zx�R\�ĐC�d�
��lm]��9����0��dȧ	M5��]�j�]IgHn�Ą���)Ȝ��x�	GYy�}��|ϑyo��܃�v�Ee�nN�z���:���;�u��+Ҿ������6�C�MHwO'
`�C�q�p�	o���O����e)�0�/�A.Z��{�`%(���D�0�D���ۤN_�6)�̠�`W�6����ti��3���F��I��k{쩏�Ύ��|�/7Ob�@����P(we�nH��KMi-`���2��R�'0�w�,����8iՈ���I>�;��{$����e���n�t�P�1l���(�â�Q,B�Y��.���Z��д���+9�~	��L�4�{{�d��������䔮a����,�`�y�ε���b�"���Rcv�jd
iR|����eY�)���=*���#�A.����븗vۻ^����K�-���f��}{+�ʘ� N&TO��{)9��i�Ҥ��@E���n��Q�4�㢦ܺ������88`/
�Uv2����x�:��n�J�V���v��n.��%��^�ʴ�p.��,�w���%2���̞�׎Y>��kq��4&k��-���&n�3�l�M�O33������T%8��k/� ޢ�m6��rD�2H������'�2��yX��N6-��BwrC��K�� �3c���A|:��J0z)N��p�B,��W�B(�/���)<��)���w\�!�	�
`�[�P��:����j(�,�{$2Y��<����{lLmji�k�/&����U����Ĳ#L����),�<_4@Ti.��N)���e��=nĞ�~x"	���`��U��~����z�U�`7�U���Q���W�������z�g>��,����Z�ZgCuU�?rIm�F�2C��r%�ӸW��1����S�1��o��&��Lk ,��;���Mz�!y��}ҽ��p.�O·�7�9����l*�3��8?,k�*"��7NB��^V=m��.p�'	Kmx��qR��q��U�|{ӈ-M�&���-��F��<����qe�#R`�$��mc},�lu�~@��p�A�8߃��SmƱ)q�eQ�K@��G�
�ۚ�PʒAG��AD~T�Ӄ{�7��+��d(�"�WT�\e�a���+��ZQ��̬l��L���v+��@�eC!�q0����c���C}twB�&�L�]�dg�_T���ڇ$^ jg���}?����ލ����Ŀ�dЙ���#s���R��\ئR�o�a��& ��!D������
��Õ_�?���uو�����m"�'4�"~ͷ�X�i�5��,�[����S����HQG�Nݢ�l�n鬩J�I��B)$�C"��P|$�x���O��DB�j��� @����u���s�Uش)��݊�����7��L��t�~m�s�V�,�9͝%bб:E��r��S���P7}�W��Lb#¬dc����3E ���W�����;5��W�cz Ihl�� J�R	5�ν��\rc?;�d��gnWH��C�H��4[���I�|��\��m��v����sS�����D3�0_��J1n,���R�Q��<�s���^��O�$�_��T�34�8a�
���7 ����V[�/����� �������aRg��)Vce���A����3�[�w��LR%OA����$��D��Yi�FM�����@ߨ��㷟t�r�lx?�1{�@*a̔��T�;��_�%��{y�jb�����⬗�?�W�J�^\s;Ũ���^�=:�a�`*&��i/l�ˑ�:�g���]�`��������2��K�_�_
�ĴW3��Y�$�P���� �.7�|70s�����rP0�����ō��A�����m�&$��&�$!ߞ��p��o]�n{C��@`��*�[�e\-���H���;V�
�w+��=Fl������nQCNR��bHALqx&�8�R���	g�L6z�]P7D�H$��xx�	��AM��Hx��Q����5bgK�:9jL��ݍ�ߴ ��a~��B�n>I��?1�g�y�瞖K'�^��k�E�z�$F,ӟ�exI����1�2��������U�z����q
a��?������n�^��RK�|Y����mK:��:
p�-P^���-�I6f����`���o�MÌQ�6jZ:|���A��KM=q?�?�tq�hS�RT��$��|c�� ��]݈2Rg��앒&�ۏ Ag� Ò4���M)���qK���N#�k`޳o_�����2�ʙ�-����s5R�%u��iB#R�JU�	�2��	ݡ���/e��];>D����Z���Y�����%�+I`n�����7o��_���L[��i�Q��@�M`fe���_Hm'rΕ�P���B=!�CQwJFT�|/6����0���z����`�G�������{-&���4t���A��.�!
�B!�(���~�2ivb�%]�(&o��)J��pZ�9����ȗ)����=�+�2�W���'���ҨSŔ�`f�_��8�S������M��v�5�Ʋa��]V�������bO�H��c՛�ա�n�ZR�Mg0��mUX�S��"Sz#���*M-V��\�pp�q���W�?�iV,�����tG�W�t=[�8�}\HNs�	��HP��z�����}��qS�zP^�	�8V�,9�J&&pc0͓">_��)�cBʫ���V� �T^��{Q�C-x�;���f�'������2:1z�f����P܆�W�S�l,�)#����o�"�m��xq����m;p�!,�O��C��$��M���]$�8�Sp5O�1[FA�/w���y��r�eKH8|�OE��L�6&>�ѣHX/fJ
�����b���d���TIf6M��fEj�*��jf�o�� X���W$�챥U�j c���54a{F�'�`M�?�}?�t^Ϗf��T�D�ͅ�̌cCc.e�lnT��׼�|�d4ҡ
`S��添F�i�_��j�����}S�-�q��9��-�����p��v[b1}<	��u����@�I�gn�ۅ�����'yІ�s
PU�iP���Pb�l��������e߄�\�㍓�,�\ 5**���&��s�Iw�pJ�{��τ7V���y�Z�v�J�)��Bn�H6��"��&)�|�����6~���Z�m#���W��源_vL�+���7��(�.���Y�,@9Q��4HQH�ղ�TP­)7	V^`4�xb����p�y�Nk��0����h�H8E��(R����N�3JA3`�R6!O��u�J�vM��8���N�]J�%j?��W�s��ޯ!�%���q�]E���,.�XT��C��,�dy�/��� �WD�]C[��@ ��S��⩵��n��W�OAχ��
`M���O�_��S��0�
�n5	�8�.+��rܸޑ��{�PV��Z*�F�[ +�x#��؀Ys�O�Ed��0
~�6�Tlw�5�Z�'���u�h�Jکۻ�����P��l3H��Ŗ���5��RI��3�%9ST :03��? 5:�M���b��7Oy��XeE�$^���őԌ$&k��V`{��[ͨ�?l�LI\$�b�1�:1��D��E���9&�R`�P�0;	�|��<�KȬ��i��S
M��N�f��%���'��;�<�g����D,��G�J_\��N��S��V���Z��yv�Z��㐭���l�����6Q�Q��ӻ��d�u��R�i��R��ҏy�Ix�?�K�O�H�0=0�!�Փ���s&�w/JC�Mg����<݆�=�Ѩf��(]?䆮�ؽ#=�K53c0�I�Z��(N���J���T����b��罡��]����K�}3y2�BY��wCSTZ�u��|Ͷ�sZE���ۗ�0C��+1Z�uR^p�ɵ�m����}��GkW�7k���D��[g�u�.r��&jaZ�� 5o�E����}B`�����7�<�1�a��KXW�L�^��/�g�"�e }i�q'�|>�hV��<Ӧ(�w�������N�����"�a��b���!?`c��U_������ gV)���Q�{�� *�:K��Τ5�Τ��"��Vڒ��C������&������S�<BZ����N�	��kw�߫s�؃���R ��>9���+-����a�E����~�>�:W�i�h$�D�'/�le�9S�@���׫�����(�C�Y�$w�e���\���J�¾��=�3]XK�@�y�(�V�k_��#z�ɐM9�qMT�ް��d��=,WN�wќG�$��9���)�QeW�WF������h�Kcb�ЅN/�:Y���¬c��b:��T�j����ǯD�< I��8�~�I7���w>�I������k��[~F��k�.gM�LƬc�`h��V ��fO�R���/�!r�C����Bgt�v3E������S�7��-�h� ��C3:Y*I��M��c.S�z\7�6\Hh����3v���3:<�faWPQȔ����/�Z�ʒ!F�U��Z��H��^��������{#-�E8&P��H�+4��[���'+4S5����ʗ������o�3ScY� .��8N��A�n^�y<��h�k���4ݿ��1@��Z��O&f��)A^�w��g��֭
��Y�u��F���Zc�� �t�:59�{3�Sv���)��{������s���KS6�Q
�_I�e��~����D}��g�, �����5�����ԩD���P@�i��~�z3�qL����Ir#U�]�L�/�n�'f
q8k7C�j�6�
��d�p&k�fhԤ�~g��m־8����V{�7h��Q�8�*_�=����U����t�v��-a�8V�v��(�F�AA"~�����t��Z����{��K��Ym����%ND���EyX�XX��qV�����4�×}�$�� "yՖ�/�ç��y����>A�ή�c�������Ss�HU)mdSaY� V��z��=��P�՗���\2'E��l�D����a2%�Fz�o>%���=%��!�}���`v@�2��k�Q�i�2ݵ�B��\C)V&2'F�3+��.<%Z�bݭ��<n�T��fV|mM���`j� <�#Uk��E��)����TtL�O?E�A�?��^B��k����gSe̗�y��#TL).�:V�o��(1��h���}+�r,��n���������@@��M��>��F�T�����C�&������n�WJF���DV��\|��l	��0�?(�	�iJk�E���4��3CZ��඲���:��{��� &�]��t&Grf���W�V$G|��`I�މ���$D~�0���������+v
�݊:'�lM�v��Bwm!�}��^���fv�� ƺ+���[/�G�Vh�8�=�+IB_�l��zi��[Bi�.H�^����{��7��ݗ�,��io{����%tݲN����kyp�m��A�_�3	���`����� �ߥ6~~I��ϝ�p�(��:��J(؞��%=M�I9\�=�
�x8#�Sp�a�{��RT$�ؕ���ǌU&�/�]aǿߦ��7�0���+S5��=�l���m���<��@�Ь�� �;v��gE��ᬦD�L�d��C��������Y]W�̈́���Q���1VW�cR�8⦿֘ۿi����S���Cw2[s[�yw��N�?��8���n�'�����h�iA�/��*�#B��{Dwj�M5�x���JA*�	rj�����xc�/�e�O�0_������F�$l�\X��"�	�=ԇ��y�hP��]��>q�����K�ذ!W&��ƥK]��
��L%�T�Ħ�)%3\�ڠF�x�{�e*�L�	_� !&�]���:�?��w{VV���z��@\�H�H���0x":j��G���i��JB�����*��j��4Y����`����x���I~��Gy��W��k���<�^�	W
*q���^����*�:�,m)h��7O4Q�G�q��ވ�������@q��J��a��)�z�b���ņpJ������GӚ&���s��	cy�ȥn��W�< r��u<l+��+����f����]w�y4���Y)�fS�XL�Y��N"h`ҵ�LS<�q�1�,AJ��Q��m�a��j�L�ˍ���<�-0�"zF�i=&R��M��ыͷ�����US�}O@��%̸��h��o��Aʮ\�d#)F �Ǻ8d�2�~�%��'P^g'���KG6�u��=.�u;��0Nyz�_�y?��Oz}Q�^d�\����Ç�������7<���;�5�r�u�/����R��^"���F�۶�<���#�:C˾��&3���H���[��Xw�&��r�6�4�<Z�H;V�T��� 5�j>�1�6� �&����~D�*�Y8�W�\�����IY-s]4a�9H[/ZYn��eH��]�k`���j�A6�}ɡS�%,�).M��Ac��6��Zuu��EQ�J��LE�j/���� �(ʮ>7m;���f ������t�w��3�ۦ'>;�

��:�}�c�b�P�-ш��R���˄����,��k�p����^�6X:�K�S�N֔�0�`�s��P:=��4����<J�0���GC�k0O+`7=~[5P�����s�Y�5`����n�h��<X�qs�>R���oƟ�gP @��ʃ�"�
ɰ*`5�}����=��.R޴�+�Z%�m�`�V�3�jl8��2��d�~)�;9n���є7��c7���9����ވLV �4������$�Գ�G�̼���=���!�������C�|�Ŋ\�����o����b�+�֥�۶�c۶m�c����юm۶m����̹w��oճ�j-���H	߮��:�_�H�d0�{�[������D	��d��M����e<��E�����LCJݑ2Ñ�4W�JS�o��1�����S� �:�0JW�f�\��WMڭ�>�z=[��^�;���
D���0��_��S&��Ⴚ};	�dY�Rp���˪�����>��F&5)����3��:�{rx���,�㾵��aˑ��[X��J���GR���	gJ�w�j-h����.�.���E0))�⃘���B߭;�S�F����[J��E;	��H�vK�公�}�p��6>bx�
&���&�5��V�<Ft�T8jXl�~����~�35f0q��o��d����q]�H@����8k��w�R�a˗ϸ����@q�� h��D ����;T��]�A�j3�R�/�_Ft���H;󛂃8~]ߋՉ�;6�cc�c��p��魑�3̸��� e1WaV�ԅ7+Jc��Q��n�7�(�L��є����1�#,ח�\�/�g3<�~��9C4�����@ܾv�l��]�R�ED:k��,\]��@Tx���I��_�%B��ży���1~�6��>�ETlD`�'����u�udX*��*�^�XƝ>��3��H� #͊3P�O���}��
���fC�y$��� ~�?ţ���7��s:>���b���S>d�*s'��qv:$w����������<d���/ ��]��(�i��S�ZuB�fL)1�)�BQ�d��J'�k�[x�~"��N�@VnFfnyܾ��]����s�݇jk큭��r�[�S7�[�&��*u��ۘ�<�x��%�'+���5�\�)����4���zՋ�ylnԁ���߫5��������:=|,����TbL�O��]M���9��t����`��ZD��$Bi�l�}~��с%��ǝ�I�����T�(������"��@g���7/ ��p�����E*�>W�Y/d�fD�r͡��ց���Q�Ѣ. P�e����%����{אU�#y�������oRs�z�D{�	u�B�G� �)��P�9���2@/�� ���������2��%0�0%b�Z�"ۖ��(�Z"&�##����hB���tу���S�=^5��J�����s��'�Z��y
���T_m<���Y����0���04����u�4ݵ%�Q�Z�������������m\���ڝ"u���!6w��- �=M3x�Q���� `������ KB+A�&S�Uq���~�S��q�>L6 ���Fʨ����k-�#�����0��eX��+�?L�$_`e������}�Q*xV�Q�ď�M~lDD	X���5�#U�D|P�l�k�=����F��k"�&�G^��6K+t:U�_���?t%vȊض}+L�r�yg����ҦO������u�����I�
�Kh:���}b��K����%�9�3H��dJ�'�O�2��lr6?�p��5���9kY�/�����ԞZ1�����̒����2;?�� JU��_��b��h�i�������hl����C�yӺB�t�ٿ�^[��x��bT0��旪-�����"xtV K�ʳ[L�������D/�����isXv�U$H�AQ%�`-�3H�dOS,�
�D�`���an�����{L�W!Pk�"���B�.P��;�R^��'�/����%�%����(���l;�1H�)�^��6�8�U�u�Ή����e�X���y�4���ĂꝄN�� f[�)>��#��\v��?\^T?��-��C��2/?[��k��ʍ�ڻ��)�+�Q��*x֋؄�/�xo~���\Aq�12+������aĠ�G�cM�+E�Լ� 4���kiF���'a>��},���t` �i�"�/�k��!��YX@�Pgj��\���'����~Ք�m�>��G#֜�z�.0�(]�!���b�t?�F����ӎq!=���>��0��ڱ٦}_��^v�v +���K��H��Q�7P����� 
�~�9�y0��~����n[I�:�YM��� w`���/$�Kz��|*!����w���s��9����V��o�{���m]"����b釟7������I��)+�E,X8@d(�������*�z�+��m�T�5Sbi����M���պ�A:�p��l����K�!��ԛ���)�p�o��0m���2�m��v���ǅ���
���Z��c~C�Y�Ŧ�"��r]����ؽ�P������[1�琑�(�Ͳ�w�е��x��P��ֶ'.��No��[����a�-,ov5YT�vBU>�j����`���Kð�kN�Ĉ��g����N�.ݤ�/�{�7�n�C�-��{�U0�S��oi�zݰ�
E<a�u��e0A�x/~J�(n�����F@�.��m�^H��@��l�dz�4*����jj��1h���2g��b��W���g�>l���RYދ�w�B�iy���pX�M+����a�M5R*�-���� ����3���9�e�(D磉ɭ%ٓV�I����E�c����	^��%Z�j��|�U^�b�� �׋�jo��A�4	W�dϻ���f����íu��c4?;��O�4��}Wv
�<�h��=j�忣�]�M�vGѹ�o���S~\�&-~���
��K�C Q����\�-�P�p,�uW����K,@�:y?�7g�(�ʴ����W��硥	1��Y��ĳ뮰Z�����O����n�S�!+Q�=[����CD�*i�X.��!��!�G����rt���vy�i)�!	[��o���Ϝ�����.�9�o�=�`�d~8k����q��zöAk ī��@�ts6yz��ǻU�Z�$���F����XF�T�Ma���A��P� �~/t�l}es�}�2!�5�I�{-��u>��)��J!�R�#8k�3V���%��B�#k;��>J�'is�1��
�7jWk��X ��%�+�脏�]�~ڞ&���Mf��Ղ1#��em�?U�bT�4|>�:�U��!T��,�{�ԥ��y�����=�-���#@��ʺ��4��R�Ϣ�#�n�!A&��_�u�%C���ŭ.�^	�s͈_H�e,x�q�6`deyW�>xV��X���>6��7�6��n\�C��1������z��ߟ(�4̯�����2.z��A�$=�)x���ԭ��p���Ew�n�~�3I�_+�wDm��޴k&To9��jx�N�@�3�
#0��.s�D�״�B��ݶG Fx8��]��u߅zK�K�m��h�j�udf��E�
�#F�,�Հ� }Y�J%��LW4�X�N�t�T�qZFqH3������*y�X��Q變+��B-�!l�G�'&��	uŘ��e�2�.
���ļ�\o��Bl����X�tU��B��ʢ��ռ*6T�8ŗ�ԫ�O�2 6�]�rv����83m������U3��'D��ae�MPɥW��4bڸ��L8��3��2_[l|A�/��n�����m�p�Gy?�a�!@!c�;ѩ����%����ߔF��}Ϟ�ڱ-b(Z���t���$�n��UN��uD����tX��N��X�y��1��7&-7�2�\~�خW۔6K+��x���P*�(b�V��`�Kl��@���������ץ]�E����9�vf��4�z��p�$)��)�@_5}MA9H���4Z���Y�w�X~���1��k��_�ywI�q�n��&h��Tp�{D<��i�����w��0)ϯf�B�+�e��7ĺ�Z���W,<��?{��f}�cz;��62�=��$N�ts�ρ-/?�ٟ��۶wu�e�����ʞ4���O�yQq�\o覕�r{Ķ4v�ȩS��[���l16�
5���A9���jb������kd�!��6y6�(jC[Tg `A<c��G9W���sC��qW�`��m���Ri��%�w��ک�ա�XYXT�Eb�
pz�װ2VN/4��ݔH�:Q���)e�fPه�Sb|aU�P�g�h�:�����t�:%\�,�a�b/�����0oL�d��v�e��{@0"�L8`!����[k�ͪ��	�"���$�,2�"� I�Q�^$���0�r}U�����Xx3`;����mz_3�
.	h��n`,M��|/�A$�/s��r$<]�ڊ�TJ\-����7�B���xoM��փ+�hC��+�Rĕ�M*�
l���/cZ�1��1���D�A�'���n"ҷ��X�VFIG^�����X:G��t	X`�膅�Bb=���Qڼ�j|p����֮ ��1�5�տ�i�z���$��Ң��$F�T��s`t Ĳ��V��]�ɛ�1��[�n�-��bGſ���O�6�2P���'�ަ�y���Ҝ���O����i��`�Fhn���������}scث����?���!)>��@4�iБH�2[t�L;�X�uh+�]������f�CB��aev6��D�X84}?�c� 8�Xa:�4 _��`ڣ2
n�K)(��G���m�<�v&�CS䞗�:�i���^!%|w�HD<��;�LF��!��4"7�}�O4�E]U**��>�y9����ķP7�J��j��^��3���1�
\���3ް�$��D��>����_t���L���y=�.���	Ɵ&F]&����yz�Ń��.��(.*���X7�n"��v.;��|h����ʅ�˧�z��Is��u��-��,tf�T�͊���;r�����Ww�Y=M��4㾈���b�`v-w�����h!W�Z��d�MdM��yDN[9�s��Ϥ.�.L#%�؆Ǻz�a8�~�/�ek��-� ;�m���dX�Kr-�+�p��mq��@_|}�ޣ��6X��t�ֻ9j�0��jȷ������%�w��!0�r)8IB�pk��D�6���1=�9�cYW-Fo�ˇ+,\u�Dz��'h�A��"E���dX�D<w���vG�P{r����z
�����{������ղ�|���\�I1�7޽��Y�G��\����y�2��¨@�F�R�|�FU#�U�bl�XK�M4c�_N��Ke]���=�3m��d�䑙�al�MA$J���2������$�Q�S!É��sy.��Wm���쭇��q`	�ӌC�XxfCd����H���o��e�&;����P��h*���}}��{Vܕi-��6�0PsE>p0��׳}�'9x$�.��?,5*����A?��C�uhK��2+D�A�0b�C�k�x¾UѶxV$�/jl�7�R�G��/�_~��N!T�v�xxkZ����fhrM��E�*�+��ݼ����%���+��'����R<�sI���$zI��>d_U솥..[��NK�T:K/��q�	沾��$�xַ0�q���*�1���cw�z�)�E������*1�ږ������T+��!T$W^��  �kno�u�4���HЇ�SƝ�&�ݕ)iz��'�䂴���ni>Ʊ�c���YQ�=%SZ�fW�&P�}�[=do�[�EWl!����k`�>'�;��Z*�z�A�K�b�7h��4�`����*�~>�07c`�$p=�ė2�$��D�	i��|)r�׹WKpt-p�F@
&�W�f>������"3�_!���+����p��W1$�$b.
D�7�kl\�[��?�m3;����+�1�2��-�ٷՍH�L�;n�ȿ=_S�&�=R}�L��s_ ��KF�{dq�bi��[�)TA��kc6����X�욋x�@��F-��_;L����B�p����:�j���l�����뵰f��*�=u`���?��ߤ�[�%N� O�Gc��gu��YSB0�~�Ӭ�]���k�$0�#<>�[��)W��PqUP��L �#�~�X!&�j��rx4�=�s{���L����S--����S���&��~�oL����Uβ�d o�o��3����y<2;��|�(}�`!�	�_:F&��4K�q'[�p&<�)a�ܝ��ɰ���ᵴ�
����w���@�.݈���)��2�4�}���6 ��sסX�`-�*u;����cSe�u�;v���T��r9����q�@��HcH�浴���t�Y�˳��)����e1]�r_ �\�-7

�p������08�ps�d0���ꁄ��i�%�Y���p���y�i��]�9 ����Qm#�� "���u�~@E|����dT��+���sa�+���P�!����)9��:���k�yR`����������S�9�{����\�Z��뀿���C*����^��d�G	s��h�����C����@�.S*��*�y���릙=���I"��N��3��m�*���Z�c���k�C�j�����r����Cs����ެ.rSl��9Y��\��x�ّ�	 z�s������Y����Rq

F�&��k����F�e\~k�����SX;=���z5p���=3�N�䝛LA�٧���
'y��' ��<H�Q]��z->n҈vk<��1��u�'����'��������P�g��/n*�P@K��+����Jم����u�.gy�a�q��U��%��Ef�4��wx*$��e +��X^H�����V\J�	� {:x�82�6LC/����뷍s5v<���b�A��\u�Q����N�L'���x�=v��k�3.�iĞu��Ʉ����@W�����0� �F��(�͝�������*Il��4��o����e�T�m�oA&�}��Fr�q���w��1�XL.���}kytR$NP�Iš�d�|�X�ܠ�5A�l~�H%���w}Ud������9�eA��Exu(�8���j#�&h�&�I�b�I�2ꌂUR<l�;��7h�+�E��vzW�u��t�$e����vfD�w���Nm��6���o�	m�N��:C�q�G[��/kg�[��^9��7��Z�vAa.���B��3R�$��i{�e|��އ�̈e��x��/x~n��#}�,��}�kI �_|tm���.����[c`�q�>����[�r���#�3'�����n��618��p����T
�0� ڥ�aW��4�xA���uGڣ��E?���e(�a�K�uM�N݇��l(�R8$�˫tsJ�����`��צYc{��o��;��A��2�d�)}5	3�h������qz���q5Ab��4�DS!-�&�%�x8��1(�+H�CZ3�|U�Y0=|�ɚ�g�s��d��|����-6៴�6N�H�Tj��*�)��a� �ȇ��aA&`���{=c�[z�q3�K߅�\�^܊&_��/D��
:ި 1 >2��%8����p�𥀰��jmْ�'�=F�S��I?�����19�|��h�.�����l����\8�\��!8;�A�W�hI�5t�f�V�r�[�FfR]�^�	.��w���O)�gP���|�/���QW��ϣ�w� ̉ �%�y؈�:[`�_r����/�wܚ��A�Ǯ�d��'�����%3I�Q�oýШ�l�N�ɧ���D�#>���K\�����r�D�)?�c�%PEn83�ǽ	x&�l�r"dnIȟe��һ���2X���w���i�%���@9�׸H[B��b��ǩ����L^Tіp/�&2l�� ���t��U��]�����ғ��#'xka��c��	�7��Nv�!�ANXr���O�Q��.���9#�|�kۏ8�-~�xvb��־8�j��M�1�������8�M~���ܷ���ǎ �������t0ܑH�������+�i���� �H]��Y�?�9���&���C�Ȉ�ϖxZ��u�*\Iuy3�Tf/�b� ��	�~�i�6��Z�����K�/���C:ፓ�� �����03|b|@j�X�;72?'6�O~-��@c�[��+V�y\�C��Jg�9ϗ�knK�H�[/��\n&�ϓ�׺�#�WDꖺ�p$:~�|��<�4l��@��2�Bq���|dϟu�hi��5 6u|PC�I�%Y.��$��r��*BN��Bx���U�r)�Mi���`p��#U����Q�ąV��V������ʹ��Fܫ���{�H����љ`�26
���.#zz5�>���<�a�g�	-�x1�2Xf�^w�>��}NM�U�0ć�� Fd'�QN?k��i����q?�ay�sc�ŪS�];��@�e+w?]q�b:�;����c܊��[�u��Φ�����kk�s4����1��f� �O����
6���P���Z�����s\�� S��2�u��8>�X�'��t���vH��Ǜ���I�ʗ��(�?���� �%K� �,��2d�<)i^���yV�y�6�n�����w�I:�����vy\đ��v���}X7��3!�(Z�F�' 㽋�5������b��O �R�p�O�)v��H��ާ���w
4
�*���}��L�X�Q��oěbV�U��T��Z�\�DH��[=���fh���|��ԋ�c�>�8M(WOXTb]���(Gت�j�]�s/�p�0��`���Y�x�@BкEf���ru���}�'/��{bRp����;�za3�Ʃ��M��(0��ĸ�)��&��qH[v(��j�W$�`$�S�NT�˙�n�᮪���H�`5��Dn�8��N`Ğ�9���6���ֻ���د� FT�K{�'X�6<���X�	(����ء���,��D1
�9|��������M���k���&����^�\i"nE��T�����oH��OS�>H�;@ٳPq�k�!Q���Y�R�z�|��lx�S��\�����n�_�P_A�A�9�QX8�!��u�Gjw����ѮRmr��:��Z��73��zjJ��6��p �BwX�mHk�\������u���@$��e��5��9���q�T�
��n<���q����=���dC˽���-n�F:0��<�se0#l{�QK�Y�}q��,?g�Fq�9���1$��a����)�6mͫC����c��
��j��(��1����nC�H������vD�Rı}u��3aJn�����`6Ӳ=�_��a",
�)Fw�W�����Լ�'�a2�.���>�bz�]o��S�NP��l�fj�C��;�#SyRQ0���{�w����31��i��+io\TVR�R�e3�edew���0�b���r�ْJ�<���d����^&�9 ��:�9N�Uk<&_�D�G0�85u̒@���l��QN��4��+i���`N'�
�s�do���,l�W�\Ǻ�&>�`�ܺ��� ��P���@�\t�S�$Z�'�Oe�ۛ�S� o�#�s)�R���,Lt����pV���G����`���v��5I?���G4̕��\h������oP�D�"�z��5��Ǐ��N�X�D9k�}OX����'������$�Q�a�����?���=����v+�~"�Zc�����3����~m(��(f=�w�%{�1�|�q�:I�ڙ������4~:ՍU�-�C!nk�3ע5`P���+��m��1�={��eT�~`�v7(R怩��mʔ��b�x��Ķ��-��ul�i-mϮ�r� �=�Y��xAk�^�u5ﲑ������j��P&�DA�*�MZ\;R��<Z57J��tp0�pr/az��\���Oo13���-'�c_���箴Q��.K,���*�7�D�f�@͝��JΒ�J(��t��|�ze��\t�M��z�':�����.��s{�z�u��q찏[�6��KHH�L7}~.{�C���H<u��O6���T�B�����f��mXi�(�N̸q0�6Od^��
d:�f8�?w}?�;����:���s�q�t'��w��z �1&	W��_�ih�`�D�ci+Hss�nZ��w��X��1��p�A;�زDcDy����	�9Q�^����ݭO���<���Dǟ���_�ϲ;��n��
G9'I]iT����K���ټ҉��-��[h�����>��V���X�p��0*���ʺ��+�5�H2�	����PVچ��0Ё�nZ5[��|e[cXt��/���x^]�鐺���26��O��~��°D>�*{���>�A�޲/;u/�T�ĝ�2�a�a�
�s*�'�|ƴ0���]}Ld��ַ���{$����ʶ���x7s��7�XY6D�8���� ���� /4��UmZ���҇�'�p<l�Q���F#ɱ�"���$(��s��ɳ�	;C���Sx΁��B>xwm+��פ�˱��\������԰�v�ˑ�x��٠�򕴸G�j�
")7�2h�!�H�E�mR�H_rD��K4�����#,��z5��-��3&�s��n�Fuog5���#�Wy� ��2oL��b��݄�)��Db�6���ŵφD��3�{� N��obԬ��xS>=�~4u)�~������{/d�0�5G�UCq��"+>a� ��՟��%_�0o94�Q�Q�����ݗ.��=t�d��N�ͅ��?���������Qn�z"�z/���X�
�j���>��� 4��l��EH����v�nP��N�TB�$��m�˄ �D#�FG5YX��3���7�OeZ�Ȕ���������e���Ζ�a��4b
�O�w]Q��7k �Ls��n��%:��<'M��e��3_��I�H~2*��<�}c��� �4G��
�<}N�%֑7e*v���z��jp"_�U�[�o�:��(��O;�{f�!�`�t���)D+���;@��) �q��D&�����j��N�q��4*�����2�4�	j�)3�UM�Wuf��� �£4w��º8z�%z����v�}��ה������2��O�^N΁��&��;�Y+����=�=Үy���������e"T�S	���-5�=�a��|/0��h Lacb#x�3��;\l���Z��r���e)��̞�ƅ�^�]�f��Ơd�6��rw�3vB�SY���|\U�N�g�V~cȘ�4R0�qg��R���,7��Y�U��k�yZ�Q?�*i�і�5���,ƚg�T=���҄(����,/�y<�;�Q�3���vl:ٕ��{��QOd�31M��Ew�r��K.�D���閨,��8���n�D�YV�n���'3�7��K����rϾ�nmd�F����u���U�ˡ gȽܷ<>��0��-��Ǫ�3���$Md ���I�l﵁���S��1��*�B�K?Ưx ���?�����m#�!JD��+|�Z���a��^�ɍ�m
m�ME]���!'j�� R��
o��\Q�<*,A�� @ɳ`XQ����)���J&�c~�@yw#�B*~��7�b�i�f��ә��<����`@��E����I�1z�_ �>�.�r�`%wx@R�^�z,o�a�MA_μ{�#�Ϟ�����[�/x���.�ؑ������5�Q}�x�a�T8��MvO��B���k����B��q��^4��3�����{a(`�0��4�WW(�]q2,�k&����~�UL����b&X���宩� ��߄bT �����Nk��U�D��F����#�k���Q�>w�٣��`����>\�����k/X���N��v��k��Bl;�T�����cfF�G	�k�a��"c��F���g*�'����H�|��N���B�o��J:Ŵ_�`U�4��aF+��/�NS�q� �7%�.t�H�}`r �ƲW�ݭ�l|��i��t'��]�yd����ƅ��Fq9<�'�V!A�z���GʙRP6���πbe����n?�����!��H���fW�:7a�χ�:����颖��e���,����L,{���+ڜ"�py�_VM�Ê�D����t�nT**��M����4T��^����A��Zgh�5��{�:����S�2�XlD&n��SF6"��K��q$;�)cfޢÛ�>�B�R���g���q��V�Jʜ�;/Ӵ8^�E��T����f�9]hp&>/��΂m9a q�K"/����Ozc�O�_ۛ,���eZ��]y��^�sи��c���9��������s,B�J2��ݖS����-�)�h��;���+� {���'Cc&#A�W�V.��?����R��`��g5j�Td����RJzQ�l<R�,��4��~t߭@>9��'�ހ�>�<�c:-��G��7�W��o�_ �gF��l�2:�QS�P7��6g���1�cͼ�b��=�`��;3���1�J��Os~.+iP�c8��ҝ���}�̥E�.�F�W	 =j���x��#���"�H/�#�{��h���K���A�)�c�!�?)it9#�a�����eg˪!B�^��g��9.@�]:��wIs��e�L.ɭ��|!���d��t�C$��z3]U���|��
��3��*.��wB�p��)0xg��c�������_Qƙ8��Ǆ���U
 ��d���q�v��a���>� ^vq�A�r$HV�[��yo�&v����C����^f%eT����dޕ��a�����]B���r��<���S �/@��
M��F��f�j*~wu1�]Z13�1��
��:�F/w�٩����H���q�z�l/ñgE�z<�S�u#*:Y;�!)������������|b`뭙��1�+)������1�'S�}���Nd��˱K���yz�6Efe3^��""S5������*�}󏵐�b�2��\�-��ʢ-Hf�NHA�^�'�ș]���p�7�� Yn��q`/�A�S3���-Q���kB��h�ᡨ1 �=������j��f�ܓC-f��V^h�~R��z�7���H�2?�&z<��%��xi�(�
G���� ZO].r���!6��:�jpf�ݬ;��U_u�D�4\I[T��O퐔A�R jCAT��"7��ݾǖ��}QS�p�bd��
�h��QȃqE�W 6��"��j��D��P��b5W�b���e�\9�Ĝ�n�əv&���V�Z�~3��8��2J�ှ��H�ׯ����DAj5��v�/���ړ�T�V���ѯoow2����pR1iK��t�R:I 3�6�0Q����ԣg��(Z@�#B���~4�[��G1�4B�t2ca�W�+
PH�k��1����,V�oi'	P��zGv3��&�n-���O�_>{�s�k���/~n~�����h��8��w\v��2W�R<"��J�ۆ����)䢳�;+1�S��O�)������;��n@���0�S��ǟ��&Jp}�^�[?��&�
�̺�=�(?W���'3<��lq���ߍ7B*����7��.vr����tH�:��a2�p��M�j����9w��wa�����dw�6���r�>��6���g�#������x��d�L�L��T$�j�P=�
�ˌ�3!x+��ϟI�; -���?Z ��N�Fe�7��+A��Af���U�<FP� w����zJ�]a�-׍���\L���<��c���#�c���c=��5�'�4�}P`tR����s��1����i�p�����cM���������FUC�Ohq��?����#�n�O��׏a�D�}�}���L����4��6o[�sQ�G�����R'&�j=|~�����Ѳ�����jv�MÞ��}�t�	����0��p�(��ʡ���"�_���Z鞫tqZJ~y������+�@�o�A��eO
��3b�ZH�����NT�2*�H�.OA���a	�����݆0��J�F{:��J�W���x"f(����6��������'�x��v�V�N�N
ƌ���)�Zǿ����^*U��'��W��b^f��=��p0�hWl�f�;ܑ��6㲇��Së]��3��H��o
-�����<ͱ�Ō\���m)�1���$n�����I4x��e_�H;��x7f��'-�������g)��ߗv�~� �,;�p2l�G���X7շ�ƥMh�Q:����$�MٝW���3,p}zAZ��Q�R�+����e���.5��K1�8����]�5T��ٿ��R%9h�c.��/(\.,�ؾ����[��}���V+Y���_R�jƠ����
N�F�q��}�1�1 ��.�7�1_��S�w���=[��%�I����v� �$�J���,�� �u�o^����{?$�*�ȇ8����a�������]^NV��n;���Bs}�>K==�0�дs�
�/�)�.p�c#�)�c~�/^�[��>2&2D��pz�P�rN(CgN��P��׭z��(F���NR��r���U�N������u��:�M��R�������˿��>���8���`���!_Gͯ��r��f��صD�W��(���4����Fg�
a<��D��r�N�`P�7�$�N��A*3�<Bk�%��8����T��*ѦS��_���ӹ�)���1�����I㴜������K�+w�}O/���z�&D���.ZS�Fn���l��]�A`��V�6�����t{��6����Y2
��nL1���ҞD^ٯv�yڤ���b~���`�Cۆ���s�;c�%h���*Z]� d��fGY�e��Nc�������E��5��p���S�[���w��̌lǤ6F/�Bg�S���Vs����V��-5�o��N�@�c��(��6KX��;bBbؾ�H��U��}�H����8�*I���8��}���a����	���ڭepQN�܅�.����.���z��dE���-��m�<؝��������6���u�rs袖���k1b�kb�P���.����s��+�!?���&��[�[آ����@D��A8v{���L�%��H5���?AVk�d�U�;���":��
Y�6�Dy��0[��T��5��&��F��<��&����uuY�F���V� ��������%d�WT������m���}�������W����A;����\CC��n� n[n�ҹɦ�ђC5�f�د���*���t��@��'�#�Z�q���͋m�jW
��b� ����y&xg�1G��V�6G��Ǔ�[�e�&��Y�O�*
�:�!i�4t���zo�2���p>g����K��&��g3a����$pIDDDi�/Y��.M,�X�fv�ֶR�݆ܫ8!������U�����G��^BH���m��E�V�vc�H��i��F���I�u��H_�f	�@����z�)i�p�e��͔h_��0���3�ط���&LqhE�`�b�`�9��j��Jw}����K��,�|���E��'�}�	`kd�G:bÍI�m�+-Ey�y2�LB�Ʉ����s�x|��������|��1�g��s		ˬ H���Ni+;g�����8Q����@�~彉A|v��p�{O�[�Ģm���s��&ٚ�|h�#����W+���l��w͛��O+�Nz��(�������⺣-u�D>��j\s<�����"�.��QМ���	�m�YQw�*F8�>�\\��g��L��]��|���Ϛ����+��an~E�%�^*�9,_~CЅ�d?lV!�	�N
���+	t���gm��ֻM�ˈ��Z��z�ա���ķ����؎��� �;=���~z,�B�p��Q����W��V�r���#�2ڔ��[F��k��f�˦$��gKG&���h|�����lC���V���V��]:S��f�R����m�}��l[vu�b���ۇO�U����-���N�ík��3��}�	�qPX�(�j���B�ó��b.�_�eڑ��!iq璦ח�H��+���C`4]FVM�F���T/
Ӥ���6�Jo�A*N{8���s�G.����	>s
3i��%�G���U��"b-�:�Λo��t�� ��F��i9������-��HJ�H�N��ң��8�;�e�+��X	�od����uwi���ߕ��w���8��A�;��=�ou�l���	w$���90����Jj�7>d�`FRSpm��^}�"I�������z?I)op趿���0���Xp��Bw7�o��{/ �4��ݩtIH���,�t�ҝ��"���,ݵtw��{���s������|���G
�*I��*F0��H@6��R�"�>거��6����A!o=-��w)k#���p*XL{�V��L{u;he<���*�X��Dzːg��v�d$孻��3�䒉��+�y�6����
	al�E�i�u�a;t\�>����#�4��Z��.�Ky��EE��S�e���3)}�&��v��]������S�z���08�#9#+�Ċ�Jw�0w?�-Z+���"�-\���������v�� l
�~+s�t$��6�ӥz�~����ǑiM~�+�����`c��'�H������!;����O�����^�k���O����2�i������7�e����[��Z}`��ê��tW��i���z����Q��3����,G[�Od�i�|��#ߞ1�K,[�5ε��_l&��)ɗ�<f=�v�V��!�ױ�q��9t����M�p�/]]ft7Y��rg�E�_}k�������Gj�����sc�6c;��-L��ޕ���h��H�]߅�|��ZM폣Iѯ�?]�Exd�J���/	�~6vNu�ѕ���6�������G!�2�}C+� 4�xq���BA����6/??X���eX���z  :�/.��}��@}���������5�x��,R^}} �/� �poZ���t~��8�2AG���U����9�jB�)��I_x��~;|6��S^�<�z���*"WHi~N���IJ��된�N����6�/]y�A�Y��Pszg���Q��>�ӱ���P*���.��?��~�*a_8�}����5�ٟw _i�_�
Y&Ǘ�>�o�wQ�+�FK�L����PO���3Sh�B��Q�U�������[��n6�Q�v����.�JP��N��N~ԫ�юN��&��6$7�����[\Ux��:�x�)n�cT�5b"?:�$�Zf2x���H�"�����������z-�#ĉD�������q��w��_x4��~U�}͖��N���2��=>�=��4^@Q��S��yM8O�hs�ba���5P7�ݭ�kf�{��$�	lZ��/`ܘ�N���3��q�ߝ����;/�)��L�2U�0��^>�6���
=����,��N�h�vT�R�ܦ��	�k.�<�e����W��$����8��]%����������#�g%�ё��g��K`li������ȣ�"`�ߛN;y'O���5m{�b��3?0C�]m۷1�A{������#�+�s,�Y5�����|�����o���uQLiT�BėW��!bc�#.�I����h�)�j��uq��u��;�����j���?���F�l�c'l����Y���s��לjk�
>ӝ{���C��Ao�N}��K.�.�FqC�����=�2�6���ӘXY��������`��?tr�d2�m��׏���DM&� �%Ռ�؄�4?)��,Re�۾�J�S���j���},�.����.��܌W�]}4iR~]�#
�b�O�/x�W����+��f o�b��������jg��l���:��c;~D���mt��C��6c��Z҄ԒS��2�������s��|s����J�xC����z��S�+�,5A��px�w#JY�}�}�mlx_���%�U �� ��.c���OR0��0��
�y�-���������!~3������[rm"�z�8�����nIJj��i��輻�ѡ_�� �o���)�U9 �]�:0��X��B��1Z�V�*��6J�q�6���O�[䱵�@Q8��N�d`r��'`���
�[�<�@ė7��]*��ȥ������)� � Yi������C����f2(Y�>Gp>������AV��9Oز��%���?K�����/׷t�1@��a����w��� ��V�+��߉w�U�'L�&�@X���:��&%N�)Kͬ)��~>��zi�����|�>���G����c9 �����E�����ɾu�[-9���x��:��<W!���+PZ\��h�n��ҟ��嘎�~���k��O����}^n��F9����/�bU��E�9]F|�tTx?����9F@��������T�cz���0���C������?/6�������[	�"r�.*��􈈗��H�ጱ�}�zM�h>^��;���KOG���_�ٗ�-*<�j��6!גJT���^�bZ����-+���LdG-��wg.���'��!��=���a�?yr��4�6h�B�Ek_�-�	�������f�rD�����7���)�h�Bf����p�&��EnN�?,�xj��B��y�����BO����$�b�%���ה{��9�Q����*�y���b��\&��f�������qyV��t�k��<mɖ���o��*iJl�:!u۲x:��N���z%7�/�ۜwU��� �?��R"�u�%}��{
���M�u�m�k�G����pA���lV*�/ g���fK���y���b�h}�����	�/��,����c4GX��r�&%`�~&a����Zcg�:0L?��@7c��w (���BZo�&�i�0��[�/$0�J�Hby���&�( ���躻q9��=�l��޷���2lʐ!ϖG�Ǉ/n�$1bYo�W�� ^HL�) ���˼EbBO�'&A]M�m�?��Ås���o��K��Fgz����,��HB�K���;� ���Q9e��>9��>����Sn����)~oL@���u���`
�nn���=Ƨl�Y$�NFP�I���R,/h�c\�[U{^��J�F�`���K�^'c7]d�+E8�0��P �}��|`����`�sV�s��&�������rw͆�4�u�D<��S���4?=�0�o�Y�����X��^^Q������s _QBYlD7lL�t=��>�:�J���x��{����'�����d[�i�o��891$\R%��!3�N.�ӷwk��(�=!Ȱm��RyW���&����ewk����}�\����\�Rw�!���%g�7���G��MC��}$m�]�b��J�z��tJ�e������l��/t)��JJ��1o�R
ˁ��NrD�(	��~R��rO�7��00�hrĮN*f���Ҡgq���7��N��"�ч�锦���7|�j��3�7�=K�_�?�vR�2��$;�B/F�������^������Qk������Z��r�=TC=آ�U-��&�z��5~~P'��	Y�Mv��}`׌Y�h�`��+wv<�Հu� ��8޷���wLL ��i���|x�J���yL��4t�#T��/�@�:���D_�LX�v� �x�h����dپΚC�^N��BZ�m�Ŏ����"��w�	`��F�s�O�w�d�i��/3��b���D6��X^>�Ar~4d�K��|]�0��ŵ
���\�ar��?8���{Y�1H��1s|��݁��l��s*����h���D0/�����#���y����e*D�C);���HG�s̕H�-J��h�&��E��:���G�6.���*t�����8������;��9����A�u���!�R�T�Q/���e2��GE���p�y�/� 6�BaE���(΅#q��h��(���Cqn��I�\{��`��jf�8�^�x:�]0
 {&F�{��o"��x�m(H�Z8����ڹ���Vҏ��s��>Ҡ��~�y�J?��h��K�r�ؙ͏��=}�2
E��y����В=f�UF�Fq�֗��r���4��z�C8���EH��V���}*0m�j���C��n���J%Y�jB��4���-؀X ����C���BN�Z��U�GRM�*� ����/��U�wI�eɔT7��M݃�AF(��{xzc�C@dc�����B�z'"�����6����w�ŝS"���yT�ȏKfʹ�	M�����Y_����h>5��U�JҔ��aT_�@��p�j���F^��8#�$�˩_�=���|���8��<)��N�������S�a-���Z��E��� ��������*�����b����&
�t�Q>ʇpb+�Ȗ����v�=�u9[�h�U��eTfK��-M��]��$�}�f!Mk�kT����򢡉~�����6|E��P[�}{l���3�2F6�멙�F"�(����ϛ�($yC�`G��tYo&�F'��qUR��f7��:b��m��l�Xiv��{�}�e�� O[�HE�o�[�]����V��#ԑo):F�yךگ|��p1�(1�[! �������rGs�o(���,�j����ɼi΀5��D����D6 ���{��N<%�o6�.6{��C';#�Qڍ[��KHɭa�$�c���F�{�Q\�j��xw�y¶�����6����XW)[��ݖ���H��aq1g�D9��������,��Q��c��֡���'��N�|k9��Ꜵ����y��̇!�h��_To.b�����u22�%�6��s��%؆)��=�'}3���_.�����H���ne�N��8o��aM�݆J�.�� �u.uC�P�Y�b�n����!Z(o�]���߾��;�)�B��&y�i���z���m�l`�Q�������ѭ��7Q1WV��+���@�h���h�ERm��!��m?۞b�#�hI�jJ�%�ݵ�ћV{zۥ/8�}=����p-��u�u�h���~����Te����a�ͤ�l�U�gi��6�\��2���'����bt5��X6/kn��2[i����o-�d5���ۉ����L�O`N��k۟g���Bs�3���;cz��<2W�L��:�����M��w�D+��w.��t������
��\~~��\�;� ��s]8�_�O��h���
`Y��F���|e[��0ԏ֢��Y�7�#�L/�C<=Ŵ�I�IC�Ά=�Es�rc�d���{���H�䯢�\���;�H�Η�MU˩n7�cY��F[�����-�~I�o]�7k�(ف;����H񆄜?ճ��IA\�0�i��0��~�T-y�Q����^m�7s6=<ZG[�=q��U?G��1W5�ϴK��F� X�m. �n�9>�T�^s�V1+��>{.7KE^Bx����d�P��I2�#?5x���ݩ�A�<�}^�:̚(T?��^�;~�1�Ѩ
��|�w]�);�)̒�&̆�҂d���SI?���,���k�Ac'"�d�c�z���)G~��cA @:;�Tw�ׄ]N`��ޔO�7y�s�K����[U� �¼ҦY�)!�)��=�4�LN��z��%y}� ߉5��v�Af������S��}�\�I6�9/�8�3�����V��r��� c�����\S �ߘ�D�&����E��	�~�[L��q��d	�{	��'<-�A�dK*'J�y	o��E�J?f��a/ڻjwϛ��D���Q�K��q�{�&=��s�u��w��Y��/֫�����pV ��5-�λ��7{ί�.��rPr���L_;"�1;��.���)oE�Q���+s�K��w��{/�n���O���`��L�u��\>���W���d��"}f�A~n"%bܛ�ij�*+�;Z��pR>5�n����3����QQ3!S���B�]��֦X�������R��Z�%��k��<K������w�<TP��{��i,��>\�:�$�µ�s�����%\�H����E+U�M#H�z��[;�8�r�= ���ʩ��Al�9:8[���6�r���(~K{T��
B�/Ͻ:+,˝9�U�����@��i�L�ި����o*/���wP�𻫻��dr��]�Fy�D�<RMX���q�෸R��p�����l�oɫЗљ�9�҅�.��+DB���@T�x��Ϧ�,q0��H�7����
d�d@���s�������� �!���c����N�%�7�p�f��_�Lֿ����~$��?3./M���qr�:=��Z�6�8��x��8!ݭ=���:�n�?�z��g�(Y
���BE;~��6u�d��tQ ��{`m֥y�L�o�Q%��}6���gjTK�~�@4�¬��gOK����/G�C|ei�%��W��wa(��R4����20�+b��}1�N+�gL'��d����v���:� �0��g����U^���:��%�]䳩fx?�up�.�����&;K�#�:es�Yr���ޡF��<�+�ꮪ*c�.���H�mtC�N#5��=]8��ɿ����Z������������/[�+F>�U����5~W"����{����W��2��\��*~,~}������,{�||�_�1�L��A��U,��U���fXP)��V@t�E��8�b����(��%��e!�U��q�b"2���â��E�=��W5]��򾏟�i|K�j}��o^��<T���oJ�9�%9G�7�,O W}HAu�!���dy�k���*���7���2�S���CJ�"�|z�_0#�����?I%�]�8N�Ƥ�8�'�n�]��f�g	��!Xm�ү=�ixOnNa�*��ۋd�Қb�"ƭ�3~aK'��o�Il!��=��ﮎ�G7?�8 ]�}r�	 ��U�vx�_�$͞D�[����q�#���}y�=%��Q���<�$�ω�~.����@�Ȼ�ρ� �����Vm����)�R��$�~� �Om�m,v64&��#����߁�)c�~��ivaKr`��^*Is��~��#H��>�(�8a�u��瑼���a�b�r)�\#��L��.1���y�+��#۷�ו��!8��ǧ���\�ן#;�c�G'��^� 0\w��pQ�2d�S��G����m\���eʥ"'������>!�PcV���n��DB�҄Q�^��"�9i��]H��/|z��+2��4^0�`֮[w F�"�r�$؅?8E)�o>��A�����M W��0ť"�9 T�0c������Y�m���:+�B�߭[Z>�[�}�4���Ȑ?#�M��^qە��n���3����O�G���v���o�8�:���nz��2���"�t���G�Ɯ7]�ݍ<q�X�&�6/_���Y�7��Ѥ��/�Q�N��J�ɵ�J������^���|��.�mvid���&9a��D���*��s��~	F;/#�H�3�u&Xv{-�S߳-|�����E+t��)Ӵ6���/o3M 2=�k�OZ̧)��9�Þy�A��)�fu����N�R�.��{�"��Cg�[F�-��?�]|��m��~IULa�(cK��Xf��<�&y�N������l��8h�;�ť\;Ւ	�f)`�#n�/6'gВ����L�Nr�P����[1��cJ��_��'�W\�0��u9�Y��Pi16�'$��T�t�{H���g*�;!�CR��
Y�@�t��t,�Q���%5z�;�:��\CG�����S�+�z7}��cll��y�pp)����,&���x�S���h���h+�b%��T���T��S�.Q�8�����χ/��	��=V���8^A��]c��������E��X��T���FV���{C۷�j�������Vt��+��w��ȧh��v�+���~?O�h%���lZ����st(��23Ĩ�[)��]-��pX�*�	|��3x���(w�E�Un��\)���|C�~������.͵7$�B#V�섺�����\&���a��/Fg��i
�Z�j�-]Ax�G�\a�/����ч�.|��H".����ɹ�����7�`3���a�fZ��Lcc�S��S�}!�W�b���Mş�2�2J	�jp�2s��?�@EW�%T[��sۉc���Ҽ���=Rb~����z�K���_tW���A$~��
M������K���N"��pOy���՟p�M�p�n탊w���5oz��|����m���m�����7I�|�V�/r��6��	�BN�V�7U����B����㑆=r$&��ؙ�#�=����:�e��Q"�(r��y�h�&���\�W5�_k-cο�u W��
=����%�B�L��ȶ�sAEJ�s�XGPM�]�������x'9ZǠs9����O�I�?(޵FX�Aår���G������JF�
E���J����PW����H`�q��K����ڔ�O�ˏN��UR7տ��5�m�ժil/���.�/#`�}؋r ��h��g>�ў�O��;gLs�ZM�^�m8��f$wEN�j��@!ئ���?���NԂ��I��t⽺�j��C;�.ޣ��W"�UY%�(����#u��4���ˡ;I�
�#ſ��Zs�:w�'�a`?��hk�[^[���L���B�2zeю�h�>	p����i�ḱ'�%�����3.���{��s|x��x�^�6��j�3 �M9
���y8RM�{i�m�I/��̌�l�Y���s�إ$��������ZU�dʤϦ�KV5�}$T�Bm�ʎ����|��vD�2Q�L�������|,��"{��R��2Y)�ލtD����(�p��,B��� �BN�
�j2�Ӫ=qr""LUO-����~�%���h�7j�08>��ey�)�w.1W~��(U*�,qʮ"+�Q�!��@"� t �����,i�����3�:U��Pxo�(�ՈEG�.��w�OhN��Z��Gk\K#��it5KiB"���6�ro���S����X:;*ZM(�o	��Op�-�����1}݁�E�YP;��������z1��8|�����1[�#:�(����?�l3���],�9{����3�-�0�$���E����/�y��]��:�����_� �S�y�<� �
��Y�	����tm��a&���]�*�����sxEkw�F2�{q�K`Ztv~Q\C�E͡���)h����N����s�<e�Q�����'�W����MNe����'`X�i�t|Q���B'̤Y�4 �g���K��j޷���vW;J���=�デ@�ɴ CJ�'m-��m��@ �����P��Q�β<�`CB��0E��r�}��'C��-�n�v�� ��&P�"e닋�b�o�f[d��]>l�g٣1��P�6�̺x3}jZ>��&D�dG��L4_ ������e\42k�����ל$���b�6_�TO��Z!�Eg�E'�\����;c.��}�?{�Ia���{­*�l]RťJ�U��]0+�O�����r�Z5�JB�M��lp!v��	�:��"z�\���8؀_���f�-�sʋajh�W5+�i8��l�JkC�+���W��w��:��;'�pB!aj�t/��Iۙ�6�|K��Vq(���N>i�ǹIy��`x�Ka?k���A㪮wc3��[Lv�1{��G��z���P����I�"[��>�u�%��o䢳�"�߂�q��Y˨����C�B$a��Uי�Y� �
���Dya�=*)<q���[#��r�ױ��lT}�,���IY�K���������|�?r9�Z�Z$X-V|�<�R��ā8N�$���j1�腡�S�D;����D_���!4�O��/�d��4z�.�מ�j�[*�.�vG��5 �/!ǁ�����EG!�
�_/���� IwG��舁��&X�ѥ{����&Y�0%<�=�-I=>M�QǗ_b�+�|ql��&��r�%��̜<+Pz�'�m�9�}C*a��\�/݄D<�V%���f�V�⠚��gj~�}��s��{�.�zD����ITy��V���}��%����ISk�bbB�����|����i��t:&��h?�j�JUI�RL�Iy5��UD�a��T�Fd�y���d�{'��#	S@�-�۴��U(�xL�_�2�m�2��"C;�U�Y��z�掗�_}s��-���.NN�|V@s��U����wU����V��<[F�y��y�w�iB�+��?���=�󜤳dv�bB�6U\Rw=f��t�(]����ף�\����:��kt���T��UM5;~�{�$L�}�ײ*e�`CW��N��W�ޱne�y���|_3n��E�E2+pa��!;��W��bSj}gN��w���Z\�
�%��X�h� �|�'�K��z��ِ�*#����X���0.S"�@F��-���T�c��4�y_���=��}l�9�2�큿�"S.m�@����Y�;U|�J�e�)E��O�Z4�}bn���l�P1�[��j�Cak��(5 �+�\�j5��!�ط����C��n�h���~�aW�Z(����w?�l�}� )Z%&(�M��|w�u�NM��)b���-�r�Mw��Xo:n�0���@&3ճd��P|�ݭ���m&.�[-imI1k�ps��dC�����9�0�8�S[٩-_W���q��ѻ�M$[���ɜ�1E@擊�'���k�׺>6���[���ײ]5��m�����"Tt���ˇ-��@�;��B;b:J����>��η�]����6�{P,����ȍs��f�1\����d��E���6��m�,�7�*�|���(b?�,�n���#�s1c��S]���?��#�e��G�!�S���ƻ��!Aے@$�Oc̽ے��q�ﶟ�Y�a� k1�}��D������<�������D��8׿�	�~�s~����i��� &�T2AKI�n"��t��cY���wn2��T?�LGO�]�ODK��*Ɲ%_�[��Q�=�o캐��6scM�&���l��\�狑O�E[WM�a�+��?��� jUm@�.�ݶ)h�휺:��6e�L�L�/J��[^�B�S���`v���9_����
������q����rAܲ���Q�>�){�ҕױ�38�%���'W�;g����'���O��Lb(0>�s�@9 )*f�a�Uw�'�w{`}x���l������*�|v��H_hmw�h@vs�n�*^Z��*y��j��|��)���4ͭ�����N9�����",p�[*��J���a��*-�����AV���M/A����N�V1x0?�1j�]8c��dS���4G���CҖ�����MD��qx��>�s3��]>��P����̝6��r&�k���Ua��*$�-��{>�������Ed��}���INX8O��I��0��ĵE��TB�)GQ��5�Y��#B���C�$��E�����4�W�qCw��]V�-»�ѡߔ�{]��]<�ĵ���\�G�kz����{*��B o��:_���I�B��U#���3;&˝a��2��.Z���Uܹt,�-�PAϡn�.��靽���B�w��\���-_f|��<u��ꩯ��t��
�|������n[�i5���a֥��VS�C��n˨�W��2v��ɜ^�d����'���yI���/��$� �rp'57�����.��ufE�:;74����oŮF��\TOD}H^U�/�
�&#�)�yq[�Sr�!���h�~��yeëH)uT;%3]f؈�3#'^�Z�K���L;c�l+-�ζ�y��K�r��>H��A��������ҡ�I8m��D����#�Q��s�����O�tSz�xH��ܜ��$���W)Y[�_�U��������ꉬ:��a'�S!]��5�S�����<Q)CM��BK��6uÈ��Ů��U��Ȭ�vU��f@,ǔ�u��~s`����!�tz�bq5y,ۡee��jhE�nS=��'a�״�˧%ٸ��Z�������Oۣߧ5�%&_	%ǜ��N��YUp��K����⮵�r�~؂�r��rS�n{�t.�W�aa�����H����3�ͻ�]�i>�'����>�w�&�z�ԗq���]�?��6��*�fQ�4[�kg���6�C�4EB����+W�O@T��\�^;�ȭ6
�Y��1��S�ŖC�<���}�b��-�#h�s��e���Z����c�V�����CyN1R�Lt��W�I��Y��L#��xfa>����}Z8�s��1�fg#�hdȀ�p��rP������,	n%U<Ȭ���\�c�B4��H���c��c �k���+�Nt��n�Z�L�h������v�o�K��eNQ�E�Y�XΛ��܂*�2+6��YL����C �J#�f�|˨A�A����כ�6}4�k7B;먨�5�RѴ���:#�ǈS[uz�t�.WJ���fĘ[�H<B����qU'�L�������@8����?ݏ�#�R?�(��1��tx��wQ\c�d�y�22>��� ��JYGr5�fo�}�J ���\�����G�-�ֻ��M;�jʾB	���ɱ� _�3#2���m��\�ࠄK���'�l�[28�懋ѡ"�a�����$i�TOe)�5"���y{����E�qRL�(8�0 �*�1+6b��f��}��+�V/v����euU�tDm�z�L1���~��5խ����$>���i��H�ة����NL�Q��m�iLt˯|`�w�b�~�]���3�� �XO�kKB[��7��%�u_t�)���Sk�9a2����v-��up��t�w{��_��6Stt2�����J퍅���U=��ސ�ݦ�/8%`J����?��9�H�`�-
N>F��bw����X�0���$�0�B�LYM���F���1n��en�{��qy9�{�=�T9ڕk�n��ቐ���d�D��=�˵��g�_���.I��n÷-��jIL���/t;k�2��b����������cjv�V�y�E.�9�,��+[~�����-V�u��{�B�o�q��x��O�8��3��6e��ۗ{WwHE��
��EP����Z�ϹY�e�>���@��u���.8/�����:c�>T�Q �|F_x��B��B_5��_�nZ�ܗ1^{�7R���+�mi���ɻIS�����˅���ǛW@���*L�F�u��.�n(�O����4��Q���.#YH�^�&�q��Ǧ��*J�$�4ɗ�d]�����N�b����:��.T�I�m9l�jj[K�N]���s�@�������ٝ�+0:�&#[�-u)�V"��u�\89f;h�������0�����A���݇��
����`�F,%��x;��¿��@�|y�	�(��V��z�8���.29L%Z_��N�zKZ�1,��.-����$Y�9�g�c�g�	�dP�����z�?ad +9�@-�V1<\�D{��q��$y��P���g�L��*���^r��R��,� �a��L�[\(=���C�Ӗm໪�M�����W�S	6Q�e��
�Mu�ǻ�����J��{qc!%�*�����%u�,��]a�
]!mĊ�z[��^��(QZO�S?,�g�v�H��H��h���8&:���BG���pú��h��8;�-�S�,̃�Fepn/�\hk�IFs�Z�$���$*�6�a!3�6��)p�Md�����:K[O,W�����@��'�p�k��ښ��g8ω)q�!p�U<{O$b?����݌d���aȘ߆p)]����%m�"���l��8e@gjB�㈭�-N��`����g!�C�u7R`90+�e㔰K�����Y�g��]+U�<os�g8���I�/ϣЙ��r|k7�p�+��Y2%#{�x� �����2&2���	��4y��6�%J8\#��bM��k�u��H�������/�}@Oߊ�O��\�X7�֨ ���d�����;�ٕ�1�.�H�?���,�@f��:І*�d�5���N250ӧ-�-{,��O��
�?�
��Qy[�M�%��$T�j�0N����n�q�G/�}*���x��T�������0މ1zU�������{'�>&qԲ%3��J��0 ��n����+�NN�=?ƨM����J�����v�a;9E^��h$r��{Rs��i��r�&�F;��>ۿ翧3�iF�C?��v� h��,�$V�_������Cw[�����������>����B�1�.��i�	i�'&fְi�Cjޥ���[i)$����������"c��K|y�\>���7"���-��(�`�o�T�<2"�#fe�e/a�܀_��V��	h��H��U-�3�B?j�t҅����Lz,y�/��9T���[�,��1�4���]|�|�-�Y�P�?����`��s�T	����w��+a=0��+���{�Ǚev jO7���/h�F���xfdI������W5� �P���� )����q˻6�sL?�Z����N�>@����UB��gH��C���<G��&����:w.h�ک�3�ĥ��$����H����c�o��c��[�p�_�x"�U�:�Ʌ���}F�XQ��j\+����4~��"UpC�| �GVd��8�эg�rږOK+�{�i�"�ݟ�;�J���"���Q7�q������E� �}Ih�{���{����JF�����LaY���4�ȉJ<�:�ǲ�il���z �O���P�以�3 %�Âk��`��G�����P��Ē���d:�b,A|��D5�&�9�*�/�[��A��a�hU��L���!Vb����n�Ȧ	��o�Pd`$�c�|9���d���9XK�� �S�s:�%G��f�z��-�0�p�mK�k��c��I��aߡ�?�xS:<�k���Q��EM4�w%�`���s�����/o��!(����q�A��@Ut������n]�h�e��T����
��M���qtV��#@��-��q�q���?�:g�8x�7+GvW}��Fi�%]%t�i�$�3YrG�kK���i ;�%�,t�\���7�E��YhݫD��3�d�"����J�ðل�{@
m�F5$fhΝǲ%�6��}�ͼ���<L��*���ݧ�?��	�+;Z!u*��k=�9"����^9�U�j��MӺo�i�	��Q�ֱ#�=�t8ܥjec+?i�e�i�:_�,�,��)�&�ʆ6^]�FǢ����fy1**�ъ�RD��c�M��Q~��F���jv�( ��}q�F�o�Y4�גD�znO�3s��K���]x���|��z�:&���K���2���r��qO�_�Ձ9�)�_@�LZ��vwƸ�a�w��`��5H�0��;h#��N�J8�v˵;^wy8�)f�!��B�hĤ:t�i�C�5��P$�5��=���\\���I��r������C=�3B1��ן�{�<|�P����C��*��]k�|������y���ԣm_#*ĩ�z!���q����S�!�5�K��#2cx�F���q��m��7{�E���l�徸[�d��4�[��絤�ĝ�n�YF��fic��n�Ԯ�~�a�ۻ"F\��� ��Ò̭^�Uȡ�d��Ղp�e�����p~�m�w��$�(��NYZq��-����~�����4,�e�;#�D�i� �̞��7EJ���F��.j��J�()���J����g,<?D�{燰(�?*j�T?����j��{��1��B�5̘�R<p�G�P�T�������9�<s(��p�hw] ���>��ip<*��gU��x�d���$j�!�I��F�b�
X6ZiKnY��,���a�Z�װZE#�O�vV��Q��qM"I!��N ��u^�*����ʫ�n���/��Ń_V]�K�0��`�n��_Ѥ]�鸖TT�;4��yo���T�����*��/�F���_y:Z,�V�*]M�וqوb��e��!��+szO�t��h6�O��X^1Jm�!����T�����g��j�u~����<)w�!�Zi�&�����!
���`����-�p�g�$h�G�K�I��U�&ovx�w#Pл�H;�)R��D����:CIN[2j4��-j��#��B2ZL��5sF�?r�-D<�&��kZ���M�+��@��j�2��a-��%���~�@��P�*'s�	x��x~��ۢ]���OU� �I������o��k�g�!�V��HtGT#��<�|l8�HE�7���x� :�¢�Q������q�{a�Fqr�;CD�l�1�Z���~����p�ν�I��Ik�P��Y�C�կ n��֪�@�êv b9�l_����
I�߰�@M]ޏ���,<�:�B4�Ӵ�|��h:�_��fgC��BS(S���5���Q����ciݯEǺ/��9A�>4R�D�{�{�b;i�6MVԸ�m�v�IccŶms���ƶu���y���}��o�9���J�A�����J
��Ȯ�C�����3w	~(jE��3x�uY�ߌE#G�*~ȴ��=�%C���	sP
�x�_Mcz�?�4G����U�]qpK���kl�\��r�`��ps�A����ꐈ��(y� %}Qo�ڻ&o���>O��S��B2d�g5��6J�ŭ"����ǮI�� �mEX�0����`�aG��Â@A<H�8�g�>�����b�Bc�l.b�ϧ��<σ��� �`����<&���ϛ20�Q�'"�&�����*�щ�y�f�L��fG��	m&�A���  {���H�>6.s$և�����V�=�+ �≎�� *UQ>K��q�OwEH?'�<�� �al�n3�^��1]��� ��Q4�l���Q6�A�'�T;��81���F}mȕM׾F8vպ�j�8�%�|�<N*p�5��Sg�5䭒�l�������	�(�����eI쒿�lq��Nv��������:"�=��}*G����u�� S~��%�@��Ϫ��w��N�j�6$��,�&Z�R@n���Rg�O�g��ioL��[S�[�rz1)�QW�{�ߨA���?�����1�Kqof�������.�Vs'��q��>���-�F%B�F*2}i����U��V�����z��.����18���c�|���#�_�c�sJ�l@C`�8R�����=�-�o��<ֵ�⏋�SDJ�پ�u��M3~盨��T��'�h��iO�u7�v���"��zh�j��-ן#�뾽�X�c���dxS�%��=lit4���:\�cլt�%��,I�Q�ؠ�e�E˕��4�X��]��9=;B[�v2�U.�nڳ�{5C��+G�ɴ+�\�A�CJ�V�P�p��f)�ʚ��eA�(�ʱ�NP��|*;��&�θ��ֳ�(�,w�K ����!�)^�óN姙���p� �k��K��9Ш�}ĉ��̃ߧ�x���pX:a_��|s�yu��j�!̀@C���Uv&X�G�6���@��QT��s��J%�2�΋e1����s�f¥[��QX���(/&��e�S�G�t-��7�q<���z� �UH$�<W�U�z/7�@I�Wu���,����i��o����d�(��*- u>�!e:�IH�r�x����U��.���ud�=.e��ڈY�_�Ų�1.�1�l�B�h4���M�-:I�����V�l�S����h�Y��%�'�E+T%*/���؀	W~;9�������WK򋧩�>rxG�_�鶰��h�l�{	�uN#�S��qV%@~����u�G\���ʃ����6��Z]��_��4�M5)m�v[eٵ�r�iTo����!������ú������<�&�7��#�l�ý�����������r1s�r@@�����<ºW]�)V�џ>y�V��b�a�[b-�=�~ʜ�V�H֠\R�L�����a�UѮR���8
��{@�.��ׁ�ҝ��J���	u:=M��w�e�7��Q���w���qe�r���U�L;պZ(%����ŜI��oq��(��f�mؖt��S�*��p�-R}d��{�x�6V�>��ry�6��CÅF�t��e���4a�1\:n �sS�yx��C��I�eHR�Ip�U�m����g�h�1�d7w?���9C�����G�Zt9kB�IX$�VW6���xH:�i�x��{��d�7�� }O&<ȳ�KGޣ'�8�߃���NƢ}�-}��|��ٶ%��g�`�}���9�M]�`\�*��x�%V��/*��ɪ��;�U�
$=a��Y��b����?��ڄ����E�on�F	G	�&�MN6�� d��O��d$�|��Ν2����P�LR���E��}�U�g��XVA*�'2A[�F˦����K���L��1d:���ԯ�;~C��_�`�ErS�]�	o�~߂Ւo�w��U�	����h��^������rΦ3)vS��n�ѝa��S�lշ�DI��F�^k����=���xn����%���no,gR��=�eSK��r���I"� L�UE��X�#����ä꽭�̐��d۝D��Ν J�JGe�DE�ccLBQ�VŪ��5��?T���%#l�o�Jk�g�c�~����6
n� �.��o��⤺�@�{��H�Y-)�Y�-5[�>^�����tުt�ԕjT*y�g9�� ���J \��P�ٺ6�$��Nm��Vʅ��m�R5�)a4��U��䧔G�y] l/���n]&�e-�dNߜ�Df�i�?h(b�)nH��rCф�{B*��i�0'![��dl����s*�*�wW��nF�{���޶B�YX�����C� �k�j+ׁ8c�F���jf��]�p�zVP�[��Զ���#bu�M��LS9��Ԩ���˳�K����������8�<��0�Zx~�1��]�_��� z�U������Qc��Њ]�� ��xSg�T!8��*l�ڜ��� U|,���˾F�E��(Wꍁ��g����-�4S(��Gـ��Q���)�[鈳,�I�9�W0�.�X�6��"�Ǧt�O]����Q���<����Ҩ|���%kU.�J�G��(P�"wcW�%����d7S���p_�挭��\,ּBN�����ؘO�|���2�Ҍ�Pk�>�,'�)�Gsh��FX�d�n~�Ys�@�J}˸2Al�9.���O���|�t��Fm(�Ss��3�' ��|��5eV���&�˻L���``,��|�������ln��dJ_��E;L��ɟm3� �	p�k��+Ao��2N�u��&0p�M�� %��Bv��>E�8Q�XD��Q&�T�e�F�(Ǟه��p�r_��j�4�,qSw�WY�˳�)���YO_�'�_��%���{Yt�c�r��Û��Y���wf�d�UM�/�p@=����`k���di�B>4���є,������;;h�>��.�_鹳]wv�K�F㻎�`�^+�.D�� oX�]Oq�*xt�m�9�R�3i�G��6ێ�ȿvm=�u_�>~������9͊��>䬥9�_�䵴Ȱt/�av�+���B_�����:�R����:ld�W5=R}��r�FG4:a��K� ��D���j�ƿ�6'��8voD�YkTP{8����qa�h���5?���޿ġ���5���Xj���0{��/P2� �W�ë�e
�E���rXfW��<;j;�}$j��SZ���|İ¦.��LHz�����'�f�Q�A�^��<w~�̷�7veoT����F��+�(%G�J�JVC����$T۪{�D�V�Bߦ׉��d���� Y]���x+R&��b�躧.�R��xf��qWHT�T����&��c��k�9���ZtQH8���/i[M�!6p1�͡$��b�^(������t!��jH1H̶�1>�s����'��V�Z�+�r��5!�?��ϒ޸]��)�I��A�5�1)#�,�W��+����+%Ʒ�˱���_�#]j����G2�dӽ����S�ׯ�=�$���T ��w�g�E8�8I�2ʒYqh���R������aF�y2j�.�.F����	@����~��ж	�-����~�duO���s�%p��Zh�5;L3t<]��%ۿB})%�����d.��Ѵr��:�	MT�0 �+�B*K�%WS>��U(b�p �_EsC���(O�Z�k��~¥��?�y`#1���S����j�mTY/�cY�&?/�Vr���;����͟���ʄ����W;i�+@5vD����;uƛnKg��ͼ�k����
�i޿4a�A��߼�{�5&����I\���˾�&��1H:��W����_�Oc���FKS\��r������XX@ٰ���Ss���*Q�?�G)�	FZ�v�I��~fq1(�S�*$��x�4t�K�7�_e�^��+�YgX>'y(��"[�7#�)%G����pjh�͉��*�d^�w�e%F�-6��n�U����&�8Mu}\޸nK��a/����+���a� ���C������O�s/A=�\b�6/k�/��[sl!>�
;���ϐb�XS%����]�h�J���F��
�`)�@.�. x^�E蠞͗6+��؆�'�{�:���|�!�L����>�I�����4���\:�7"�LG2�^)���b4*?W�i1��2����*��tdC1���uMu-��ZY&�alйU��Z3ٔ���֔���K��nS��œ�:\�yn�T���f�.�HG��$mFX�,�۵]�=C�����N��i��1�7]�}T��ʪ��{�]}�~[�����t���43��{�߱1ӕ˩7�Ұ�M����|��l��������Au#eo����,��� ���ʠ�>�H��2�ǒC���Q���Y�S� ��7�v%���k�ve�8�eBF=3wC�i_|�ड़].�#�s%ז���̙�c� ;Ө��V��÷+�o�x����\ri_�ć7���x��X��]��' 2�M��&X}ε����5�L��r*�1�i���Q���*�4'N)BV������.�tH�H�)�k���j��ʑ<���[���y>�f-�"�q�Mu����iq��l�6ИFF���R	,�ZFH�{ʤ�2՜���F��+]+��n��=�:	�uE�ܥzb $FU	�g3̥:�M���ӗ�.K��b��a&٨zi_�N)Y̝����@����}AH�~��0f�OА��y�rǽ'��Rx�L�'������K��%�p��'�UȈn��^��hsd^{H���\ٝ6�A����*�����y1�0fز�x��!��7����3��8����9�sb �#9X�@�r�\�A��ji_r���?�)�
챬ώ2[lv�l~��U�I����qH#�U��Pu�w5xVe��Z���̴�K�T\�!�&')���؆9��d>T՛d�ߪ3J;%��4U]x�����E��&�C��Mr�S�۶��D򕇳'(�5���W=
�	�ɬ�a6y~;�Oi80�������ۛ�o��)����.��)��P|v�u��pЭ�ks@;��=׼��J#��\�VZ�V��&���y�7FX���8ޗ��[w�=�k[��;}m����3��9D�7���T9�nG�r����^a��~Q�Z2�Qj�\���6�LWhO��cf��V��b!��RJ-�I�γg)���[3�&y	Tŵ�]=��{,�g/Wr�Z �S�6n��[b�OCJ��� ǚT��H��0Dc��N��;�LƇu!�2��C�;R����mWb�-(ɲߍY�O�v��!M�n�Kc�"�����!����ǐ����H�����)�U: Cf8�^܄~�I�lL�YK�\:��ܸx�Io2�n�U�z�o�����eY��73�B���ZQ��[�}���q�x��-�z_�k?
���A�+	�����������6߼�v���c�-i���Lj�qZ�^I�oOX@���Vm�38n�}�w����.�RV��4��ro	�P
�Mf�r�@V��)4�1��o�}����pE��i�(��"��][��� �"�M����bG�0W��)�|J����[��[�4�;Ηk��տ��d�}�"h?�@Z�0
o<׍:,���?�\��u�+=&�����(���n���ώ��;�HN���<ڋ�֨Ӄ��#N�P:���x5�5��W�Tܶ{�iC���I��4C3��C����9&���F�k%��Z]<5��})�*�b���_��PW!Ba��Fl�a�V����/��a���a��s����,T�Y��?�����a߽��QK�=8蠟���yY����H���3x�wr��" ���'���m{	��/�g�/%BmRӏ-�=����*X��p�'<���,>!���d)��<���s0m����	z���Hxƒ�`���lj��W�� $�f�s�����	����؇ŶM�LX��
�������M.]�&�ݽ�D	y:�����S��	8v{7�q|݅���7�I�0�NW0�f�rs�A��R�.zQe�jb������4��ᓞ����ʡ�9��{��4�4;U������5��TP'	�C���!fG?iH�"z	�TT��O#so���������vD@_��%�Wn�9�=�!p�Ú��MN�^\���'�mZ,���#됬�@�K.p<���B=HGU���b���g<GH�qu�2�aS���}�%U3n�$Kc�t����;锝�B�~�����b
@I��Vk�}��-��ʗ3�'?���F�\x�w��V�o9�����u���y��㛔(�~!�aR�G2�w[P�F=��G������\����������~UBU���J&_2lY���-���i:~����섒��)���&�"�$����֊~���SF������=�|���û���r�FCs2C8�@��L:l�|�Ϛ�%,�پ�`u�����f�g��e�X	��V�ip�1y���)�g	�\��\w�H+�T�@�	�ӻ3�
{8�C���D�L�D�Fk���Bm�,����!��)&]�8�Kǲ8)P*��a�/�
���MzS�O5��>�6<�������\$�(��F揇n�ͣ�H[��:��G珅�Ht��E��J�{�7������PB�u� �0�!�QNY2��B~�������5ax£#`i-�~���)�����7�)��P@�n���{��ݶ���R���c�����o�,3�c�I8�����b�1�
m�pW����@:�XIv��d"Ȕ��}���c��)�k-�U�8�P����P8lɝm�ƜZ�����ً7�?�f�f��q>� w+�M|�b(�~����ڿ��2���(�P8�~,� �����~�C�����Hs�羱C���U��A�#m�.H�2+TU�8��dЍ�Dn��6�=A�
϶��+�W �id����<_��V.����\^}�����v��.h�lzB�O�y����ព#��v��wt�6İZ������ղD����Y�(��������������?�+�ݛ����mi�M�k��܅�ݳ)���1�9Q2�%/��m$���ڛ!�&jй�F6�������i�B)��}��^+��Wڴ����܄�ͧ	$�x���*���昰����5`�m�ef�O-+�@d��%�`����;YV}PF=B��{���/�}����TK�_q��nN��0���Kg�@�j�$�u̐��(�]���HeF}�D�{��]��K���F�Ӱ+�vEDX���(���S�Vt�;T܂��X$@E����H��oAC<γ�=0\��,T"n��������i9�Y���?X���"&���ù�+��s9t�+�"���M7[1��K�OYI�!�]�VwWt�Hと��ǌ��1=��{�O
���*���=}����4����_��{����#��S�?���<ª���^+��.��ǭ�� 4|Ӟ:�ΐf�KE���h�Ւ7���X.'Z�ź��̃!�C6_H�MK�P�i�qVﯽ���+:譴X'��bi��ͣ�7Y����>>�4�b7PK�B��^�GX����B������O۸B|��� gq+���s�W���V���M�%Đ&|K�#�,���.��Qq�hpRR�q�'!0(��NP��W1ՠ��o͙�Ց��M�+lD ��u�n�E������~�d���!��:/��������E
8��WL}���L��*�64^�����^��h���ʂ�	8:�ˤI)D��[���mP����5��ф���q��ޗ��-�8*���"�=�2�<ƛ�>����\�ͭe�����{T�����&vi���d�
�����g�#��Y����v3�[��T3�v���|�Ifb�4?�����.��ke��8#�:��kg�r��"���WV@'��^�����Y���6k�*:�HPq,�fRf!x�AY����H�	%��{����+V |�ZؑR%vJ��ח����8���[�%���6)Q����W��\�H-�)�*<��)|j2ɋp93uGS���m����CT�CT=��BVO���9
譴d��2���y�
Xvb8LO휑O���'ے u�%���bص=�^b�J�k���X[i���l�6Ѹ�h�!������KL�{oy�13�v[gNՇst�%}*�WE�7!K��=����X�-��c�����y`6�=J��x*&F�,��ą �J��*�@���y��|�p$�Lo=�ͧ�kEN*�"� �ߕ=�-с���l���]����΢:F9O)K�R��R��^��_P��ocj|��B:-72k�p�>v���H�[-� ���3��	24f��Ù=�g!,�����!����^Kxl�BPI��:}e�b;M��<v�LX�f՛%�4���wݍ�=r�<�Xy㩕aeW��e��g�u*�!��*	]���Ps�HCT[ϰe䛮��=.�˶JOÿo�J����"���h<������
�nֽ��gƇ@����B�ƱR��p��Z\�ϵR�)�IƧl$�c���ˣ����{��O��h�Q�g)&_�m��UF1˙��,�%lQ
�%%O�(��){��_v�<�l�����A�p;���@���~���!s�{Q�V7���FX�H�f7Cs��#���w��0����|�!>K���Պ�ò%�+�|s�/�Ţ8>V�>^�=9I��MS�L� M�ʹ�KY��=yD�Ƽ�����h��-^���L�9�q���dҾ���)���s4��93�q�x�Ơ#�x"���`��JKCA�o�N��]C�5H"޿f���[U�����4�3�N�K&m��vP����B�v?}B��!��
ܣ��#��$�$8k?�1;�o�Ȃ0~�P�����Kq=�ߙC��[�s�9�B�$�М�ѐ��9>�}Ak���`���*E�^����	��z��h���-�-;C�Cd�v�-)>:<������f�!'����Q'D^9�!\ٯ#S�d:%R�[��W1�������8�e̵0먊�݁F��D죿�������'Q�|�(�f��o�_�O0��J��(�ub�Ϧ�dȇQ����II��_,0�z�|�N"��G�B�73�iV��Q�<,W@0��[�O��ւ�6���_����9��0@u9�����1�[�rP���N-Is��#:fN��IHž��A�/"�:���֕��mx����$U���QAY-���z�\�!�������!��a�\��L��b5�U6�� �m*G�N�Ex�ʠūg�HnJ�����ÜQǪ1�%��(�wN
v�y���@������؇�	��&U��P��J�?>�������
���ml����8�ޡ�����,ke�(@6�r3����Ϟx��~��q��s�����_��J������t��X��\ط����d���~��2��ř��L:?B��Vm����`T�Gh=��(��)1Nu����q��
3�$&��������t�3p>S�&_'�xj��c��������l+��f(�Ћ5EM}��9�NH���$ؓ��{�[cR��,��L����Mcj���*�%��\�	��q�C�T+r�2�:��G�cۯ�M���t��I6ԣK.J����5�?�q��5�
ҏI`���w>�,�ꍕ��J'3�'���@ߗ����Dk���J�޷|�n�}�I����q(|�!�f�\��(�O�@^Ut���Q�ݥ�aQj��2��bu�xL�R�[ >$CNq�Y�,>�oI���I��7��l��.�4o�M�/���ύYkI~U�+�O�z1Qup�����r��wo��8�t����\��pTBu��T��kDe�<����c�� �{!���H�YC���5�����%�����bئ��
��.=��S�fq��#E�����88�������81{�歷]�� �g��&���&���!,�&���]v�ݚ���wͣ��s�zk�	k�[�K�)/=hx\e����vѕ���]V@*b��G��e{���9��:<��j����4r>��6�C��jT��X����C�M�ʶ��Nvm�+?Y�б�ו�e@�0'����C%F���@:��k1�D�q�uu}T��l���֙j3v\9w�ؽXD��묑�,?�!ƥ6o.�
W߉	6�����dh�w!�Mu�?�+���K�S~�� -��y"�JX�������UZ��r9�-��y�Ӱ�T����gC� �Nئ���
��j����߈�L��z���q�&3�T[_��/(�f2��Ӑ���#�(�}ke�&6#�]�pm'&������J��/��:r��d'u�1\�ž���T�\��$b!��M�|QŶ���*\�Č�s*����R- m�GG�<r�����l.����2(ulN���1�+��|Cbr��K���N!]vKis�/Mk���D��_ �~�\b�y���΄l$�i������/�w^���>�
JD���
��{�Tz�����[�ws����t��}��{<Ζ���d�|�T;9I��dTߦ˦M��Jr��#�˳�Rq,�#F?>���"�Z�
n��hb��{��#�I؉��'7��8�	�C9t�ԗD��Q:�к�S��իf�{u��&��.�4湒��Y� �i}��/#[�m������F-/�"����/e< ��?Ѿ�c�vL�M��J�����41w�'?QN�ױ��iU�&�R�C\pZ��)���OKп��7h!l=�ukq��^d���,'����<j$��%>�#�%86u��CV��4[1��o�E_
�ԛ5�w��=u���BU��/7F1'���WL�ֶ6զ�I�,��#�,���P>�-����mS>�Ύ��������]|���T��0�'Fs%;nӍ����K��կ��]�rhDbՒ5��!?�m@V�8����U��J��G�c����{�q5˪��i��.Dx����w����tU3��t�`�|��,�
��U<�(�=���HbI4��*�({�����ֶ�Yf
��t�w<6���I5�|
{Q2*>�L�ZEjf���M/�[�f��z'+es�Q�v���EY�i�Po��aCS��t�H޳�v�*� *]2
c��l�X�=���ˢS�
D禶K�B�F����\ 4���5������1:��ӵ[��Cb��ܖ��c�p}w����Կ��A����~��|�����l�5#�W>�^Hub�G�7��=��lw��&Y�T���?��"����˯��3f��ه~@sߴ� N�!�B�Ƴ��Ț^�жU�h�
&�Mѻ���ܸ�T��T8��]*i:vw�H�+Zɯ	o5�O�uz_ЪHIߎo�	V�(��2�:���7f�޿4��d���;�z�A��u��?<Ŝ��t�����8G�����jk�O�u��ğ��9/��?��9�z��!P�����O�jXeøSOz�ə�ʣ�����>.�.��	�f����)�.a���O'���@u�)���6o�ٺ����a��x��i�����^9�Y{����"R�dǿJ�._��ӂ*X< .�����PI��h���K�Ɋ�e��24a���D?�/�B<qs�����Ɏ��2%�ve�TF�7n^�l�����;���ނ^/{>����rM ��Q�����{R���Iu���5R��P4���:F�o����6��7�+�$�Oi2rEn��\���K &G�@#���������8w�Ugk��X�&���}9s��٨r���o) _K/O���q��F���RN)�|�BE4�����IK?�\��<S��I�ܘ>=;_o�5�w�:b����l);jc��؁���'	<�c���!]��n�u��х,��;��.���x'l�U��>I龛�	f$Ʌ�D#�	���bVO;���N �Rb��`q���q�AQPz�#���-rg����ř�z?:6+ ����Y�Jb�F��,��8�e�.l�I����|oǢ��8[R�P�"���qV'�C^Dwl"����("�%.N�bs��*R���1�¼z�z��X�[�]�Ђ����';XD�/����0�B�,��GXoV��1M�%��`���3��֫p)��q�A�������*cq�}�d58�X ���l�Z��2SSqA�s&%,bv����U��E�/���,k*��׵�4a�_A�6�9g����U|���5u�&.H���5�)u��?���,��X�e����F��9�?��A�����Qsf�����%/�}W�	[_M);}8Q>�;�Mf��,C[����T�Wɖ��;No{֪�����Ēza���k��/�Dk��	��cٞ��\k�	�����T��N��e�ľ��~&�$�/���^�AV>���گ��\|��S^TQg��jo(�W1P�<��٥>�-m��������Ƕs7QB�����7�����*��b�*n�y�`��}�}9�gק�Ta�$"����
V��g��E�s���bG�gM�����	QM�����`����}��&�4Ѥ_��J�^i�U���{��@�s��C�L�C��_̀�م��v~�k�(Y:���'��=��-��)�-�\^g���s$ $V/:�M�U�D6�,�nY���\{>Qa�)��%TU���p�G����T�d�Dk"�Y�貦��6�X��T�R��o����2.���VdZ~��k��P����
��k֔�0W5���[F%T?|�?�D�hn ~��Y�w7"�KMi	�L�	�f��n>�ӎ�3�C@�=V,w����<(k���'m|}�c�X�}s=�Wj�:ˑ9	��;y<��G2'���U��R��oax���� �r"��A��M�=�^z������m�Rz��?����ig�������W��<�}>^���23d���-Lpz���F� H�U@�5�`;'+��_�q�p��}QI�����-�{��rv�肋V&�?ϧ���*�EJ�ʃǺ�:�7�6�1G����w�q`��`������BP㤕��`��}>G���#h�2Q���U#Z9��'��6jN�����ysة&)^�j�q#n�.�Q[�Yf�i�^m�{HC�0�(��+��τ�q/w�4e��4�=}^:��Y>���%�ʇ�t5�4��Ec�ƞ���@ҔӀ����;�1��+�OFgG�o���}/�:/)��#1Zy�A1���̬�dz�������.���@MUO.jO���l�z�2!�i�j���Z������|��9өV����M3Ϟ�9�VtvM�-UeL��$��z��+_�������w���c�����w�'H[�K��Cԩ�����ز�:�pbk-"ᷤ����D�&���s�@M_�@cm<}��������o���%��[�gP�͸�~��|ڽ�]>g_z|sv������!����^��\�EU��u������ �{DPb>$�c�bp�_�X��"�=[@~7i�j�ܕ�D���8t��#�:kZ���*�[�*��C���u:�_���n�O��0fj��b���.������ᗹj�gZrF:+���Ǉ'8�o�:1Fvy5�IIL>�W6r�ԓ�&�en{w�u*MF�}u��o�53~�S3���^��trbUo�q/z��Z��g��g�*C��LѨ7aqSY��_�6^����ݻ��[�\m���QoM�%]�����c�=���������4�Gۿ���#d��G�R�k�;�BNhE`�z�A��;j��d��{�>p/+�P9e� Pqʌ��U��!"��2��n��u���&xn�z"��H<9�T�Ǘ�W���ʝ��C�d���?� Y4g�%]��\S󠀤T4x��<]~>�X�<����6�&&Q�%Fp�G3G�x�m7�k	��g��a*�X�)i������u�J���9��3At�(�`����H�CN���3�v�<V��\/k>_j�)C���x�A��|3��RIG���Y�hh�g
x쳶@�\#E5fv&�@���|Z���#J��d1��t�N�k�ݡ��uo���
"�L'�r[���۔�W�5�sk!Smi!�ǖ[�O�&�XG%%x+l��p�6UY7��ӿD���H ��Ќ��!�d윟Z�9+E��'������Y���k򟒨G�pۨ��f��׮c��n>5M�w�m�k��O׻�PS�?jR����6����zs������(Pgzo�'Z��;�Pb��m���\s���G![�%���(����.
+����P�������n<%m��9k�p�G~ r�<,�#L7��)u`p�
B�^}��R�(��U��i1��%κ�ҕ��e.�\���@j����,��>���\���N�tJ6����>�ڹ��5��
���R�Ƌo=l�aa�T���X��Gۭ۞�����'����O{>N?w��=/��@�ʚ�I�X�G���"h�"h���������N_L�b5���>�RR�E~ )�v��N��d��-ih�L�9�+�Q)o�b�Ͱ�j�6�B���xv�a�M�,b �M�ۍ�^[�� F�|��A�ns5����6�41ad��R>2��~B~%vBL���q2Oo�[��,�#�+��B>q�ܿukB9;p>dG��X�M�:c����o�F�N�-�ߟֶ>��=�M�����Z������&+���"�̓�}ݥ�$�}S��E�*8~>���bЊ�Z�K��=�1fqljX��:O�Q���x� �:ZB!���� ������}��D��Gf�,�/�o�����ڤ�,[�-Z�8��K%��]�=a<���,���W[b����ՙ�XFXm����j︎:�6v�1
��x ;�s7��I��:� ��;f��T��y�\2MMS��(.z��f�D��*�˙�$�M�	5_����C{�{���Nȡ��=>�-�Ǌ�,�3����]�O6D�ǋX�)>�W�3\�l�I$�(���6���./d���O���4�H��<�(�~�12�/�%�[6���{���:Ij�>�+��e�c�Q�i��)j�X�{���|KD�'�I-�v�"7=p�� ��QMr�M�����}�ep��Іm ��)X�W{Rv�Bil�c�Y�A�>%�S�h�5ԑ��T1Ħ��V���_	�>ڹ��� Tv�w�``Tf�'g_^�{Ԍΰs_u�����NUF��5EMAЍ���v�/��Y���1�K�n���0�M�ps�'�?|�z�1b�^�]�R��/_TX��`��S@],��E�%�RT��P���[��<�af�I�[������٘�@-��#Kf-�dF�
hq ���ԗ��m�����$�M�	F��zT�K�̒fM����P[V7��Y���}��҄Q%�X����ۏ{�!~���˩JU����A�����O��f��斮�iI`�?]�G���熖��ʃ�P�%�阔^�%l����eD��h�A�|I6�J�n����]�$��i��_��Z2�5���A�_��_��bl'O&t`R���5hm��t�n�b�|�������t�7�Ě�B��cрl�i_�$�G��"o�Z�FrR-`�y/3�be������D,=
m�Ձ��W���@�(Z�?�1-&�C�]�MF��
�r�8O.���\"���kE�W�eQFp��B�>^Aqh��]'�XTT�bbD1����j!ӣ�RP�+CJ��S���Q�x�\�����	t%�����'�N^�d��y�H'�N)�2����:l��ӥaf�J�	��߶eQڗ���?ٯs�
�~<`?R(n�5��Ͼ��vΓ�ڝ`͕�4�!�$��L>3��[�T��`%ɜ08�,��LYkJW�A�%�}�mL߲�����_���4����E����S�T��6փ���/��3��Z��z^'��&.g��� ���E���\�,Կ³|
�,����#��&$p��P\��M����K|{ħ��Շ��(�+|Z�(bf�7��ў����(.AQ8v�q�0�GtQ�ǯW5p�t�[=���Y�?(�ֻ�I���r��VE����NR�X��ٗ�$�U���R.��%J���&��}��p���kRޑb���W�����٤q��Fc۶�ƶm۶m�N&�&v����u�|�5��f�G{�s<�8|^���da/��,(�cQv0�!�Pr��$�j����2��2>�17T��46u�����|�q��I�k_�c����B�;]��}����Nt�%E�x���{���h��@[�ێ�������`��p�Cշ��<͜$�(����,�Mw���k,���7�+��������Hxw�n�H�=�_�Y�ٚ�I�/-)��N���*��ou`��x�|�2��=�db��8:�e���3��m"�w3E����3���9=���%j����3;^W=}̄4��} ��ԿIoק��8'��3��B�-�Z
�RD�F���[�z<zT�Ԅ��&}/�ܜ* �|n��3�E�;�#�B�I����*]�lܹ������u4S[��$W��6cL;=�c�#���4ѡt�ft��n6��W,���������&�㲿�skxق���ī�'@h�
lgifq;xf���&!���G� ��.H%����e�=x��1�H�����h�j�o�����3���H����������I1ƿ$�u���������v57wŘ��?i9ZP�� ��med/Z��_(��g�H���»x�me?�Ow�"�J���3��X������w���7�`.�I�Y�S�sӥxH��l5�(��o/�~�W����f2k���v���f<�G>�["ʇ���|4�P�N_�曻krh�ݘ�d���Yj+*Yj�b/��d�UF��T��A���!�#����
?����D�`X9ԩ
�t��NK��䀆�!�Kb��Wa̜<����ƾ���x���P�9{������2@�28/FH��r��:b�����v��;<�p�1Y�^�l9��چF�d��TP7 �:�V$`~��[LuW��R[��3c�a��
��rs7g���oW{t�7*�H���ây�ȫ��1���"���ώe�B�~��*یR|P�a� ���C+V\>�궺U$SЬW���i���+����ҨJ�!H�4��M&�x����w0�]�|�;Œ�g�M�O�ӹ���KS�*)�ܽwUӶ��7TW�$��v�݀>Os�vo�mFXam�g�4��z\��0�"�����}���j]��(Fxy��:�c�T値Icз��H���L�􋗚�+������[�ŏ��M-s�G]9��yh)[��9U�	�6X{&jß���\�����?/D�2 +��0���;d3~�K��P������J(|�������=&7�?���� ^��k.���������s1}υί�i��i뮋���c[R�g�N�w���ؠ�V��q�_�P�uꮥ�؊�9}YR��e��N.uk����98m*�`�J��W����kW�ntM�=c�p�`U_=d}�������q�
�?��a^[��A�
U����>g3�
���U��G+3�r�.Q(�!�^����7����j�X�&����YC~�������_`�^Ԗ�\��A�X�($���e�r�+�����^Ɗ�]����('� r`�z��g��I:h��&�[������I�'陶L�����`��Jɳ�!���Jo���:x�d��Cg$����+y|�(-s\�せ�/��T
�q3R3_E��{ɓ4�Oߑ/5u�2�l(ǉ�'��ޑ�����_uvh�l�+�J�ˠ�K	Mi��YIa~judc��6@= ,V���w���ڄ
��)�n���G�U�V���7�����E���D���&2"��qZ��6���8������T�/��{��-V��eǱ.���'��o�T�����֚#�rF�*���a�TYuP&�RA��.7μ�r�5� Q
-�?3�M�<VrРJ�Nw�e�$~2N:�X��q)]�r��jL���E��4�_�s�Jׅ�K|a�eW8��k�>�?�0�����}�b�џ�5�����Q�XRs/-�1]�L�
���
���?�!��J�(yğ�~����f�s*��Vk��=>����=����-k���za��������}�z���e�/��BM48�G�R��;����&�0J�Dkq��b�\C��0cn�v}p�$�fsO�l�+�3���(�V�]���3�tW�3���𔽋[)�������v�1�Q)ݝԇ38c;OdP�����Ɩ��LMY]��'#�&�s��~��`��{�]'|��ҍ*�b��R��|
H�2"�K��>4̌$.0eL_v='��]p���|��!�u2���7����N��L���Q2�[0�4=q��G2t����1�v�Ь���c�Y���>�� ���E7"(��͜���b��K�~���'3�tRU�l��P�i;�ik3ڎ?�̭�ғ�~�:g����+fP8�M���Y��v��K��~}�W3���F���.S,_M���*��L7+���<�8��G.�H��>�"V�S�/6)|�;��M��k��[?p�,��J�Y�Eb����&����J�#�r�BJ�v7~{or�"�<��䝆���r���Rt�2�`�s��y�}�p^���Gv�2;��mo;=O;�v�I��,��X2��6Nb����<�\7g.���W�̐�&��GG��Y��<Vu_��^#q��"����i�:,�Dڪ��IQ�P��dR%�.x�5k�����D�sFN��)�֏I)����"8�?������/���j&q��)��脱,c����q�)jЫ�~���f���+g�(g�z�B����������F�r%�
ik-h��` �\n�֐���2�ܢ��{5���@o,��OA�����j��������u�?J���{lS�o��&�rd7N3�a�]��g@*���˝a�3~�,#I?��1~�j6�6:%D�^
PB*J�n�c��i�Z@��]P�ׯ,g^C��u��s����T�(3�,(��)Y<�Z����5}����Um�-��Ăc\����H�����x ���5l"I�L�61���^?1���w�w���E���~1V�ʵbe��䮩��8;ٯ|��^�����P��[	֕wߦԽ�<�>������g��Pq욬͟���4Jܴ��s1��l�9��&Ce�_Nx�D�sJ��Yf���]{�xTʰ�%:�D�lԴ;>���m,mT��8��}�pR	���?��ȕ4cN��.��7x��.��M����U*������S�[�����4�)�ș�/��2��xt�*�S�ێ�2���g ����봠'N>��{��|��|���L��R�_[>�?��w=�����L�Ġ�:�ľa�xz�Mv�*C�f`��C�L¦$�a��~Y[b�
R�D���? �(oz";�(QQ��'gO�ڣ�Y��d>�������̟� �q@�
Q���7�Ϟ��G��Ǝ��Ӝf�	������Xf`Q�/��L��*��K�r$(qE�eۄ�j��PQ��sc�;���ΒuC�ΫR��u�
�nonN�䮡P�%����������2���=O�����y����`��H��F}���ʤ�B��#��m�@s��`ԅ�Ѹ�)��8tBf��R����=«k��ο�n#yV��?��J�q�*5U��$e���+�d�E#p��
2Kb3�>�BW���G͟�A9�-ŖV�j���>����x������8�(��Gv��f����e��Lp�=�Sn�o��Z��/�<ȑ��4�UQ��Y����7/I�?�"ٹ�}����f�暸�|V���[�`��;���O9�������HU�d[b�ӧ��R��ٱ8�/Ck�7ӡd9�V5'�al�v@��gM2q��V��>(��*Li9���]Vk���;m���[�������*QD{�*�1�5-R6��
p�WjRu�5G��{ޙ�w��A0(�cq�%(�o����k9���Z7���9�M����j$
��km�,P~	9��E�L9fYz�dlE_R����85�R>ݮ,�A����{t�K�꒙+�-i8��H+I�Ҋ�F]/���(�6CO�*�ˌ^b���x��f*��LP�6.v��dM�!���t�Xg_����Y}�O���^~O�=M7��[Ag13q]��J���>�5#�Xl(w��N�X͋w�!��~�5�ܔ�c��`��~&i��1�� obݼ�'��Mk#�P�<����z���c� p�{������`e/X�)����W�����^L�h���d��bEG\�N�uj�>�.�b)幨���n+��|~��-��|i �L�3���0�m��ـ�<�,rT;�A�6����M˟r��\��cC�Y�����j�>!��f*��f����=R��C�1�Ki�ɭZ��f.N�%!�����ގ&�EW�����3I�ܪFw�ߣ��/z	���9|u���Ř��	߬�u�v��i������i��8~~�܁�4N��@��Ι~+UzM~oc~�\ �S+uя��瑾�CNv~B�	���UI�BUHxk�s��x<�mI'�L�A��oY�����u�\?�cZU{^�)9�>�=�J����_�F�ҟV��:''�&�ʁѯ�'.����W#�YO�М,V���j�B�L�2J��;���'�*���;G�%�,��N>�5v:��\Gp�[}� �Ta�	&�ƙd��9Cd[��~oٚ��n�̽�<_�Wfs�_o����nQ�̦��e��\G�s���m�w�씳�%�?�B!����XH�����$�$�S��K�Jj/�����J��{~��:�˥��y�n{���N�_�j"ﮖ������P�[n��g���Ð��v�c�ed�탒[���p�j:�ٹ�Kz��#eS�M�~�P5ǽ��X`�Иz[F	K��:�M����U�5q}HN}t�S3w�r�mIk�	��á
d'Ҷ^�3���o�lrR����]�V��k�Gi��Z�����UE+����ZX������Fbȯ\�]I�"��|J︢��*b����T偮�v�5�:��S�?���1kP2h��* f�~�����^���Ib�E(��(����q�Q����?����ֺ'�1υr��	��~)��@���eHC�,� ��
 #A,��#K�_*��|��A3K�^o9�qڼ�3S1l#�b��555!�71Wo����ݕ��W~��彏;��,5pl���VYy�P,����v�W�ڻ��[��]��Ψ_:�׎�Dm�q�pT'5#�H��܌�ځm����Q���9z8�����	'%�KY9"p��b�b�\�N��ly�e����sx�k�]Bk��%3�l$��2/nx��MK�^Q'�bWgl�K�%K�W�X4ڇ`w���@s+�
���Y�suEPS?m�c��S��¯I�����z$���\���g�����'������.��?��!�=�]9�P$~��l��6�`��+,����O�������jt�$)�B����AM���g.ڜ͵�5�KqP8�Y�k�ڌ_)�2p��X��V�ɷ��I|F*�8�JnI�
��9�nO�QL��{G,���ʉ�5ݠ�u^�F�5�֍@YO�H��:��""�Q��c�nL���@o�j�~��2}C�DR����.Q�* �|�x������Rɿ���&8���^�}���#�ңY���xϤA�u���~m��v�݉Ҩ�s�4��))Gs[e`��s���R����m�h©ګ�ζ�˕t��l�x�%�E]!:���mb�4�����sq(���ʪ��V@ga�1@p��^~�����(�������S��tU�7w��3�h塁���_E����\��>Ϻ��qm����U�n�.k�}��~��GU���즖[h�h�"��Nr�;�$�	_ҬQ|�V�֖Ip�c#�A�K�RB��.�l$�7ќº*$(��-����诅��sj��tU)�������l��B���nf?}YȪc�,�|,`�����ט����J�|v{�m_n��;��3K�Σ����vfD�M�2�SS%����U�jlt�9!���S$���ym�Z�!���r���S�ʷ&��/y�/g���L�"2��÷�Y(2ӑiE �=xp���X���0	����%%~|`��'���fz/5�y�}S 7��)��$b�n��w|A��@[�@�	��3	dH2���yŌo����^�:�����nȮ���u��l��&�]u�4�L��d��/��"�!���� ���2��� @�wvc�M��Q@J���6�:p��;3����dC�z�Y��9Z��=6/��Xs�(d��:���ܦ+�m�]��-;
��_��5��9W9@p�f�#_��=��L�LA�J�~�;3:d%r�C�KZ�7���R�"�h���*St��̑`���2��l���b �bުdT���J���X}��O�����}Tp�7�M͵�d�J\�2b��S4��V���dǾ��b��o6����.�����HK7�.���6d`�]����U�sծ�Q"��@-������{- z)�Gu���F����F�I��^�1/�$V�$)YER'3W��*��b����&d�r�d����b����҅s�+򀱍�E��\[��Ff��0)2D�y���nB�^{.z&���Q��bħ����5��$Q��i���1�jN�ʔ��*�X��0T��g���xjm�jA�/�����Kdu��/sm�!�Q���Ezv��9\6^[8ij"
<8���A GE'�$���db�.��<#$gfi+1�\'��6_]�_�L�N멫��˳���KT�yF��D[�E��d��L��eJm��,�$='�Y������o0yV���!�>�otD�Y_�,�E�J�)ez���OB�T�gsz��利�G�52�������{��:e�(�`����y�վ�:}>���O�M������|m;/[%���D[�m���Eʥ����'��e3�t�����~�kVJi�HKU��h��$�Pr�[�s�&�HbiO�Y$$cv�n`��df��A܈JT�n�h����iIlZ[j�}*��f<+�T���`o�a�����+�P��O�&_�<Mg�A�Ɉ�-9��D�y�;3�]�T=�6�+�4�<�,Q�o4���qu�gIU�>��|�)|��G�����i8e���*U�0Z�>�K���uI��ɽ2O�c���ᗥ���Mk�)��뺗��?�ٍ��^-��J���8�x��wֿ�z.i#�h`�K�A�Dl��r%Ŗ�|�S�</xrﮰbͧ��Q^#ʜ�}�67U�V��)�����5�`[c�WUe���������y�����'��`D�������W���a�ͫ�e�KUi-�*a5�Hr}�ޮ�K��|��j�|��C�OG)��J�F����M�Q�$�g���@l����"=�?�@-���� ��jC�����D����ts܃�gK`^�.m���4
\���*;��bӒ{�^�<P)�`���67�Q�[�g��J*��u�M�k q����o������D�h�[}����
s0Er�!�t����^Cf��i�N@��EWӯ
WI�R*�,~���.,w\c�∿~U-x~��R��Q�ߴ�'�CN��jz�0�`y��+��
�2�xm
��=���9��}G�ۚ�^��F'J�w>pΎfdmh�v��h����t2]&��>�f|dN�_��G8g��}�C����1�)i�C�����&Y.O�2ȕ{=^��i�P�F�AH'_�����Ԗ°�����&PӚz:�T	�=+�r�/���ΖiBȮ��F��l����Uy�8Vn��KW���f�f���������ڶ�֠&��mF�ܸ�! f�s�&�oz0����et��ǆ,g얪Fo�y�d%���n^}V���%��D2��&'�z�o�H�FI$�%$�������:�=,i[�v��3j�"k��O���28)����n;Yh_"�;���ӓ�ˌ���L]k�2ᵑ=�����SdzG�[Ls�q�/�Ƒ}��g�E�kϚO�J=�~$�x���Ԣ#�Uċ��r^��zH�A��^�M���(oxt�@6��vY�ej�~㴖X7�����L.:���"��Y�!�W���+A1���7��ټ��kN<dCV���\.�o���P���T�1�z��Hmz�6�u��>Խ�h/g��Pzظv�ʆS�:$���a�+w��c��]�����NI�G�;�d�������{��:��՗4��������5*8�X�+=�������6���}�<�M���h�
?B	VCc2�����ՃC>�'$����nM�5i�{N���_�=�� �'��1݋��_��?���(�j�U��(�&�}��B�����X��1q�K~^` ԥ�B����)P�6�@�*��iR��+=,��(m#��L��B��/Oh�P6��t��W�o0�6ȓ�2ɓ���;�=��Z�����b��f,���
��-}(��TA�zC#��IG�ٖ}��D��b/Vt <|Te��������lG����;���7��s���˻��8��0�g��c���fi��lkk�d+��{6��%����8Eg98/?C�y&�U�JR��b�G\g�1��	lR?�_n� :�5UX
��� U�Ϧ��uSx,cٓQJ��^����o��@ct���Dn�ބ�%l�ÆI��^>?����r�L�´�#���D�f�{Z��qݻ��=;͘��P�0�4��%u �+�����&|޿(]˹(�`T������	���$�NY7�»긜�|�y��}m�U�$�J�_=�:Ь�ڀ���O߉�hR�N�Yt���|T�:����e#(5L���n$s#�vP��U1h)<��
,�O{X*�o*u4��hMqsk����ư�p��~I�:�T�Y�r�TE����P{�1��A�Y�`�i������i�jBt�~�ȍs쉅�_� 2�*���T��=�^���WxZv�f�-v�`����=�þ��O6�:A(/̓Ց�,Q�>ݿn���fdȗ@���{{aD���匶x��6r�T-��������}L�%���h��i��M%��7�����"(K�&�5U�;[�:��e S�7n6�t_��)-(��8����ҝSk����:����@ɋ?�M�f���Q���zav�	�&Ơ������ѡ����)YJŃ�?-����]t,��w&�s�\*��b۪J�Q|�oz�nn#�%�1l_��x}$��Z�a�S����� ������?��d���n�lT��h�2I{&�Oㆲ+NVf�C�y��D}=�X?��Ք�2E�&C	��ÿ89p��������|�ʐ�%@�k���,v�R��5V�ef)�K�~)/����v�^�'�iTs.r$��tTk��[�Tށ�Tw�@R�)��-�=5S���{:"�Y�t�W0k����6V	,����B>�����0��d�w�_'U^XY �υ?������27Xw��jY��^��9*ў|�;�!����� �n5Ɲ���5UU��\^��x|#2��}{E��s*Te�����v9U���޺R�A�;�0�X�h��lt��|
cJ=q�^����bt<o���ױ�ȴ�\ne��X�>�;<Ee<�cO�B�e����
�(L�x���8�A�����msK�W������!�Ua1���2��E��s�����&�h�y�!\�)�`���J`�C ���C�i�d�j�D��������Uµ��g��e�@[�Jߞ�l�C�踷�K�C�P���mQ����'�lP������qG4�j���+�R���x㧼����&�,������ڗ�.A�p��.SOQ3|��&r���.��׌پ��/�����Bյ>0Q���}����s��Т3D����;cpY�*3��8
����u���5VU���0&Q�Y�·�cA���H�9��0�RR�wJbÂ��*��S�3�)=v~*'�LcLg��4��w*&�n�2.eg��8�4Q�eQ�Ȭ��J��4�'��H��4P� �3�^Q���Q��]%��?�Дp$�а/��(k�[:��Ә���}
�Gu�4|�cr���N �9D�B��#R�`�O�1�Y������T�rh�a�kj~j'v�a���*��:��:	{���5�\���F�0"�$>4B��׏l��t2xC�T�بb�Z�X,�FK&�qM^�?�F�ܿ�rn���]�~�dM�*�8�}͙0�fB��c�K[�x�9\���"goiD�l�cǴ�d%�yg��̞u5
[l"�0��S֎k3@����L!��~�����s]�������Q֤��͠W= F!{	V`�P�^���Ւ��R��6�S�B6��F ����D^Tñ��A��6R�R�V��|��"p�3�������k�D'�<�T��fU��������Ek���o\s��ї�u����>6-��Z��ՑA�;'{Urj�ؖ�m�Io�hOmJnq���ҒJ'CM��A�a��᧩4~��)t%�P�qk�6�v����o�c&�-|�$��X�n2�b�8���WN�B��Sn�F�{����Z�}ޒW�������8�f6�F�y$/N�/�E���h<�EyW��Vx�r�᭦&	М*0�ȦsTh�b[h(:��S��"�k��ޓ܎~)�C�5�>���@���
��L�����������y`�H쯴c2F-�����v�V��k����߃رʷ����nU��o+q&wh������6^k@ˊ/)(��:��:�3sL�����cԊH�����A��J99��D�?P^4��Ǘ(���ho2�[F�0�L2z��![5�N	V��CP�?2�M��t��a��=��~��p$k�z�*O���i;�JD�75~+%X��
OaR�
)��
��ニ���Kݒ�CK���h0�3-LEyK��aeB�����׋E��_3���O3�l�2x�ܫ����K?�F�]UU��ڪ�����^u�'��fi"�W�=㙞^���!�s��W1Lݙ���cM��t00RX|S,�$��{OV܏�D�c���-���Iv���G�*�V�ݛ{7�mgV�c��8�?��?��(�)y@L��k� N�lA�Z���i��]�:c�(b��R������./��̩�dd/r�u�g�'D�#W�.��(^脯���ht/ܖa|k�:Ǎ��4���-;�rPz�Ϧ�@�����c�����l�ׇ���L��(A��R��a�C׃�:�m�-�|��-�0:ߘ�zޟm�s��\�1�1�8q`����"��&�+B~y&\��fQ��b6����
��YN�.R�U�Z(�=/C�s�s��cf�zO��UOf�,����ʸ㈻0Hg��!_a]��~6���Y(�%����$9� �I�H��8�.��0�9A�[j*a<�����'��$�'�'�!�y��]9>�?-{<	�Ǐ�Bf�f`!��X�x�����R��>�k#{74�>�@���͍����8������"�jFnOVdt��8q�t=5��	��4�zD�p@d�g�m���?h�#�V�������dY	��,�'�rg^���� �Fq	Ȣ!���!;S�w�<q	�iX��l�w"��4*��=�0�vgK(HŔ����ր�xv�M��B��M�/5�� e#��-�}a�!=��.4Gs{'�#�����bN����D�h������p�]G��7���MeD��Z$�m�,��!��DlJi�lצ�)5z���W�y��³�m�Vu��T��f�ઢ��=��4���P��p���Exr^�D��n�Ui�����8���(�42^4�ֺ�?p}.�1�:7��s�(~�����\ ���o���'��ZSJ�D�c�PL�;����4[o�C��u,��6���Qs�l�^�i������s{�b�$�s�J�7��`��0.��q�[���o�u�2�mr݃��A�%��xZ�'?dm˹�����&d����Ĳ�%+A.Q�P3�~`��gX̉���`?zѡ�;4<��. �Q��
�]Q���*��-��֌�=�ϏM�z��ǐ��H���Q�u'�~��
�W>r�D|tkaI/$�r�����nݭ��/��:�A��٪�3�d�������y�L��Q|1�k�o���6Dqˠf�u404�ؔ���S)����͢�UG�jD���0'3�zY^�!���9�d���a�}s���ǏN*��U����q_�%C�o�F��>6Y�a�{iB��#�)Hy̗t<w�3>I�Mo����-�ML$\V$�FxE��8������R��P~�e	�2�T���g�G�v�����������E�S;ÊE��F���߆����A��C�GC�:���a��`!ƤU;��d.��v����9��>a������]�\yy��'�+�{�������%N��Z���z��<���Xٽmlf�p��aɬ�Q����� ���ٚ͌���C�u���c��x�ˀ�_"Q�C�AsO�� �?N�T��Ǵr8*�S]N~iy�����Qh�-8(�q~Y?�XL�#tmgU�vG���h�j��g�ծɝܦ�ԑ�}��������_�P�/Z�¯6.��xR��~�+ԭ����ߏ���@�r�p��T{�+�x=p���a#�����oX'��t���{T ��G�U��ΘV�M��n�}��'��)L-�de�3�[��V�j�3ː����}�VxSݎR��6�<�Mck���F;c��0�cI/�7S�w���Sclx�	k?;������ճ���Yם)W"�皞�e��<����t
���0r8��Ŀ��l�5;� ���
�j8�u�^�vvtɡ��������}��q����N���Q�Ķ�ໝ�P�bMS����йMG��~t��1��ɯfh��dN�������F�:+���M�����s�5f�w��Yׄ��VwÅ�q	pvW�PNX�~���y�
�#���%Sa hKy�� x��s�(\�s��I��N��:�J�]�!5�r.-�g*m���b��0����	��^g��l��rU �wY�����rz�M[��Q�A��}�����D�[
���Q&��>n˽���HU�
���ZQr�΃.M��1�/�Չ�ov9�;�W���8�V}n$��!���	?� h�TҳT��s�n�6'����s����i�U)�G�A g���P�� LH��3n�$Ő�v]S�0?��%X	���v����G>�V���8������Z�Z/y�c�TrMy���R:�~1�aޝ��M@�X2����$��ů����1�m��֊N���Tz���� A������Cb��X�d�C�8�_���|"t91����H4K,�`�lY�����:w�jF1��Q8���S(�R�Ͼ������p�yJN<n��w�?\���A��<يG��!&��.����8,x<��
�-[[p�>��^7��Aj�
�����5��_(�����4���s�~V�}�����������[�t��j��Y�|R�]q��/�8�h�9+�hi�����K��?�7c��ږ��5�.<X~��6���&��@%r�	2��9+��޷vZ�,V7���T���yh�3�oJc�Gl4�{y�d��	��.�I#���6�`7�Hh0;׺���d��\�)���7�+�QQ�:v�1��h.�Z��i[���s�/���/�� ��ٿr=��uވ���B���z���	n�N��pM�z4��p}]u���t�Ї�Ϳ�%2���i�|$����+��nu��<	��q�˂ѱ>�+;�	�K���e�����R�J�$�
F�9Dճw�m(��۳n�=#�]1��1RY�8,�U������z��O��q�`i������.�:<��GC���X.��LO}l�#���T�&�B_�i�#�M]][��]�}���������۟�ج�R�N�L�ڳ���A���y0`{O;�*�J�sp�6�e���f6�%S�r����;&�[�:� 9������V1�O�X:�z��s{[��J��
`�;O�[n�s���r�;�=X�K���'z�Q�a����
h8���H�"h����<��9�	���?�z"A���7�VV��[8���/��!������Q�؋�tG�M���ƾ���������I�H��B�{�U��1��������ߞ����hW(�A\�%�T��k0�Y�e�F���PH�=�i|��;!�5!ؖ�EȜO�'�ih�!G3�d�X��x�Q�����E@�X#��L0�pvZp�:�覍z|��rY��I�C��u�t!;3m(��$�cU�4
��x��)8�?#E�(���
�(��xk�x�uTyH���'���QS�����'}�D������h��%�T�h$,J [w�of�����k���6Jt0�H�圌����G���N��Z���ՍV�j&�9�5qQ��%	�B�<���)���2t���g����<����<����Fɹ�a��e���P����j���i�U~��!�~>�Ǻ���=���*(�,��q��d��j�	����)�� UO���D������0;�e���Ŀ�y���Bb ���K��j!��Ij��Ƅ��G���kp7��\���.����f���v"� �r�[?�u$TRH^�K�TD�BS"~�ή���[�A��mEo0�~5�s�]��:(����5B��nY� �J�}{6>ͩ��u����]�E�19o�жM������s �_���ѫʳ}ΥU�IB�~�w��Д:�1�ϻt�[�@�	QАN���W�Y]�Zk{�4��x��ðh[��l��y[x�r�N�c������1G��Z��_��,
���~DF���\��6Z��k2��^澓����{ʣ��fwjX��eM��t+���������O��ԍ#<���'���u0
����K\O�������=�̎�%9�;��&=	=r����S�%C|���#�[�B[O8kb0�|��#����"��C��w���o�idUs.�i�l�(�%�Յ�5r���>,�ͦ����A��Y7-����_�&Pq��-�+���h��
h�#Y6Q�]�~�ڜ��������2����ݾw�q�E@��s�%��!��]�}�b'�G��H9�SBsS���y3�HXD�MCᦽ���H�f��h��yBV��[�\�Ť���T^l�´���eͧn�¨]��������$��B�&}��㯐���2�|v��4�C��"�}&�[��|���Y�����Lh�Ў��Lأ����V��#�� ���_�d��ۧ��:���,�0�BHDh"�� �$t��]_,��H��C7�7�V
Xl,~��{���E�\����$�(m�}��(a�(T�$1?G��&�5��h�P��3e=���us�r8z��8�Nk�tĞ�,�i��u>�:�Ӎ��8�ޞ���>�!w�|2��BE�R�^��>�1��Ȥ����ä�ҿYm�}�D����ˡFo!18�ױ����M�n$4��w�>J�y����NB2_���{R�,{��t6�0G��hc^�+O����u��k���-�/�����/2������HX��XC�+�V�����P>U�e�Qg}��������8���C���Q��}�m�<��$���ǣƄ�i��E��%��T�7B|�f��^H�,��V(�-�M
�4�Ezb-ԔL�Uf��4�7��G�X�D��az�9�.r�x�Fj�Q͏	�y1�����)�Tv�������!�`7�K�[�O�*�
D��u�y�k�d��u�Q�g�cOGYvys|����
��}��u���F!|���*�Q/��wd�k���-��7�SE�k��D�����x��������|_.�DݨN�6��3	�æ��띹m�rEV���P7DLi���:)�{b��7��Is��X�|ZF��Mh+V�	�Y2վ��ľE���b�b�6�>���`�<0a��Yl�m��~�����Mߣ�&��v�`��֋B���a�+���H�(���������_���|@Ґ����;�K� r֛�� �]���t8��
���Di柑D&6Z�@�)�^��{�xC�e]�X�F}�W��	}/�#^��
!���ǰh����r���r��G��s�;�*���*��u���� J!��.�N����2����i�|�+B]��bb��؆G��0)��4)I�G�IL�e�����{�矱<r0d���g������s��P���Dvʾbd9�X'	��)e)[v�X��,Y&�(�![H��e�V��!��]c�>c3����	�߾�/����~]�s���x����`�y���NZ�Ww�S�e�l�Yۓb���p$�O`K�R�-���^k���"Oɻ�qW���[|�{cn�<]M�U�uto����+=��HD5�����(���@=&�zP�X���s��:�7>@��=���:sҲ?�1{1�[0S@�L��l��-�:Fb|�(��͟���uq�%7h������xо� ���<�=��e�é;M޸��g�ݕ58)�/3������$mɨk�%�&U7ٞ�d!�
�$��u�����(�zu/��dv��h�s���l Y�����ˣ�_��?ڱ���bvx�VX0�^h�⠆�e��q�|�D�|fʧ�Y'C�x�@L��T'�Ju�,�:�t���>������������VQ�z�����|�ญm��%3.����ק6(8q�X��*��ዑ(?���:��H{���M��<�e�\?첞��Oq�Y
�:���޿W�rwD��lp�W���doց���0����l�����U�e{S������U+.�[��}BҢ�C�%Obp��vZS�F�N8H��&�I�O����l1������[s�4Lx[�2]ō�R��R�]V~fv�r���w]������S��)Z�869nuځ���y��l?b<�=o�w��<z�c�(r���Sc�4��x]ߴR���P(��)8�{��n���L��t�.�
�鑶9�mF�����������R���<�6�P(P��c�Q�]ւ��;h�O���W�Ѱ��"��
�5T:s�%�`��
/z1_��sw�j�x3_E.��v_{�Go��)m����^,����	�$��ֹ�n>63��lnN�y�Hd��T��g��7��^�c��PN�_��s�c�}��Y�[v�W<����%�rc�b$l�-�1s����`�1,�����tyK�P����W�*j .��D�r�'L���dN��X���y�:f���x������)�TH��ө(�t@����뿡�J�Q)ޡi2����1<Қ<Ŕu�%���Ԕ
���)}m�
�$����=�)��F#�!��;�Z�O��_��,t�,�Y\��D�N`I�@�Е��Jr{��[���j���G�^zi�ݧ�Y�/S�^PS}}��9<����FiLt�fL5���h�����iՙ�������!��4 H�xq�moЄ%+g�^���c^u��Zѐ�	�h��45��Wkbp���r�h�	J�,�A���<Փ�0Ie��d�Y~pW��[K@O����c��l�Oާ���G��Q�!�*�Z�_��Ĉ=L8��Y�)�G\*oN�}c��>H f��N�XԤќ�t'��[-T7�֚���j�>�D6��{�����ڣ��wn� @*\:9J����S]NTJ������)�gn.s;���ƿ��b��ҽ5�}�Jb0�I�N��;³����n�b�~�ZR?��N�4n�i��� �%܌�7p�ʷ!Y �ƅ畉������Z�yR�����$W�����J��AS��l�R��������{�Y��杼iE�F_��>�c!�e�yg�xQ<���� ^p�� �DD�M' ���{{|$�tG�7���K���Ắ��p'Z�R�H��DA��������̚�
t^h��f�����*~M�;j��2�v4+�����r!	�nU�-��-�h��Ѐ0������s�ؖ3 n_��R�~|$��ƌx��w��������/2�s\�l?��>�\Q����D�4xɖ����� ݃7�x^DR�_W�/Z�z�����g�$7~��	ٚ�����d�SZZ
ٷe�b�\d<x�x��U*��mih3�;�(yS]}����J���,��v�QTP0��aa�5@�U�> �c���?�F�:V��c���V"��j'����`�Z�����̬�j�>��RE<<T����]�U� ������a���/	)g�4ƹ*��Zf�9��Z�Ly�
G�M�b~X��C!<���܍�Dԯ� "'b$��|P��2���kv���4�����xd�u%�oH�G�&���w����������ޭfҭt�0_�4����Ʋ��3qº�r˹f���]�V���Q�;���/ŵ������9s7����57�~���i���,jܻ�h8�|�1�r���|Zlѭ������I��w� @4�f�7�X-o���oWPn���Dm��V{������ߕ��)$'���k�����
^G�	nF�X^���B&FґOg�ջ�~�.<!�Pd�}3>1�ަF����}/׸��*4:"S����t��Cq�%$����Ro���I}.�D zw���i��;� q88R� �Dz�� ��ťu�����6��C{����b�J�2y��z a�|���%���8��+Ӎ��|I�p��%7# ��[��AH�,�dg]!��o��'���m^�QC�}]*�]��x.g�X��Jh�5'H�ʖ��Ѿ�跂���5�>vS�e>�w���D~��sP��1�*J��&��E:��`=0`���]��ѥh�lQL�낮`��E!����2|b��T��>���ĵ`��b���j�Ǯ��-Ϧ�b�I>f&��'�/dHڹ}���j�;3��5
S���	�2e 8X�U��5�K��2l�L
Ox���˘��=8j�y,��9�/'E����*@�z�$� �Sǩ�a�*�z�%��SԞ	���Gv�����1�b3P�5rHއ՘�ޛz{�݇ �BW��Pvդ�/�ʄ���$|T;S�	ww;h����F�ݓ����ݔ��Vd��Fy��?�pp��>$/V��U�R�6��>B����*d�9�^Fl���~)�F"�%K,��	H3���w��c��?��3�_�0`8H�a"2yxz>�G�K�)�r��Wt���Y��'��Z��6a�X]��1�9���Ï=*7/��Rʈ�!�_F�$5��KJ�ȇ^���k��yn2��л�.��0�U8.��a5��+���S	<�q�b���ĉ'(.!H$�)�3+����R{k��;䣽�Iz԰㨓x	����*V��w�!���'���n����[.%��r~�� 	2����(�l�c~q��~�6d?Є3�1�3o�$%l��*�����9�� ��*�WLP��>a����|.�(�g����b,�n���x��`�f�O��FV�J�[�\q=�pbk�����%��y���B�8�gH�x���Bm�,+$!�Nʯ�U7�6P[�?P"K�U��&����� �k&���-Ǵ|l�)�|ʻC��d��4�ϵ`T��Bo�,���C������ԟv�4*Fm����=,TT=��X�i�����bڟ�e2į�cܚu�#��T����Q���H�i*�S���4i������8���еgH<�󑧸��ޱ��vڠpmng͇*�K�V<�*�:�N(����C��7fJ����H�ʲA�����l�b������n��ɇ&&j�x�w,���+І�ҦmT]�����Wc����-������,�ҷ��N��h��IS_y�r|5���&3\�\��ثߴ��R����o1Ł���z	R�i�#��-��?Rʫ#`FC`�c�~ʐK� C�R�{�P[� 
�)s[m��g��^�F�A����u��PI�bKޠ���c��qC�;S�LK�aI�kR��������jJ*�J�L�3l:��uF���@�'���M��^crϥ�滶��2ngq��P�Y���@=YL^wy��e����X��e�e�^��2B)� M����դ�Z-�`�I�e��X�sݓ�z�w��-��8d.?�Z-ßo8�B��Z���5��iR�h��x/�i}����D��p��V=�fH��O����^�.`��'�ϗ�O��$F��Ok�Uc0��Js���RKbyF�oO�����J-��=CqCǳ�<�P��G���5t@Oko�4�p�dh�0��g�d�R|���P��ȃ���k.��>ח-B�Ѩ��Ǵ���u+����q�@'/����3*y�)�vxm���� �w��ǀ�>��x��^���U���S��O1��Vf(s���$���jJ&�w�kiT
���D�c�W����x$y;�1��d;+������e����2��?���O�f���6� �6\f�=L���<<]�^�K��p�&�z�-G�Y���f��.��7�}~9p�g4����Mg\sC�����������qFE\(����An|�n�?PK   �X�Xmb?�4 �R /   images/9399b738-9a99-483d-8480-139b77408719.png��y8��?>c0!�l�d�%K�G�B�5{vB���L�ZB
�d�:H"K���
٦�پ7������?����s?�9�>�u^����]uFzz�P5�@hF �C��J����������	>���a5�| �g#Cp�N�*���:�������/����co�u��vJ^�����`T/�̍�?��}��k�D<����Ws�P����ɂ�[�F���3&أ�P_�#��W�<fsc�]����W�у��;��ܒ��~j���P���X��b�R+fl佄��Tp�Z�I�J6��_c�]�#����F�ͱ7�vS����x�������89�K?M����Z�]`�C�+���������Rf=��V��Q�=�i�ȝ�G�ɰ�Nw55��$>{�Ֆ~0=9@=´�풬>�!�����e��U�c�!�D��ջ�?)�ԫ��|m��2!ڧ�t����
��G���}˫9�h5\���L��9;��C5w�q,��`��M1DK���E��(�?AF�v������R/����M$y������s�ZD֏�J��P�)��m=��φe��Iꄔ�f�,�8����'�T��O�.�ܹvIQt�V�6"��L�^�>��#�As�c��\dU��K�,&0%*љ��m��>k&�+w�d��7�l���?.�K����{C�*�"^�A�ѩ�P��]�g,r,�!j�֏���!��!`���z��>��`.ǉX�0-�L,&������z	��]
M��H��IQZ��9-&d�i񹻟_�[���߶4����-7a1�� ��GGڸ����
���U��Ԅ$�Qzz
$=��)�-�����E�n��h�S	��{t,�4c����=�%u� ���w�9~�V]{嵀_���S���G�1�2��<���;M@a����=X`>�'Z�����?��?W�l|~$Rɇ��������"��QC�ŷ���H+��D�%yy�F�`[s\��(cջ��5�����T��U=�R���[�<fpJ�y���1JJ[]�)��|>ؖ�J��`4������hU|C��an��]�ӔӶ.��UE�l�k���
x�왞��;RM�H�r<���̌2��,ȑu#���Q�����0�8Tb<��U>;=��(����p��5\ǡ�p��v�����u:�q()�'��*U�"��H2������c��6V��I��;Ae�bJow��Sp:]z�X�#�}R�t�9M����>g�!~������r[�9�6��#��iC��g_��(�����H��D�F���Yd+a5I0*�x��V5H���I<��SA�/&e�V+U�5�õ=CŠb��N!:�G�Z�0T΅=�~l��}��[o?S���R�\��ʌ⺕q��ບdҷ�G^�'��G��2TPR&����k�U�$?�"����Q�~+r��Ay�׹^�S����8�',:E�Y�ʪDV����ѻw�c��;E)� �lZ�Κ1#3&��Ҥ)�d���3}���L��2�4H�g�'��"��gf6�qa��p�X���"˪�lj��)UbxHg��ʴ���	��8�$O�PJa�J�϶����/�x�
���#�I������I�N����W�(�i�D(遝9MaK�x�Pt�u5�P=(�������BR�)5�N��x�Zբ��&��]� � )�5���x�EM������@C�i��U��1�_i���#����[د�A��kv�I�PvAAA��%G�ޏl����|��N�e����<D0�����%W �s�Gb6;j�rnp�.���eΝ�-�����+mv�$��!��Z(L�7�0��`|;L4#��OC.���l�>�m�T��0�vgZPU�����x'�{tt[��ۉ��<6��<j�� F��2k����|��k����38xS��2�G���(((�D!r*^`���� +��Z��?�_wo�/k�S�v�$~{�����
��H�k^��K2{6��!>h��� Z^>�L6�t��;̏)z����f'�q/lE��}9�(�<�a��u�C���=��`�M^oj()��fo�n*�^�M�����6+�FR�b��'�-�}B���_��v�I$^0��ܣ�(�G���R��z0�^���{�(���|��ɉQ�ᮼ�P��Q��"�@%��0��g�����\�G���{ةc'f5I�|��:��q��7��.�����a���Գ��:�>�������2��x�U����'�<��+y�z�Y�DIK�?&慴�$N��+NC׷��x�̘T����-A.��8Cw���V�|hծ>_?���يLH��ϟ�S茹�����HJ�#�`����,W,�`���)OO^ӻ��0z>�:�6�X����_}=�dLOg�[�|�M	nM9K�>��m��E��Y��r����˶�,lwGɥ P5�뭈�:H$rs�%u�ϗ�����h�w�������>��Rd���R��uIk��Ԙ�˞��kq������;��iQ�/��sz]J�ȷz%%�%���L}�����U�(�w�wK��w��u��q��"a�/ިS9���~9�@)�;t�^}q7�n&�o��<��<��ۄ�r���E��̿�Pd�3]�g�A�a�G�q����a����"*����XLOO<��zrY@�;�o��`'�1�4Ei��QuSp��k<Z�;��M���$�W����њx�K��s�;���EPo�7>8����O�'�Y]4���W�sB��:���2���`��S5+���b?M�����y�"�
�Q������hC5w|��v�U�,�#�R^t����2Y,O�@-�3򔱾�Ӕ0�Lp�t�Q�"�L|��=eA�䊕O픸.X��)���cZ0�e|<D1��KD���u���Oc���tg�43�Ә��8)Y����Zχ`�~�U=�i�Ku���D��D�G{�Pu���TM���H�^7��\�G��!�������tt����7��P�`�^Y�&��;G��n�M������v<\x���A/�(�Ǥ\�?__$7R��sQ�h�|�çC�	��,ǂ>!�C����mN���5��^��q�@�tz<H�K5��?�e���Ia�2׳��Ԥ��EEN�S���uwNtUK,wq�|������9y��6pn���-�daK�Ł+m�pU@�����	�$d�]���`b�2�e��Td��G�����dzz�~�Êԗ�&����k�ܣQ���Aҧ��	�DTG��@����+K}�9rD���83~�W��=f���ɜ�|Ԍ����n���^�O�X�������`��g�lc��	��[Q�yC�W<����PtX�I�I���C�r�Y~�J!;����ͽ����z�V�\�K\����Kv=Os�q|�W$��s<�����H-�Zb�f��()+;����%�84@��y\/�Πӿ��[��T���
ߒ��d�NFb��,�9�a6e���@���w�1��Eߥ�Y���^���-Ey��"�-j�n��=
�8?����֏u2����iGDǶ��1����JD)~l0Z�-�`��t5 �e<�T�%*2������-�6��z���}��U\��pZa^��5(ذ�Æ(��b���������˦è����J�a�mQ�J����M����b�@^�?z����eh�g���VZ?@`�"8�J �|-�:�3��jqQW�ť|kNa�Z�Qc�t;�lo�q�G�׃��y�r.���*Φ�!/D��-ίh��/�y����66P4{�_�T6|�R�I&�FL�7��xq��/���k2#?ݷ�	��B���`���b(���SV �=1H���_�� �&�a�ג�*��+{dYNk��^9ʙ��0���R<ÏI��s�1K��9}��;@��`E�T,�YEǏ_�{��)�^�m�vbV�Ac��o'�q,�g���5{A�k0��,Z���K]Sc��
�~�����MD�j�Ȓ��3y��<�z�����[V~_��s���̵S2�i3� ��e�P�E�O9�g�9��"7�97���:�C �g�^b=8��a�ܖ�&>�>���Px�΄�z΄G���g��{w��b�ǫ;��c,�W�9��U���)�f�8G+a���E+sw��{��jnaa���Kn47 �Ch9���\q}]�R��K|C����]���_�$X'��7X�ș�^/���U�B�sЛX�T�{�m]�uZj��3�[^#�.� Zjأ%.�tRC�Q�[U��2���KB�JKK9�ϧ��7'�ܯ����zn$Z	p������z��
��O0KʖQ�a��+ZG�LQwM�ie1/�XW4���O�����\cYo�����7�?Dan�\�C? }�)�)1�=\Y�,���[n�j�d���W�屓A�������\]+O�34~\Úr��$>��}�o���C�����8� �gc
*�lս!:`�0sk�]~qYz򨦕H���<�
�9���Hm�J3��c ���FB�������1(����*��X�E@ǐ���+����(gl�Kr���ĩ�Z�S�A���f�V�G�3G%4<ҿ��=�r!�pQ��6��	^ɷ��	�ڋ��S�O��za�L�����p�;U<ߪ��Xt[�z��PC]slT�<�5���n���.X�����,�(Y���������WK�g�285?�ٓ�'�	<�J�9��Ї�J|,�3��"��S6E�"wݞ��4?At�K_��<���<�(֯��*�o���#l@�3��g3��=�����w%Zl��(T�(�}�]�Õ���Q�AR���~�55V3���{������%�9Fy�;��Ɔ�\��8�J���Y�[�ʈ�7�"QΜ��x�=�J�����+BAK�.e�Pz�"s�'���4K|%p�P6���'ߣ+2�VLÔvYe��~H�忦L�*+y��`�S�{�88�?>-��}W<1���� �Ge)-V"��k�gh�A_���*B3q�C5�������Ѭ�v+~ fwe����y�br�E�m�+Tr+r_�>^.R������xӳ%��F#���)�B_"&x4��jQ��{Q�����l

��_h/)D4�<h�+`|�#���BE�m��^��Xo��b5�gB'�>���zbW�<���c(��/?��$�����On�;��Ѳ����U�( �	���TY�!�4��oR��Z�}q�_#iڣ�����V�``�+zF\�LT6��Ly��D�8V�ս����m�^�>�[�6y#��io����N�?76,E�)�SU=�Lf$��.T�������k�y��e�������@�� li]3i�h�WC��m��߃I��+�����ؔJ11��>�`��LF������x��%n�E�в��u�:1���5��YB~����H��)L��@��3#OF�{Hjg�|�~�=H�}"y�����j��jw���W2&r�S�{K���ʊH"'�L��0���%��-���-�
�.�a��V��cc5'+���
��F���wOG���1r1�Ɲ��[�^/V�{�#Q1=d)�6�ͫ˥("XX&�����n�$�Wy�?��9����%RO�P�߈�z�N2��8�<���+?{;O$.�߭�mʹ����k��F����k_?<�|��zw ii��`�Sյ���3T���Q}�7:L�\X�EY+8��h�hʂW ��g `�Ҕ�>fu���T;u���ɼ������;��n�D&��7?��"Gbx�I޹�U��گVu�oݺ��rF�j'3��$��rg����q��p��t�V�[D�d�/3�݋\p�UcA���k������s��~&��QgmjR$}�W5��g�.@���������Xh�0� ��1'D2��~uuNY	A*����[^©y/���C,�hg���fy�|<}1rS���Ƃ}Rat���Q����0���>�r5�.�RY��f�g�Of�$�Ő�-�ٺ4ɁE�RL�L�尦�Z���*ۥB��*Wgg���f�\�C�A�oXX��g]M�X�"�ɊEێ��SΖ(L}�S����8M�r����n6kB�
��1D�L�r��sX�7����`�2೨�9UTy��'�Ϲ��WzY�LѵF��y��⩠LK�j��K�P
3 ����l�rn�� �m����&�T�h���͙M܉�F.�X�A�v�C�x��#�59)j����-�pyDݜz&��bcÓg����4%������p+��?����9~���W�-��;���&��kk��j|o�(f��ئ �U�����U�`��;n���#	�ۯ�&m�|٩�u"D*�4�gH�^t��Z�~��eJHjw@/�\�����e=puww8}1X��g�yI�|#���b˻��6xC��9�,�(�F��ޚ�����AeU�G�� ���oM�����t����짖D��bgC\��2d	�2�����j�E*��:����"��=��@���3��<�ʘ��jn�ʉ���9�:{P�҈B�<�/�-��VC��"FX�yy�U�����4���(ᅌ��'n0z��K&�A�{�wwu�#��H	���Dt��-��n)�<Ő8	2��c�b�]�B4"Έ��a�}�Afg���369�{IΤ����pۮ,�\�dtq)�g�8e�q�@��=.�c3 7,S�#H���w,P�><dyzΞx�Sp����)I�����a�����~�i�S�������_�p�O&�Q�SWm��4*K��K�<i�qF�����À�L�,�ݒ�mIR���}���% �F�0��8��X�a�Y����N�g�W������wЄ~�&�M�y�a�B��cI��"<�#D���[Uơ "㠍�_Y:*�\K����P�s�K�t�ȅ���=�9��uh�i� s#ER�d��	�3��p��{t�O��o�?�,󼸸2�8���G&#$-��'�Z����#�T�W�fu��}��I�c���Y�nB��b�dy� �P���5�oݸ�;���o�|-1?��AxL�֏�:�ǉf�f��?�s���f�ٷkT�cD����V��ד�}�^��M�(���*�FL�~h���h)���J�]����X�=|�rF�����p����ӳ���L=�|��S�bx��w �t[�����0�())9��U��n�����vcLwB]��?����^|�28�����+`Կ���󦗷HEo��R�Ԫ9�E cO!G�.B�=����R���������r(.%����πm��b{���B���JU��0ʺ-5='M~���Ē�dS��Ǎ��Y�$����>X����r�aK�.4,��V�~��`���<7s<�(qq���0\�Ɏ�����_�T�qt0|݈_3�hɁ�]I�F���<�3E��c��c�]�G^TWo?�#5�R���t�>�bB�$�|;pT���ւ�
a��Ӱ^}�d`{t�չ��dQ�h7jQ*E�kF}|��K�4i����b��7	� T��p���BL�̲��k��6�g���Xʮ/�Q��;�����*����Nд��Ǎ]*���\v�ں�ԱGI�,o3Ce��G���tf���@��`"�u�f�]����,�fe.;i�=�{��ה+ug�)�i�aJ>�j��r�,�6���"��p��jt���g�Ko�B��*jU�7�K�U��<e��EN_�i �j�-��p�����������\_+�H�}'1�R�gy����)����|��[9��ɏL��a��ߙ��g)2d�x)��ߋy�H
���d���Ǥ�~�?	M�ٯ���X�+M	"�����(�E %���to�5J����C��b0&nKp��{`����\	�w-$�/H��3�%�*�A؈�;�_Y�>ѝI!�l.h��1�B���%�Z7��� ���ĩs7kY�ff?{�ȳS9PZZ����;��+}�\�F��A�5H�a�NYl��[%�Z��<�)d�!�����eT��Qu�:��)����V��`<�g�ġ��sE�|�8���h�O��Kڢ�d*0�V��|���)���뻡�R�گ����:��Y[*-�n��4�m��9<���L��B�	�?z�~�r�G��PVII�O���w�ha����������#Q�,��:���"�~�w�QX%�JtD�ǲ��3c~�ʬ�.&����D����h�%(�,�xs���/I���Y({�}�_����j��g8VaSidW�]x�p�O��ag�?p�+3ρ4%�����/Gwk�W�c>��VAՈ��
;Bv��BƇY���<��}R��0�>�ڄq)������^eKΌ�vp�ш�\�B�W���N��_���K��I	,�^/Z��P��d1����q�#�
�ģ��5:_ʜ�j^��V_J�����g$�6Aj�<:��b�AΜV��H��g*�^Y/����4%�w3��-�,�vst�c���W�����W�.#��;^�O{R)�F��PT�<�e�
Qz��wak��4��*i�ܮk$��JR`v�&���Ф!������ښ&�'~P%�&�>���9/��Lno%�o	�?H	"y��Fʚ>�d'1l�X�� �F�R��hU�)�B�*��ÏV=�h��u�R��1��#!��±r��HD����.���'��9Q:9\i�Wa��y�t�������h�"�ЃG9�fC�h�������BX]1ho6
����m�pa\���4�ns�CEYsR��R���S�2�3��u�؃%I?�c��Z��ӆ��L��{�f��ᕗ0�r�ˌ�T �����@͗4��v869�g����=��S�r�����L�\p�%.K����XM\���T-�8���#F'	<� �P�������-�'�#�e�QP�=D�P�����G����eǶ33�r�9`�.'�ʶ��k�$~Y���x1hG�?uYm�PEV��u��6ٸ��߳-8Q>��/L.>%�3��:љS�-��X�_8�3,7������q�tk�:N{]�ߙ��O[\aF�F�4u4�3���$�&�Ro��!i����q�!�����"�)���qܧ^׳�Ū�by�9(R�������r+�szp`�%�Ku�&G�U	�3���c�0��҄��@7��Y���:���oD����G˩�A!Fԧ�I��G�=�:���[X8I���6�X���)��t�����0v�J�}o_��h˷���ߞ7/!�`|��L��|(�f8!z:�Y����0�/�s�aǀ�ak7�(��Ud����ϐB�CNCy£��sR�)�q�ɦ)>p[/����0.�?]-jI����/S��	���<���E�I̶'�x/5ѧ�<W:�n��=�j�p�4)R,�e	L�.��S��N�M�b+^�L�����{Qp<CU��=�J�[�-��k���E�-��~�C�ݾ�ň��l��I���&�sLU��pcr��QJzO��%�%|DC��n������դ]�ﻞ|�Jt?�4M��Q�/��*�dJ�0:�_w�E/����UHi���gC�=����6?XZ�J�r��d-�h�#���z��z���P��J�\�:��0��a�����&T��ݽN&�����dB憾e��T�w�$,�6��"��R��/�fJ	ӑ�����.���ni���ґ��c[^�?v���� @�X���y�_�xF!�%�ëb$�ΣTE����蘆Of-�������Ѥ�K�����Hm-�ބ���+te� ��K�B��J�LC�/=;\ ch�Z_���)�_"���e]����7�6�G�F̭f����:�63_8�Q�5Kww'He��8�����B���v���ƓB iН(�ŵ5b~�i
�2�o�o}H�*qtF�O���*�X�����=�sk�Y�+S*Su�W|�K9n�b���:eA_�tU�t����B�.�jd�'@=k5�x�!H0� g� ŵeMǇ�r�(��I?%���6��K���ޑ�R�L�p�����j6\*&����c�5/^RuDE����#Lui"ۜ�/��I�ͥ-*n�\@�$��B�Nrj?���Ƕ%�hH���T1��O�p�{�lM��5�W��Y`�{�����b�TJi��M�J�%[ί�4�lCV�1�o�)k!l�!/���s̆4/�d��*�s�Ke�<V�Ǯ���q8JvwȋD�w��\�R������?���-
����@��MAB�l�Es�)`��0Q�A[��_�tJ7ve����k!;4��i�w��8�1Y���j����	z�&ؐ0�9^iv-<�4Y,����4Hx%F������I
��n��E���.N5uO��׍{��,6aA	1=�e�-��]����`?G����XE�"�{~�!�.x�R�ҥ�rs)Ļ����xD8q�����!�<�J�!?��l�aJD����r�V�j-��H�׎�x�IDF��4�zL���Q��}ݹv�9���ߋ{�2:K<��y��	y:��~���x/�A�t�]�������R�K�J�%��r�b �O�ݝ��,R1� �W�Gg����aiQ���������v>�w?W)���2 �H��mqUst�Ч���\3a�pYj�u�:N���kvT��G�%�b�ض�nv����6��P�&Y�,N~4K�i�����9p���xB��P��(��cj�	�s����<�i�1uW��N�9��� �}a��~[�MzK
��7�V�ч���Gp� ��4�0�{K�f�ٙ���˶�H�*���²Nq�����2>�?|w�����Uzޘ���f��o[F�Q� ���AѼc�߆C�M�DG��P�&���ǥЛTz�Ì�6�3a�n�e�63T��@�ã��"1���Z5拊���y�#%���fC&���y��������kZ�y�P� IeZVe��Lx4&`�,Wbz�W�9�d���/-e�o�,ֱ���E�����6���E��<�����G^��	�}����K��O�(��1ckS��>v'P�� �9?ʜ��5�kʦ�|s�od���:Tzu\���(����7vȘ����/.mɍ� ������i�yf8wm���#�U�ĺN���jG}� ��C���^�3k�7�n���
ho�/kr����󢍁���;9߸J]`k��0`�M�AMg�~y�����Ǻ�d|�ò0�h���RBؼHj��>A��O�����)�^/��
.��I,����F���؝|��LxM����4!6�I���S4��#��|���|`O˭;Md�(�c�r=����2��>ɂ@�p�7Cz�$6���R��RS�Cˍ#���\^$����uŪHQ�1t��T�vd�l!Ƒ4���[�Gd�З}(m-D� �wu	�-�]8�eGvjs(+)��O*ꕎ���r���2���|���V�zQ+�����e�Z��q,x���6�7I0 ��]s)�kUtZOs�cǡ�p�PK��a�W����!��v�*�hp�,m�ƒ���B����^;{CAYk*��4g�~�f��U|#�����h��SmסJeEv�5>q��yr����*G�a���!?2QV�I��{%nb��[<�=<����������u��y ������MqVd�bD+�FV}jJ��z8�gw@���I;)J����Wo��`:��H���$�����%a�3�䢿^�$瑒���8��6��j�*l�z��W|���@�������:\���$�yT���,adG�~���[�.$$�	rHuk}w
U��,�#F�ܥ ��~'���_�4�r���Ґ����3 hY~��ߦ�H9�B�v4�R����V�l��&��8(�M�1�+ga1��N�)SM��={�G�r%n�>ɏ;����9>�g���P��-��q��������S��N�A��zd0R-��K�
��w)Ƒ?[��	��A�v?���74�
o�З�O��s���ƧhvhD�ؐ�b@���۷^5P
�G� U'�P�p���1���|ݼ��&BR&��-И��#Xq"�G*�!�r�-NBr_�E�x��5N93�&9b���XU�#?���E�t%`��-�Y�Z�Vؚ��tXJ�9��{?�:ɛN�+�DR`l���U�4R�B�\ �5��/�q%נ��=�|�P�hp�y��퇜w�EX������x��O��T(�%[+�<D\YؖC+�#8e�}e������O�/v>D��wB[����r��߯2q?�m�s�)�&>/���4cF�_���י�5fK�@�����T�#I���r�������m��%zX� lF���s �Q�}�6�ސM)tE�x� ����ΣB�������i۝��|ᕑ>BP��a5�WG�/��p=qU�b#ɋN�k��[9�`9Z0���~7�U����{8N��wp����u˸��0�Aƪ�HFc� ������{���q��	[�Я�M�i���oQ�c7���=����۽!	E����y�K���V�[m?�Qb�u�����L�:r�o
��3i�bU� ����=�L�r͐�8��9^n�K�DV��W#�k�2Q B�:q2Z^�2�$�V�?��b�iV+�߽���A^��z��
߽=:O0�sj��{}v�0�ĵ��Fg����S� ?�:��_�G���E2��!s��������~#�t���{� ����G�=�r�My{�<孑�S&��G��`7��<p��}'�G�q�B�y`�9�������1���� !ǩ=Ǿ��X�� !��E>��M���\ab�9洏�!�qWY?Z"`�� b
�ņ���p��7Hq��
}"���� ��lU�^�هũ�_mp��vl�a�?@Z�R�F[�
(@��� {r� 7�X�v����Õ�����{ޞ���4��b }�>�;D�Y`y��r���!v��}{���]��C��:�|#A��Թ���/;�M�C�����^4
�^��+���e�=i)1��s�������!|4���@YJ�q����z���?��:x-w�����*m`,������QNE"�-Ͽ1�ݻ&�-,��x���'�N���7��@�>�+Mz����t�k3� 09rʃ0hE4�4(O����n�C��2����f�6�|u`�ǀ-7����{��O�c5	i�#���w����|ds�ӥ���cA� �b-�m�:	(	j�;�s
��Qr�S�9��-�w������V� �˝�����N!d<���3!��;0�Ņܥ��}��k�!��7X#�r|he�P����.����+O���<\�d6eSܽKUl7�]��T������ҹDp^�\";��zS�o�@/.�A�"�_�[T��ao
��?���G��Aq�ܼP�Ȋ�!�'��GR���i���wg ���	��@�p��2THp!��kD��-Q�,Z�{I�Bl�p��^���8�9<���u�M���|<�`�P�銀"��&p�������!a�Uzn}�����I�U�#O��e3x�ݿ�ˌ�D_c����b��V�~���"���M�/s}�����"ӡ;��>�'m���K����>� ����ۤ� ab���G���O�O�!�S��ʢ�� �Lf0�s����c��7E��`�=V�߳Tj�᭼���xO�~�Ջ������ܿ���<���{�'F>��Ғ� m�qa����{�������')����t���GtS�;����"�Aŭ��֗�mn��Y�n�~�La��g��������y��w��>�X���,@����D_���kX���3��Ϳ����L��*�O��J�b%�#R�RdNo'�P6��yl��	z(;�9P%Ϭ��A���l��.�_��\����9b~�W���ρ���nkv���L_��1�+	��Hl�v�G؎qք;ߑ���c6�;�y�o��t\h}�{���Ώ1�1�맫|~X:������������(G���pFS�����V�>I��S������s)!�.[e�F�e���Dǰ��be����օO�Dv-!w�!F%��ڿ�۠?�$����ҲP�A5�6�0M�/�4��}�j�a�	ݿ�q�p�z"&	�Lv�������Y��'��K#Q��'�Sf���L�ƈi�	�9	͍�zAO��'�0��h�ج�e�q���K)Y���h�?G�<�!ܑu8���o�Ԉ�"�!��c��н{�1��.!$[�n"������k#宐�m��X�cL�9����='��)���K(����7�������Z��R�q�ŗ�3���+A�wEe�_�E�M��/F&DE���{zpG������,��Χ��+н�ٍ_�ʲm0ۺx����DR�D�#�L�G���o����V�j�V+�R�Q���k�%��S3��FF'BZ&6�R��x�$�`��-���q��w�M����9�5�7;��ʈ��'&����@�������T��}Ϡv��o���9w�ڣ�>]F�6��&fG���0u-5�?=0ka�l!����ǊM^�X)cb3��v�TcC��(��"?#�6˅�z��G��Y/Z�ې��(��b�AOϯ�vF��H�r~\�y��;��K���o(�Y�ޝT�/o�N�>Y~����~�!�U�InK¶ə W	d���.�I^%�U�<*�6c6��F�b����>�R d,(F���Ug���(���-eg���i�zRԤ�4�X}����zq����1�2˘h���o7HMZ�+ ʯc��r�b�D��۱Y�P�I���C�g$0"m��A0�^=�Z�G�-gd�\�,GYvYk�V-*�Y,�ܼ&|��^�fX#1Px�]��tN\�
�\��{�*s���4��,5!0���⊻^Y���B+4��9<O-^YT���7S���0��,1Ẹ���@��{�w^������WB��<��"	��؈�'Z���s�y��{tՂ6�?zH\�}�� �&ddԝ�6�ya2+���{m�g�����j����A9n��[!�Fۓ-�������^����+�j�����+�l
�n;�-Z�-�j|�˽e�tH+\*��H��o"��F��s%�����v��F�ϏZ��ƅ����#�i6���w���u3�8���		�'�3����!x���;��V��nw����:x�F˸|&��Z�.�b�%�ꢖ��'6S�F�S1��w�d�W1&�b2�	�߼4�fkUP��w�v�BV���Dj��:�S._{�,\(�uD��ϐ������,�R�V��\���Ɯ9�z���`��ZA!A���ݍZ�[�� �/s����%(�3���&Dq\�@�@����aO���~$Q�.��|_�����J9��G[(�?Ě�ԩKvvv����S*�'�@����h�����
�d���j`Rz�L��g�}�$Ig����_��ԗ��u�?ߕ飮��Z���X���@�#&�hj����e2�1ۗ�s��v�OH2FP�\����K���F9��^6�����Oq��G]��W8�t��i��Wv��������y��]}{��Jn��ٛ7%3�%E·���A	�w����c@T{s��|~h�uؗK�	,Qش}�
!3.O?�؂;��us{M�ກ��@�{+|]�\�Z�}p#f��}��\@Z2��!��-��z$�\�y�5=3���K�3�& ��+��::M�#d����7(�"ͯ�hy��d�%ςw��,W6���х1��QEd,<ĉJ<j���O���sVy��#�X��
���31� a؈���nX/kIγ����%�В �W9Z�4�1�Y��ǵ�:�.�))���;l���Q�驺��S��ɏB}��(@efd�6��f��������~}�=$����/�_?M`G(O(�N�$FĢt��<I�?S�����z�ь �b5��ݣ^{@5�����5�jjj����z%��z�@�C������t�^������琸��M��1%.�3]/�|=�F{�-d"X�?��?2�c��혞��w��_���P��s�Oտ[������'���Y×�H61��^D"qy�vw�*~�`�������L�rq�W����=\�.��٣l/�£�KݴI�������2\���U�ݭ�G�t��;����Z��G+�,>Ҿ����B#�{�����^ǳ�цC�#��� ���f���S�$+��%�t��;w���͇XcL��@�����/��۲�M���q��ccc��ل�ݷ޼�^r�9V]Y`��k�M��r��lb&����昇B�E��J9y8��Oa��L���߯�Dsm*P1��*󛻐�ڪ��D�/�b>?\���&l��ƮA�o�jY�7пQi��8��� ����vd �����O��t�
���Y�
F�^���2�Є����5�Ł+."V=|KЛ'��Wx����<s�^؏��]�
�;;�ܜ�2�"�����/�G�;�]��~�=���]�f�Jo&/�����C��Q�p�X�2U�.9��0bR�k~�tO�S�a�����Ɓ�.z{�x����E�����T@��������r�s�W�ۚ��<��3W>�W���\��-O>��n_��|L��k3�QPw�ӎ��HR^�����!S������'ܤs�#88~������G����4.�V��QZ��5x��0��q����?�:~��[��ݔ���i�n����/u���B����\X�'���!��i+�_��W�X��P!)��d�������ߴ�΅�d�v���KgP���3i�I�u���[�u���+��G���vyz�B�B�はC11�Ɵ��n���x�'��L�9hB-�?�u�%%G�ex��<��:Up`�"G������;��2���ʶ����"���AC�kQ앁��%�����ޏ�+���C��g�^a9�+Y�v�$��4�$�6�Y����Yƛ�o��+CK�k��������� eVRFHBn�ݲB����eoR���.{����mo�����>O��������t;�3���8�y^�6WXz$*eD�q����|��3���5��Zz�3�ٚa#���b�)���7��7`��Ҧ����<' E>b��1<R�O��Y�FLɿ'�yÝL�2���\��80�2<���\�ם�!��ɬ�=`\����Ԟ�������<��}��a�*1�0ə�V�J���7I��a2-�j��3�ƾ�A(h5��ey��Y���Z�ar�T?�٠����#{?a���;i�[��㍗'́}/+h�����+��f1�%7��%�pz�w�>�:��珑vc�p����5I�8����u��F��e��<��d�f���f�c���	p9���{.|��QN�u�ŝ��y�R���\��{I����j�2���]J#��������q�\h�bM�-��A�p
���/�Y]��"����2�{��5��z�C��~���<�cp�Z['ZR���v�^����j�)gTH(��1�ڢ�8xӠ'��M(�5�:��.)��ׂ$�4��A��ך$�r���#�:EI�z����A�ׁA��1��q��>$�5�B߄��<���Y�����(�����2y�]}9ݕ��?�KV���e���	��R�\`@�c�Cw�~��E��p:Q�\�����,��*Y%;$�	�b]�$�5*��S�б�E_�����b;G�����v˃kL0�,J��ل��&-Qο�+rss#��2����6b,�0 kN d`a��"'�f���F�LϽ��󳯭ZwDDR��u�����GU-��FR
}�+9:�@?��ChqH�1����x�֮V/$z�>7��JR�35K����r�N�N^�_ܬ��X�Ǐc�1�ջ++*��Ww'"�53�ej���]��8y�$Q�SИs�0�f	c.)E)c�3S�;S�Ӈz����EV�����Oݻw^��h�D3���*�k4_��>?���(ȌИY)=�ʄ�t��<��Є^{�a��y�n�����ţ��-Z�'s�]�lkЌЇ�a{[EE��1����ij�� ��e����;+G*�(�n��P���5Ec|��Qi�R���ٰ�Y9�n���`�
ˋ��T�1�dz�,$&٩S?��u�XlNgwY�X�t�b|�~F'��$���D��������f�yX�[�j��f+��z���t��Ġ��&;5��=ﳏ0�[M���p'���df�l�A����0�Ř7����t���}��7�E��gM��w����p<��Ϻi9��i�PS��w�G&Z�f��륬H0~�yej�C��C�6@�[*n��'tOtuu���u���:K��x��B�	-�S�6Z�����ͷ��VB�߿�v cUm�<��=�f�W��$��z�V�!$���P�y�bAC Ƒ�`����h������P��o��՝]ŉ5��n���Q�Ŋ�_�(�3�`���5(3�5��Z��l������ӋWL���ԙpE�t�"�o�qW\�&�ǟ���?����RJ�<���9�;q�i�.��t�]��l;���$�E8L;5�?���Uyh�ȓk�z��W��?Z1��8n��%���x��?N-����
g���S�,%+��D������0M����r���' �P4��3�D���I�=+��$u{s5�g ���X��P���+V,r)_M��X��(�7��	 �؄C��Z�3����TW��0>Jk+=���Z[��l�Sw5w�������\S�r(��[�1��n���EN>�&�tJs���s.�j��Zy�[�O��ސ�﬏��;���,�l�����ĎXfq�HA"��Q��J�'���S�o�J�L�H�5�����?�Ett49y�����-�t#x-�;w���pq�A�ܹ\�xP���~�x�C�造X�-�|T�t},P��c�&���+򠬮�k���^�m@����:��g�TTG�fXʊ�A��0�J��檃�A{������o���}گfk[����&���@n0k�]M���j�������\�]g�]IX���ZM�ۦ�Q�}4nz��=;2�2N�ߛ����~�<�a8ݙ�=J:�6�Ά�  i���A�M���Y���;��uV	�Z��xfV����h~�a~�B��d�I�jC�,����~��
wpfmIr"������bc'��:���g�v��Y�B�:?b�f8�yvlo�G���9��X��o�N��JZ�:LB�'-d����d&",�k%�Ѥ��y�=��(o��9�o�נ�.�?Ĝ
��M����Z�Q"�ׯ_z2-��%�șd��.�߬�Z�����te���lK�r�7��{G/2��$('*�J�b��TMć�ph"O��|ARij��ի���dk�@F����G���+h�������1��"��$�k W�M������m=� :�f����Ս�o�x� �9�ի�YUs[ϴ������z���k��w"K[�M�@��AWM�.H��,;���g�RL,��;}�6M����?\����� �xG1c���/~�@�Y#����;)O���'U ��5íQ���µ-ޖ9��\��t�%����|̽���J#O��}� �\�D�'����F]�555�%��nߖAv�K��9G�};�iɧ˒������m���}�U�j0��3���r�x��:��	d�������!!![#Rlǎ��)�|��M��å�5K0�n/�zN~�uV�C�~G���m���\IyT项y��t[��V�'i�߅�7\v�� �"�9���~�V��\p|>���iJAǂ��Oj��\���"��3 51�w�հ��bk�L1����yKS]=�;�0ad�q[�Fϓ~�44iIr	Kx�EK�j���ې��ٔ����ݭ'�cD�R	r�=�7�p�N����p=Y2�Z�����eč{�P����ٜS��e�}C`m����:B�,���D����u߀[��wS�7��;��O/�������$�/O&Y�[�-@��=�u떹Uo�d؈%�i���_{{c�~&����_���whO�3fp�5�1O��T^}�4�����% H!��׸��5]�O�W���{����Q�2d��ߋC�RR�=y��O�`�E
�~�sssw`�W�l�f�La�\n�0�����NFFڜ��WŸ;G��2/*����ց�t�|+�UW����c���[5~"bbbE���
-��ܷ�.���)��>>��ւg���G�S�M!]]�^�G��!��"�|�A}&Jzzz>؝%�4��Hw���w�5>� Y1����Ot�nL��Z���ne���O�azg�m��t�'���۵�����
���k���dw"ƤPN+�M�Vl�Z`��)#f7����޹S`%��%���=�"�="���3y��xzB��p�u���\�9?ۍ�-vM�1U^SS��EVS��a=3��Ȕp�|OT��j4ν�I�OJ��NC�p����W�3�Ϫ9Oa�	?mM|�h���F��<^[_ U���0�S@����|��VYU��x�م�Y�����/O�&�	��wă�O�>M~�64|��X�#]�B}���*l�2�(�C�E��!ܴ;�i`Ѿ�����y�aI))$	��办��<6}V��+aA�u�M� �e�M�n8��r�x�cԕ��q:�Um�-e� �߀0;m�4���o�J���6�8���,'��a���>�����H�$Eu��c��o  �����|N>� �I����T��o߾���>�<d5�)C粕)��;R����c==���0N9x���$:�=U%�nm@3 e����ζ�@c8��%��@�(�z�gM�e�Ç�o��W* 	q�����Z$���#�uh���k�DT��~O�-��F��7������dl�oJhw�W<�m����g�;�o��TB�i�Dw�tU���m[lb}�}^�;��
ɍQB잕<+?��eȬ ޒY&���PC���@$�>P؛�o��4��T��-.�Z4��(m�[дzW����Q��~���3���K
�(���R����H9X������ԫ�d�^+�*�3j+u���d�$������G���J��6�0�?�rW�+�����v��+n�~u�����J,<��������i�a�=J�e"|6�ek�N�0!�M*w��V8�ǴgG��ٺ�<��m�K�ӧO]Yq���i��K6��}������q����M�i{�ic�]�^������bRC|�O=$�;Z_���$�~�t��h�f��U@q�t��l�4�u+������ ��d@�Fh�dx��\:�|�J��,�� &���_������6��f�,��9h���sr��/�aADd��O\X��bbb
z� *�?x����w 2q=�8�(S�ů�9��t�{����(L������/wvV�Y���,��f�R����ٵ��]6pQ�#�'%��(gF�!g	J����^
.ߺ�E��+�^̳���:֮0�ٻ9� )I%��hp�㳥��4|�@+L`�G3��n8mXr=�1H�V���#��[Jʛfw�v�����|}E>�H%x�*_��e}^����W���%8s�z��dZ[R�����AOA�����t�ۙ��l�� 3��_P�hw�+M���~}�	,�"(���I6 x��_H�?����;W��*�1K����e<�e,[��T{�2>!*��$�r�+���3�|�6Y1-���S����J��Bp���ͳL���`'�8��yl|��eAAMN���)hcO�ȭ\�.(Y&�Cwx�(װ#�b�$A ���>/�/���P��Tj�a�~���D+�&��B;���]Y���å�Db���@�}�����SS�D��B�!�tд>i����İ�P;h�%�'�,��|F���C$ԉ �Дv����k[�;3u0�l�ǛX89�N�<���ِ뺐��\���s��UӪ ��*
J>�T�yܳ��A�K	�`*��!u��)޽{g ����0o�T�5��u�>5X�����A.	2L���W!����j��7lf�Kww6�!]�7?�C�A��r �\��ʹ���Զ LWfz�۟�pR�7�h��8G�z���ĺQ�KMڠ��d�g��� �3g�0�Z7-'���o~:� ��k]�gl��6��l{E-..���_���쁲��ׯ@3���4��+ӟ�����.�an� �BK�(?��3T�9岻9�ۤ����J��/�l�2	�0���On��X�[���Q$G-���1���"��.��+�I<�r�1��b3�w6xt�/�9���.��ӞD�݃9���%�r��4��-Y����b������q�0a\&�7�כ\�k�_��r��]k0Ȁ�JEk�Ps�"����i��V�޾�'L�!8�����ח�� ē`�L�N����ا���^�Z�eq2�&0D����7�Q߁B��AP7����`���dI�>F:���>~�|r=$2�O!���Z������K��j<.��lPX`����q=��0��&>~���3�q�m�D� H�{�>��5�7F��t�'2����r��ֶ��m+u�q�?\�@���u;$$���i�̉w�8���#�B�}#ds��@���X���ҝ�w�Ah��2J��L�!���ݝ��wg)AHh`-~X�/���À�lK)���w�k�������X���Or�A�������_��e�W\B�!x�ɖ8/�Mc��.�g�pUN�|��Z/{�f�L�@:�1�ʝ�M���U�#�0M
���"�2�6�9��%ig�C>:�X�q�;�4
��a�`�0RC�ˢQd����&�=|k1!7���ՒJ]ŷK` UUUv���;��]������qK�q?&��y̵ɐ��:zk��oO��E���]c6čd�u���BfHP\��,�� O��b��C���bhD�AWe z���>�KE$H3]�X����tZ����o��>0\�<��ԟqW���ppȼ�,)���v�c�_����1�`7h�}}ϗ6ʹl�����H�W ���K�NK'�Y��ȕ��d��<?P(X�l����ŋ��_�n\<v �kw+ԻQQ���I�2�嵒ϴ�a��y�5I��ny�x���Y�j���Z�+����{�c\OWN�u0�E0�d�\�d�u��x��.�2���p�ߩLG6ֈșG�%B�ص4��@[}�G�v�5D
���W��D����@ɪU�;lQ��Q�.;%e�,N�mJeg@u���b�`T���*
���$��H.?G��$�^��_�j���vT��tM��0��Uu��������nJ��'�b�8c�y��Ÿ�3j#(���_j>��Gtg�z��l�i����v R�<ȳ6W�[���ف=��@X�~�L�<J;�c��y�>48��<�ڠ�F�KS�P���]f�;6��7e.\��S�����:�6S�lM=Y�R�!�Y��r�w�[S����G��X�����)�/�C����2�8i���L�����|�Y���Sp��2�>��s�a|F�a�8�ȹ��_�����|)4ނ �܁]��B�}A�tTT)�.Z�������-�R�A'�@�7,x��1�F��:��U*`b��W�?~����(!-mc=��ed�2�$��G��~L�L�� ?�������,HU����5�Y[�.��S�	����))���>�T�=ʱb��[][[�#��7��DL�YiF��63�Y0N������7�eB�/5����߼�!��J� ئ�Դ=Y��uq�J�W >�l���Y����;�TzӲ',����Y�`5�y�)�*�x��6�O���.���g{S��l`'Ї���٢�Z����w�omsj��M�ն�HkS���Pb�j��*{�ә�O��>�@K�������e�+djWQ�f���s���3]�)�00��i���pP��/�"Hz�6���)A��T����:75Ea�AJ��]����+`�j=�ImC����z	����}����5��f�@'G���1�Im�Z�˂�^
ˈ��}
��qj[&��[2j�b�r���.'�~U�|�I�-���RǮ��i���|�E�L�s*������S�upĦ|V%yF�__��'8�3��ڊ��h�|�Я���^���������ի�Lꬾ�M.�g�9�l��|�|�����S�b<������P.C��I�;u2 }�<��ږ-!�zX�,���q@~1v�cv�4~<h��)�^����:�f[�4]��z.bt� N��>�eĝ�����`��IX�ؕ���01�nv�좏���>���]�p���6��	�/���'��>h3h��z�m���1YZ�x�xNcyD*N;4�~�?� ЋǛW̓���V�rm|}g^�3зAB���ePV�(���v;���}(\�&�***r��h��j��Ԗ@<L��x�~��w�`PJ2��#b����=0v[�3�����k�>�P�����fɇa����ev�q�a>�Ɏ��%��4��#NTE�P)X�[�u�L��ĵ	��Ea�W|:z����r�q[�.�kl���k�-F���Μ��T��rN�5��4���߸���ͭ���\�Q�ND����U���.�I���3,��Rΰ�*��.G�F͜=ς���<�����oy��W���&[kR�
�6�.&[���˰���>ve?��	u'��3�&��?>�G��Yu�WM4�YA�x$�܉̫e�O������f�-���3���ų��ā�e�h��ZrFnUǚokT�����^��GW�A�% �Y�W��������/�� �E���5~����TK����_�
6��&�]f���|�������<I�o�r�u��@�W�\�EHG�!�C$�\�z4v���@���IZ�"2}P`�(ר����L�)]Zr6�ƺ�Yz��$V_#<\8Wq\FF�Y��G	��d��,7��-g+F�z����e��w繥�+>�ڥ~!u�.(d73]S��r�F��亄9F��ށX�l������pP��6~9���ݯ���h&�s�7,U�|��7tD1�<W!�R�ݣP1O��E&��̷h����gv$,�B�q��o�����O<��>�UH��]α�%��������E>�����p#��h)i��=����؃��HHf�ZJT�
�y^kB*;�y�M�E����Ϟp63�o���;��!�%��q��н8�����M�gr�����G����,D'��SRZ4Q��!�ikO��vw!|Kg��m�l=�`�˦9:X�[X���O������kV��Nk��叆�Q-�k�A%����D�*~�槇\F�&��֘�.�$ۓ�U����E̎Aځ��fϯ[��5�$��9��A�5Q�Ċ!�"`*�Q=��9��|��� v�Bs]��ދW�ֳX[���OM�3x��������Ik��C|~*^��.�~-m���λ�{s�.�������`v%E� <�Iǧۇq'�N��j~��u���CW����.Lsw���n����0Z�3t�;L�^���"ϊGF�R��8�L�F:�t	9���H�ToO����7E)ݻw�l�L�?�7��Oe�����c�s��|��P6U��-MMɰ#����c(j��l�c1.��->����Yϊ���v�+�}#v�?F��Z��~{e�U9P�m�s��r؋��]�AS���-WG��7_��rIL)]�&�8�Y9���Or/mM�>�|�r���|T���ن�b��`�`�M�1o)p	3�!�OP�͡ӅZ��{O�&�`�������Ç���g��l�����6¸�M�.�Di��v��n���~�����rrr��~=�-��_5m-�%Q�lUv���<�zL����]�ߏ����{R���ڜ:@��ˤQ��6�}�S�lgD<�_���c~+��W���{+.�t��
)������8nX]Ӆ���Q1Uy�SA�5�����St��`�`���� H#Mv�p��g}aTcG������Pۃ�|�"TKl9ʟ�Ko�ڨ�uY���s6%��}��ht�t��Lw.:���bٱc_���:��0>Z�p�#��fuW��H��Ũ]y�A���JA�n���������� Cp�l�i�D�㞥ہ�d�2l�t�I��e�reʝB���]FS���w��������fI*N<p��eG��|�@�����53���
��9�Uz�~�"HǪ�Vkכ�f`��6�H���J����X"�(������Y�sA��b��s�[���D1O�QluG��'���oڟ���c���A�������	���I����g@L�ݪ����^$�Ǎ�Qv��-[���qg�<	�;w^B��7���r'B+4����%�Zs��w��4E"����58�
�S����z��2�q)��jzsL��Qޙ��' T��P���\���":��:M�Y^��Ҍ�u�N�β��ȥ4���klEO��C��It}tt��~~t����K�y�j�e���aI��#��QY���N���֧��XpU��˗'S2�d��R�JH��\&�V�D�޽�_���>=QIx� ;�͕�B��q��ؠ����0s�L�K-v�_w��&��U�68.J���O��&���4s�X��U�F9^���P�{_JO�PS���;4�4��4��y*����]�R���ǟ���ݫ�����
����x����ʜz�~�C�h�b@}�[ ����ԍ�����|'B�Oy�?�is%�~Pi��,��Rx�L+(Zn�bk�ʚ���b�B~k�N�CA��e��(5w6:�C}��mK���2��<NOM�W�:���}n؆e�<@5Y���U��aRE�7��ע�d����u�X�'�zY�7H�{�j�����z�mO�}�ž<!��1�� ���t�3�A�;2 �OG�ߡm@���4���$�Ff��H!X��.�����%��zb_%UN<�X�F�y��} �E�5b&���[���
�=�D�|gm�������U�Q�<��E�0S��R��<���A�Bdݠ9 t�:�����h?�Cp��&#Y)�yfbF%�c�/k_`���T���	��{��䕕;s)(��>?��;��E_���h�V��~!���^�j��E�I�7�� �8oqqq�r�ןB ���h�9�4	�:�5	YN���%�XV4Ck��r��0 n����Ϭ�5J헋V槲hh�y���eV�m�G|TY	:�|CQK��T����L�Z��&��o�v�#?����@3�]�%�C�L�|�G�4l���KU6Wf��p"�`�\��G���h-�n��$\;L{��������2�/�u��i���<�6�+R �R�;��U���j�j�Uy��"!6���<���z,��')�M�/�ޑ .�����2VM`{��������>�����ҕ��)�/! ��3�q;:	r����4���,���m�
,�[O�D�����w���g9*�-h�m�/���������}fR���.((-	��ǜͶ�����C�����"�Io��qPpcJ�n����i��)�FE�[��6ĕ��7�,�������uxc���_�***��een`.�WVN�n���6tۈ�Y��xQ���WX]N�����;C&p�V��ui�~�}b��F�9�?�f�z���BՕ���t�f��V5�RT�2�Ւ�>�~ȭs���Y��S��4�]�\ 0�1��#���?�s���F��!S�P�B�%��iy��v_���[J���&D�05m�@%E�>-�<���<��E��W�If�Ͳ��"t��D9��k� yh\�I�΋�g�M�+�`�{��cD$�״T��<\W�zU���E;��>��q[Svo���ͨ�R��v����~��$�t��L�+�l�]�d��G�µe4�s<�8/q椏	�.�X��Qⳙ�AS�m��|qd���q������p7����1�h��Yk��MT�/��v��J��[����M�� ��\vw s�ֵ�� b�G���5yK��Q���~�p<����B���^/)���r�.����X�dy�x�W��{�@fq�P���<��-�*Zo
��o��e������Q@�	�|H}�~��� ��ߚ��L��$��k_�5�1V⬪9��<k���~���Į��I��9�$h���W��S��%�I8Ȯ������Zuߩl�A�3\��6fѡ?��뺵�7ovZ�ؕ��S���^^�N���DB��l0�Fk��芦��	TH�2�e��>[�(U��C��IL'��e�������|'�(�OԱ��Ô���$�t�M2�mt1��.-Y��]��nΡj��&�)����%5Ir	�.d��lo���S�Z /bzL�%KV�D��Z�V��b�#�"
}�t.!5��u��|$�Q5-�1��Ӵ��l������zi)��>���s�Uؗ��'�D�J��gz�tVu|���Q3;;G�^z|�}}������w��K�#�\�Y4�s�F��_*�1�E�������N��C������8t��u��L}�Suuu��`���҂*��
��W��}��_Q|�5F�th:H*((�%�@U�0Z�X���{oFGG�����ŷ�m� =�fˢ�v��{UmXi��A�G�m'�� z�����r��4*Z�o��H�]�����Ql�TP hx��>�G��H��4����ن2g��aoΟ�_��n(%��&HG�=}�,�*O��K����*��k��oUz����p�֭��N�/k��*)�U+#��켔�&%�$%�d9�dГg����R^���M ����8:��� W����{6�\�\J�MPs��qx�����]�eM+�۪��zy]�DW�Ο�q���#��s*?:�"���]֊��֧��~��;vV�kΌ�p��E�#O|����gh�:��o���8_E�e@�����W�� ֢٢�T7'C��i��;�R�6��6f{	�e�k�%ـ����f���K�~U��ɥ��� 7�	��O��p�ʱYt۠3��s5�������J�vq>+��(�&�Q��=��1�A�?�Py|�Rs�{C8�\aa�fD��:|��3n�:ۗ��,�m����8L"� �R�'�Kk?��ǲ��fn�x^dϓ��s+��xA*�|�[�P����"���ȕuv.�X��p��S^��:'gX���L�@�Ũ�Ƿ�
U��rq.w��{��W	�;-�a�}U���C�櫃�f䝈Ao�3Ğ�M{%+��~�	W��:�<�L~�Z�#*��kg�(���k�Z�7�o-@3�>.�oG"l����}c�t�lk�@*PT�{����������M��3-k����2Vh�#�Aި����+!���^Ә\��
86�<{K�C>[����I�d�����)p��oS�Ne�k��~���懛�2����]�Ro<�U
ݚ�uI]��LB�,s�^Sd���'ގA0�]AI#���+�#(�v���y��j��r���1Q]]�P�'> y���XeOZ�DP�dD�9F]ׁ�3�O
�z�f{q��{�&~����:��;r�|s%r�M��Ph�~�ws`<{�9��5���y�����Uyz�^�>Wo'��ĪN���u��ɤ[�-���Ӝ"�ә��<'__�Qt��]YXJ���ҽ�AY-v�\/�%
���p�-$�i����g�������փ/�byT��n�
�f��`�r�%{�*	��`��QD�M(z%��-A$�����D3+�/dh� ��Á,J�n�������]I������o�DE޸�#��{���C�*�ɀ h�P�:-z������!m� 5��y�3��X]m��;��<,���!D���w�/?����I-I��F���Vl��m�V4q��ihx_���qOn�l�8�Lmw�m���a>��������U��rS���D�����X�fr����ZD¿�.�q�u�"����9%������YXnF)�/mOr1�b�9Lj"�ӶW��{?w���LJ\����o~�ֳ�I�:X��b�ü�����[n�cQ��ϲ��j�{X��)S���C[�ϝvѹw�F��ڪ��w�w6���L�#�$E�yk����Y����.�ڕj�l�ve'xS���G
8��5P�lHq����^�p���n�c,�ᔜ��I�ʭ�*舰�!Xz�V 3��Z��9jK�QR�����3�#J

�O]�H�3�GC;,��殗�f��o;�=+t��^��;e ���{�l1f�'Ezo �l���݈w�1Q.;�:N��n�>������G�ܹs�\�A�^�wR���~T�YZr�Z��֐��#��l&&'��<z��^�Y$v����<�5�0���F������"	TH���i.�5���q['�l�N�����L#�3n��������f��l�+�mA�V��N��9� x�:����'��ܰ����~5E���k�[��5 ע�E�Aj�u���y��)���Z@�MMJ@�3��|s(N������gA���63;�#1���\�������I����%�V�(�ZKW�S �^:�r���� �'�I�B;7���Z�5��'�$�7W��M�����ٍ�De�RXB�Y���Sh���%��`[��΀$�Bӓ��q	Ҧ-\��;�2@����;q�hV,61Qq�H��a͝8��x�M�I��`�!�c7�4�hJom�Z_Cc���L��I����c�N���cg��xu�^�w����f|V�,�@ 3�� ��E��d�H�	�nL�?
҇
�2\�ST:��D�݄T���(נyx]_ �6��Q�sW�Ű�	���-g��@���X�����:������X�
�d�aFz������==�$�	x�>���\<��ڰo.8\V�<�s3�jZ�	P~
����}�;s��^��;��4*�Z���zHּ#s��]`Cᇤ,�LBBZj�&m�`�C�%b��U/z0r���������_��Ջ� ��>����N�X&�-����@�+VO�?pl��\����s�ׇ����EѲ/�`�[Lr�|���BKQT����R���<���^8F�Ჽ��p��|.RH��\�׃��6������Oq�B��ޅ�:�
�����C"+��?���E���hK:1��R��@�"1I�ic�O�yZ%�����:�şAbi2%c^���k4����С)�+@�G�k}�q��B�9����ub���F����Z��ק~�7��#������o��U����.��	�z~���>�t#��+ �+9�nnn/W��;
F���U�}[��z( ǬD���<�6ګ����h������X��7S�����ofBf���ѭ��Q\���������	~��Yyٚ���C/����˜6C}\Nt�f��1�8���5<S���d�TC�����C����o����ε�yI�:���ކJ` �n�?�p�_pp������m�'O�X���e<:-CK෵��p1R"A��W<��}��^����C�N��}O�*/�:���>���������v.���d$�T���6�1l����ij��wa�"j>�@���3p�&7�߷�����Q;E�r]���Q%E�xrEtA�I��hi���m��@�Ħa j'6�nq,n�A�'o����8+�����9�}=�j��|��,M4ò�Bo��p�W,�����ݥ6���j�5����6	׮C�an�*@�`A��ބ�ƌ�A"]�q�҆0���x������` �
�Q�JT����rZ0�t4�ί�N5W@X����}�u?j \M�},<�XD�)R`U���~�/��KC'6����Ըg�u��ai6֛\ҹ��I�|N��֊��lL�RH@���ZNˁ�е�:p0��.�W>B��W���h�W~�a�"� P�BO�$�u�l_1rw�������q�c�\Ec����f�s9��`t
22�0�b��*$Al�ǆ�S�,��j��3���\+��i�O��,���h���yu���Ur��s����%[b��_���[�/�8ͥq��}�$���t0#�R22� Z\/�ij����qȪ^;;��*�C!��i��"�ڿ<H@��K7�<��7�N�1�4V]�׿[�9H�9��؆��؞��?.��]pp]�Sm@99�*��q�~a%�t���U�3�9|T����2<��%��I���Y�%�y��-�bZb��x�:�k����1Ϧz�3���D�u��k�~"�,�!�
}�8I��cMQ�"�����R<���yջ����ń�6���u�������6�u��K$�(��Ur0	�$�聕�6$��}��J4�%��<�~��5����oB��|cscO��H�����6V!�=}�/2~�sX�Ee�����|6�瞄�b��{wA�{�e��B]˹'��Q�UsW���BY�=��yk�Z�
�ϳ���yO� �*^�ܿ=�]����U�QO������S%wH�QΊ�(��%�^�˕~q�ضTsy�KY;�H��b��6��;-�GD�:2xh�I���/��$%�J�|���3.e����w�x`&"��W��X[�n4�����a��g�@ܡ�?<�o�� �쾈0%:�C&T��\R�?�w|zq��d�����<��X!� ��Ԏ�A*��I����*�3�f�����$v�lr���_&.!�T���_8�o��p�˟6�2�x�z]��LܠO��ɤY#�a��eŽ0tC�\�߿�B&�������K3������Ŗ�!3ЧB�y�m���b*a��$s6�s�uy4a=F���y�s��G�oe���M^R+Zm�(�k='�+@�!~E��;�!�I�W2�Ӣ�`Ɵ�i����9���'��ǧ۰��0I�eN�v����Χm����8����f��n����*��|�dbb)4���#f:\g����5��sF����ߓ�fX`ar�{�,���f�9-(�|.�u��W�'��aIBk�^D��e�2���c; h��
�z���:�bTڼp��[�C�_�kغH����V�����%���!�o_j�{#���w�$���Q�.�y�W%v�����L0��f\r����Һ�]|Ɏ���ƽ��������q�{�k�>pT�y#�y�̲-�qQ�u���K��Iyi'
;ߞ�zo���:�qpU�?ױ�w��i�_�E��'Wt$��
�4h�SIC����ƲzE�����"�#�Z�O�d�;U>@�8�ڠ��\�鹰p\\\mc#��w*􏺙�]�$��0"���x�G�������i��K�.4�9�9����+;�4���،׳���0���,f��~y��=��V�_�yO����j��-�NʍU2VQ��f/s�hVDt#%���	*�7���~�܆h�[�s�P-/y\��-�t;SB��s϶��E�%�|��,2�9�T����K���w3�걖��B�_���<�="��*7S�p���`��^
A��d�̟���4�Luڅ�M�q�{�3I!q�
�l��%-�1
�CڽQm���z��a��\]��q�U1ߪ�k�n�.���ss��y���}<6��Zr���5z�p��j�ؙ^�K1Ό��SOl��v����ŏ�<e��D�3�,�%������.�N��&�.�Kx��7r���8{s��H|5��Ӥ���v�Uۊ���7%k����;��d͚���bO��9�瓢�N�S��:�R��߻��
p�<���eQ�S{�f���6ǝ��˸�*wpG��y�~PkfBl��߆�^�W��O�	H�:C���m�FC�9)�u���/o��T�R1rr翯!�B�D�y��q�ꙫr-���͚��c�Nǹ�/�t�/�����7���8i.(������p539r�_�i���){����/���it���k���\�?�ל(��P�p���癝,�[�r��f�`Htd�6q0u1�~�d"/d��v�j�2)������I��X?����-vI�b�Wj�lK��MK�=�xy)�mKQ�to�X�RPQI��ɟ
T�l&WR�DBC�{�0%�Y6�H������.����ٱA�;������j��F[1��8o��D�7ә�~�(��B[�^D:.�Y�t��~C��K��̘1�u�,�y.J��s)�+L>��d��
����������Ī�.E���<wi�(���S�Ւ��w��&�t����S/��{.�N�J�n���Z}��8Ű\"�{l}���K�ݒk�Ī�Y8F�ק�A$jt��*N16��~_��>��d�:�2I��t5�����#X�"��*��ME��r��Kr4�R}V�W�`�,Qv�Xz��{�Mot|���y����k���b�g�:-�ŉyWN�n��dwn�^Ch����/l������g�__(���G ��!װ�1w�b賡ξ�Z�������c�������v�c}ҿ�q�(��4j8�~rҌ����Br�1����O
��gK�Qo��e�+{���Z���G|Vvv���Ս"�3~o��YT�&�d�Y��x{�'Hp=\���9:d�}��}���9�C�{��3�������?ylVS,�(���U#��ae0��3E���+=�QQs���b�h��;�W��W^t��ȗ��VΞu �/��O�*� �k��|�
����z:Qͤ�������L����1��x���7ݤC����X��o(��4+79���TD�IO�zz��Xbr2s`PP��RLI	��=>N��������"��V���)�؞�)Zl�#'rudE�9q�q��_���P���Os��<���{�f�%���G&m5�,?�|�K�k{�S��QO�� #5�9W>`Sb3׏N>B�K� M<���^p)AdTP';�R����K��6�C�K��WT|�QJq����p��.��\���J�6&`[�����i �S���r��+Kf� #�2��|�r�1���hG�%�cku���\�?��*��{{h$���ABR�Vr�!$�n��A����R�����K仃�����K��{�ϳ�>�Z|��6᧦�5�/���q��Yj���b��̞m�eڗOΠί�����
�(����7���ԧ�2d�2�A�{�8-�Tz���+�j��$��%\-���Kf��f�ǈ@?�]�ƋuLE��OR�WFmK���m������݈�K���up�gt/��c��|�!j�R�'Eam���։�yq�������q�)o�xd���$�|�m�zja8 ���ӹTU�^)R���Q��@��fggS��*eX^��J!����2���ڐB�.gՒͦ���`d���k��_|W���ϟIɫ����_�v��n ���$���`��vu�{��L��a���Z��[����Y@a{}��[����л6�C�C�*m�]Xf--r����� �N�<%Vs��@Ų����竽{�B�8a	 ��Rk�<{�F�
����fJ�	��R���%E͙�([G�� ���u;��N ��(Ӵf�aTV �S���A��u��n�.mJ� Z{
P[�Y�Nl��	F��\��P�V�遇�j��UO�;��ǻ�M� tw�}�V���é�9˴T�$3���3���-jm�5EC+� �4ğ4���H��pd�P�%P�$��H
���:ʙ�Ն�վ��U��bEp(�������&�����r`�FUt�����(��H��?�h�*,����U��Ú��1���	�բ@6���@Z6EB\�t���ȋ��FC�Y�gM_���uԫ��NQ?�m&�~�t��v����� W��S�M�,�W����U���E�M!��~�B���&G������&�+n��6nV+9ik�zGls�>�V8.�؝mx���y�4�XՐ��d'����
x�U�9�R5E�X_����OZ�(>M�ѽ�����܎+��df�]k�;ِ�q�J�L�
H��6���6`��J��ȥN9�͖IHSոo�Vy�����������^�I�\��L�Ʌ̓����n���J3Sӝ�QD�ϟ?E�>�V�)�<��h����;�_�JUQ~�^�^%����n����wh���%��*��3;c���IWո��灵���|���ay���	�"��&��	#���(l��aԘ�/��[�Zv���ugIa��q�xw���[�O6�Xl���3V5&e��>����}:���JPgD�ɉNNN �xܖ�J �c������j'fN

�fggwA��n��F��'L;B�u$o֣�7rT�C��G"Ӿ~	���ruk�$-�ˠE�R$1Y��2�e�7��㼰���U6�?̒�I��tz�MY��9�-�>���>�X�پ\�*�4ף��Q�HU���$�A��xm�ٌ���^-�����%�?2E���|.j-��Q���ϻ���7�~WC��=4�\������_�!��'"�[u ��ł����­�����UY�Y�^�zF0
[��~�#a^/
,4j�4�N������_���?�#Ľ8���G*5�tP����q�k��QCQQ������x $* h������۱WFcf�=�:(A�J���<(�`ȳ�0�u\��^�O���=B�^D%j<߭÷��s�z��rCff	�
�d&��Ȭ�G7@�]a���Z;������|R�|�����Fm�j:���Ws����g)�)��V�!���J]�O�۬���f�߉\�T��\�_]t��۠�V�'���y��^��`h����*3��ǯ�3B�S��� ������I"�?�(�puԟbȤX����a/�v>�/��2b��@6��m��'q�K!f�#�11j�RJ�l���}�s��X���SP�tF�m�%�E��t��A%�#��X�+& [^T�t�ٳjsx�@���:1��R1ӏ���D$�(b`�������ە6�A�fɔգ����8y�a�1c�&��uGU_e:e�"mh�e�I��6{E�#�F`4��7
.C��G%A���d���ޫI����W^�����
R�<:�����#h����8���������GV���T�K:y��)�o���&�"�I{�Lv{�I�$z{{�8�����57<F�w��E<��9Ur�<�ߏ�-��(Zf�U���{����Cm	i0����ݲ8�ij��@g�!�ou�D�ifT�T�]��V�V�wl�Ǧ�-�(����n~��N�ix�2��a /M����$�5^?x��"�o����L�@��o�?m��{�k6Bz�ӄM�
I�I9�aRN�K׭'�D�&S����*�=ب�)GQ	����=�0Y�|���]�|�Q�iGh�r��G}7 ���L8�̴�!��O�)ww�X]�x������Ns�>��ᥣ�S���c�Ԡi���ht�Q�Vо��g�yD�B<:'Գ�eLY5�����5��K	�ͩ��'��3#�%���^,��Ɍ�X�� `<��-ˠ�_f0H��Dx������P��1TN�����ۀ�A�>��Q>�j�<��e�R�_P��U���#%�������<Ə7��و4{�}�V_����h0�G)�XW�`��R�(���#tа�������~Ӿ�ͦ�?����{qs�kTv�jo�]TD
�:�u��[TXh�P�ק�*D���(ӧ��^R�B#���<I�\#Tp�������t��o�~�J{�Rŀc2����	׌������m��;�e�H�D���x��*�Sj�y>��z-Ow�*��j����x��!�+:-��t�هuo����K()"���xٝ��]��
긆qZU ���I�sT|�AM��8�T|���W�i��\"~dFKT����	r$BN��[��k�4�>)C%�f�b����'�n�!�T��orW������9Z.&�$�L��I,r�z�_�5�v*��V�Gp"(�1�P�����p?�p?|�&M g�K+�E
��f��d�̿1;k{��7�&;���Dp�!#@��Q]=􀟩���d�j.��W�����Db�ʹ� ����~.�s׽.19({.�yqo�԰�}��a�`)/g?���$S���:��x�y����ڂ�gȔS�&~>��23] ��
�Д�]������<��/eKj�mjC�kDt�<�P�-�i��.������u��u�R�ev�&��\wֱ���*�������	Rg�o��M�V����������K�N��⯡�<+���\/��?�M`N��^���PWP��á$���v?�vL}�ù ���ϓK��ĳ!��M
��Sq^8���j"r�n���|ұù�x�M�^2���]��f�g� ����A�S��s�]UvG0������8uz����r�]���/�����JǯG���j�9�D�,��
���c���4zb;ʪe:222��H~��vW��B�E��E�Çx��+��T�8C5o}������aw1�vj�U�2UC#���B���V�<3Oc��C��C9���S��G�-�F�,2礚�ΑSSSQg�Ǘ	qq_��κX�ّ(H�O���^�� "���@��EA9NqB�4��
 7HHh7��Ce{�@���5^_��� g��@}���7��u��d7��V��k�:,�M��ߝ�L�/?8��c��q�Yۻ9�=��US���i����B�D^r뿧ฏ������@&.��?�y��f��o|��T�bلjq���� ̏�b�J�����K�4�WE^c������1�I�:��R1� V����hE@�`J���}}}��u����m �����0��/=:v�.�K�M�}R&xEsD_�����+�|l�W�������֬$3ϓ��!6*ỏmFywZ��'�����㪟�|������X�G'�^QU�%UK!����_����N�P���*� c�-������)"D7�ۛT�T�h8o1:/h��+F����F�`�P0d�О�UV�0�kC��'���d�㐠�O�HQ-�ϼy ׮V��P�p���V�+GH�������n�݋_6�K�����ӓ��g-��Z�rt�g)�*�(?�bY���Κ�&E��	���ŽNb!�z��㡨D)�7B��H�Ȃvr�g-A8���,E^�	�׈�2W���j��Fx�e��q�^E�y���T�Z�)���)����X"�X(�޾���8��L�c�x{R���V.���C�w3[��n���(#]��6E�Wd���@�ȉ�+zt���vkgN�f�9j�`1��
m*�"ZF�1 %l�p�� Q���.6����xZ��E�.!5�*\@�����;�>z��C�|���>i��Er�v~6#�$\ �]�.�=H��y���_�]%����d#e�vhUR#yp�xO2Q��ZcF �\§Q�)�^ 4O�Q�F�)$��o%%4�U��$(	;Y�95�{�+�N>��1���Xkiu[���Q�����C�L�>5]{@�e8Y���(fU�;LLk�Q
��R�U��n����WLF�/���  @�[ �Jb=^�>�.��
X�X���TX��v%�7��	�Jco�Nf߇S�Jn�#��`��:0���Ӹ
+v�+� B�<;�!P?ߛ+c��Y����V8��^#4[�J��$�d��Z�EtM�( ���{=w���DY�t��+�^:�Hi���0/ ��u�N�e���_ q�W�DHM�/�T���C�z܅���d�LU��2�*�j���E/���+E̸���X=Ч�,\9l��\U����l�d�_B��d}&uW�̮b_4^��H?OL&/j.f-�1Nii^ݕ����\`6�������2Χ]�����(��~_\s�,�Py�Б���W���l��9���y�_�%���nRn+�~/D�z�ҝO���j͉����I.-��&"�p����t��{&��B<���Q�_Qd��~�,�@�ҟS7p�͸z�^���$�<�?q����O+J����� -Q �T�@*��j�P"���6�Z/��v2Z���Od�γ�*�\m?�.O@�c��f��lKOȀ�m�M��M�Ɯ�F��W���ʡ���5�E/�����|@��+J��Ǐ��2��M���V�gna��e.q���Pst�\CFO�}팦�V�=OZ~�Y(.������B�
2K��?�Y>i�����l��=!G��z�)�e�<�$�C~l1"�FZ�+��>��F�Ƹ��@�n�1�l/⾛����/2�wE�����*c�g�I	�>��f�~���SiL�쾥χ�eq���|T^Ia�VmIa!|�vŏ�֮��lu���j���&q��U3�)]}°�O�g$�񻪜S��m���N��n�������|*HL(�]{z�9�g�Y�Y��t-7����,����{�]���oe���y�`��������҅�뭉�̕�_u�.(6�Qz��u%E��L0sN��0��Ѕ��m��eĎ���~�`"����y��6׎���t����ɏY��E��,�_c�@�B�Rm�	:r	欟��r�qn�h�6��o��8�*$J��#�U����i���a������`>����.�	R�r3�K*ψ�IYw�EDr�3m�c>�9zu/ٸU��4�#C�
�J�=��d���zՠ�k��g�[#EUA6�S�%j<W0�%G��j'n_դ�l�B�Ц�<V��'��Hc���AX��b�C���"J^r�!+:������_�	�g��¯��P�|����.�'OF6��I%�b\m��*]��q��TP�4���Vp�
Ӂ��<�V����Hf�22�ډ�',Pn��g�}��s�*�H�=�o����GS������&���<]��c)B����WH-���6ݫV#�Zۈ�Tn<���J�A��*i��ѩ黾��P��uz����g1��kI̚���]�o�g!�u�v��QC���LΕ���o,~\I��?�����^�(��=�VB^�C��DA��W�����주,�&�2Acz�����'�
�y�kL�ՑL��H��Z>����<-@r�
[{RF?�K����OaBI%TA��d��祜�+(CBj�iUz��]�	e���.l��u{܏|�T˽ɫ�L��ՍU&���$���S��j�1�N��+씐f�44�3����+�]G�������5K�}jP 9z���n���Ϭ�]��_I���j�����h�"_?M-S��Ogj��1��C���Z|��}�Q]Ҿ����υ.�����zA�O�����f�M5�^Lᇉ4o%���w�M�=y���]b��}J,�Q?��*X"�x_�����/I�����r�̢�����b�-:5�1��Z���������4+-�61�,�8���4ae]�PN�H��_p)Į���(_��4J �S�z�����k��*�	b}���Ww�H<�����?D3�FUp��,9r�Zﳔ�qN^
nE�84��F�����D���>�0�rBZ��Pz��6�doR���؀L�ګB���ȑ����y����4�����xZ-V���k�6r���!��r�U�k�	(�_^F�������4\�}jE��B�w��/����E.)�8r��z�Q��B�w�W�������B��*�S����ɫ���pp�L�"3�\��N�	�M���w�ڊ��EHS���u$g��@:{}����[��g��}�Y$-�����K��9�n�F\��f(~
Fk7��BuӮ���#iZi��2�������(�����O�K$���*�RQy�\�r��k�����rg�<�b63U؄��%���~1�~�����uWLl��؉�f~$��[ԁ)���B:jj��<W����DW�q��Tm���I���E�����()����8H>I��1(��ѻ�R�H�LˎM�E�Zi��K񨙉������{����X���S⋳���N�'�� )N榺B���\D|N�n���s���R����%q��$!"j�_Wr(�;ȝ�f6F^J�f/�2:�j9��H��61Y�2=�p�0p��D��`�F�k�����$h��V���rך��l>d�"&I�W�+��77K�I�����?�A%��� 0��j�:�#��;]��x���X�]� Tm�j�k��8ӧU�.o2���M�c�{���)|��tm�v>Z�I�����Ց�l�h@ ���1e6%O�b��F�����ww��P��g����N"QeT�q��s��[sMu� 5�"��؇���9�9����}�������-�/>ɛM����Bp��iցa�2{WVV&|�D�,ܷUY7��Z��[�C*1��������ejBd���/��)��v3Q#�o�rO����@B?�OU�6�����{�/����.tǦ�  Ҩ|a��WF�5��W~e��¼�
�~�jf����x{q�b��h���_���=�<�%���v�|ew�q�{fP&���J�y�;S3]�U�����)C�+4��1FFSSS}�M��&l�۽��I�LF� o�oR���+��)��
�^�����=(q��/s7=a�K��Ck�<a�ak2����ֶD��`�5Ǩ�z��p�'�V++'[�_v�&ΪĒƋu�&�k�ڲ��仓_��bxe
�=��2�e�����0qѕ��]Tb�ЛӺ��v��Y�^�W����|;�����ӻ��y�C��UŎ�6�J�#��!d���?~(�2��ç���2*�ۢ���o��|�E ��O��%碛��+��WJt\p=o�෥/����(�-$ت����X��^�VB��]o�М����#����9�rR>)3��m�?��^A�"A�����U�$�4�A�wO-i,^A�;e/�et�M�ZDޣ���:9�{rO>[�灣�m[?a��Q�	ٟ�\��&�m�р@�R�暶�9�נ�g�'^�8>B<JJ��ޓr�=	ܼ�c��Ǖ��>;�gV��&jw�d4;�	ygB����#��w}����ڗH��jq�T�/�����D>�S~�I��H� ��K=�QW�v�tw_���RB�i�:�uЁ��ۉ�<ˁjg��&�x���Y�x�߳�	'��^���r��_2�E��Srs��A)��:����cx�Z���TD��t�������ଣt�U��{i�j&�~��g���1tRc���BA^�~M\�J��sL��Ӟ��m�c3������O^�����yǼ����ĵnb{l��}�n��W�����H�~#�R��L�n��nŏ� у��1K[����[x,�y��D}���c.%�����/�Q�q�y�w(-:�ž���Oiࢮ�K�mX��*��<8P:��'��"'yyE�y�'��n_f�L����|�PI�i,a�5�zE甕��)/}�n��~��)Jl>�>�j0�L;F#x
*jflF[��? ��V���d}?��
�?c&|�֖��R	��>]e����׆���d�����lLI�.տz��?`�5�r��כ��Sђ���6�3FBcW��5I�l6��F�5�Py�us^�f/m��V�K����~MQd����H�[
r�z�6j��ِX6j���:�a�1�~��ҷ^K(�v��}��a�8���s������Up�\�����Sh;���戳\c�L��|�'P��1M��?�U.m�;s�k��5Gƨ@�x?�������D�c43H�D���@IF���dvv��W�U`��㇓���K��򩝝���??}j1���)���78�3x�Ӻi;[)<�P�8�+��xq]'N�dg��G�ŋ��7=����q6���.�Y��R�:Ó]���~J��U,��&ӧ:�F�z���#dQ�=x��[�g1|bǄ��ޒ�+�!Px�����A�i��܏��"�-\$���Y�f;�z��:� ���N
�sFޑ-�)eM��� �`[����K��G�}y}��y�9�|��߇�Cp���X��:ȍ�Vϻ���3,�T�?`�����Ո?t}�&p9U�O1�c��I��b	?�p�����t+z�4�m�/W;��1��ȴ���0%xq��_�e�;���<�M��R�4�w�p�2���ʹ���/a���������!�Lt
90df�G�@.����-��Ņ��m.�x����Ϝ�o�)r*��d���5�
������Ʒ�hm��:�Cڠ�n>E<��f�ꕼ���D�£m�����	��J�P��N��-Z���叙����Z�H��8���K1U\������.�/����p�O6��S�[<ߝ�j:y����B�!a�o8��g���6�\�Ȏ~�f҅MK�\�}8k�1�]Bt������Jq���ű�W̑=L؃�-���z'O�ڭ�|�t�K(��L��mC���Л?G��m�f=,���K4�!d�ɔ���KyFR΍�kg�̭��/����Tz.�P^��Fr�+�7n@U5�fĭ��W�5f�1v���&��60��lm#Ic�Z�ic&��,��
�ߚ�H��@������r1��̲�o�)��G�{ ho�tq�6�9v��+����B�l��|ڱ�f�~�V.�
��a�Q�X<��_�E�7�j�����?ԁ�#���)�ȕ� �r��ϓ��{���q�-�:��,�i�H��A�k���A����CZ�/��I�E �v�s��!��o 4�v�S~��f�x��io��8���n8]����F�Q�U�<H���-/z���;�����H���D�� ayC-$����[��������A0���W���K���W[E��g��Г���Nb�� �<�̴ɕE� �'{��>ŅN+g�xM!m�	�	q�%�@&���^��O�.���p)L�Rv��:��*}��q&㲜������U��2y��0a��0��
p���p^���/�k��y�Z��q�D������$�L��z��,�+�y6�z������T��[_j����Lzc�A�R�"�>�'�gL�+��k��wl����>{�5P�h��_DGx~!o�Z2v��U4낒p�'Y��/gF:o��l1��KX���KB�eY�����'O.O�$����v�T��7ɂ�aq�W�d ��ԁ �Ƈy@N��'h��ˁA��-��fws}�WXȾE���2O�gR`��
�ʀ���Mz����pi��)Zyw����b�Gg���X��X��W�YV4�]��10Ì�ۇ�m鞽��ȋ�|�ƺ�G�,U��G��`�g�Fx���L��'u�ꥳʼA��ف�U���������ތ�vtP�g�yO��sm�E ӝ[��!�}a?�N��х0���RvW�^19R�:���M��z{����Ӝe���]7�zo,JC�c�)g�0db7f��]�e9ט�v��ˡɣs�>�-u�S"�ʕl��F���7��u�D���h���Зg�G���*�Ww��V-c���@#`%����.�4�+����}�1v����&��I�x��P�ff��	���m)�����)~� WI�ˢ����d��@��t����������Snf���-�����U�R�::6v8�H��0�����Vlc�]34�����U��aQU\�l� ��]�1��ǁ���~ԕ��gA`q�H�oc���+/���8k?�Dy�X�<=p�-��-9 �W����dfVE�����-�$��?��b-�"#�����g�\�� .��I���	"��s1���E2-�t�*h���}S�=��wD���W�O)n�{��[S|��� N����ǡr#��_S~+�*�:��X��wcA�4��}�q�̴u��s�ċz�`���S���,%�x�3�OL	�_忟.
���m#����Ҹ��{D_��
��`(c�;{�`Bx�}�k��;���D��׳���a껷���;�b���޺�D4o��pE%OOa33�k��o<��R�-*x��\��,�+�s����E�E%��r���OI�x�}_���Wg�Tc�%�L�}F�b�|�䆍��J�����at�����m�K/+��v���Z���r�_[�zz��y%I�_�\j?2\�x�0�\d�q��}"�Œh���y�`�v�7T�(7[����'��;g�sD>��r�#�"�]
L�cb"D��V�2�7��� �O���@���1�k|�d���!����4RD���&0-��3�=�+y0�;-惣���+o��=��Y��_��읮��6t11܎��ޟ >dk3�حe��|��6ev4��ӯ�n�	N���8u/�������_�'C1�d��o.����a@�f�  u��A�z�LX��-�/���v��������X�<~c�|ΉZO�T���mu�i� �s�&�{Ά�B��!�h	���s�
n�a	V��ij]��HO��
��%!��2�A&����)���5I�%��r�gP�h������>%᰾e{u�ٱ�wXӜ��d�|O4��M
��>�/6�Zj�Q*����R�����H�th�p��;�ncc�=���<���8)��^9�ty�^H�I|'�m�����8X�G�Bd�)0]��֟pG��NW�HZ�7����q�(�n���7���^X*���i�Oz�����ݕ�k�C+�-�k~,�>OQ�G/�Ay/sZ[%6��n��r�v�+�2��{���Jݘ\khq;˥{� �{���R�� �`G)Џ�ﵱ'#d�����b� ���>%[hY�J�[XPB�|k+�W3K+�5	-�8� ~�۫rZUt����j ~2�9����4��Z��o�1�l��~*Q)p�d�y�u���Hپ�����	wC��XH�b=/�o8�V��Se���M���QU3���ŇL���Fi3]�f	�Z ���zN���>f�>w��k�L���M�0F�$�A���j���"-tu����g�����J*7� ~��}&s���'���)=�Jӑ�(�FA9DoQ##��:�wg﬉�@���8,o���$��4��	���޻
�t�vE���1�~��jϔ���*|�����59���f��ݍp���rq�yh�rpqa3m�M��];5ll�~8'EdN�������ׇ.`��R��o)?�m�?�*}����ZGKK��"�Y��h��h�s�}7�+E�~W~�V�S�ё;;la\G���ISǟ��AD��Q] ɱNހ�U���e�	�lQy���#�������%M�a��x�װɍ���_��Cl��Vp�-u�O�����ܷ4!a��=9�H]�%�R#(��&� ����c�է]#�+�;Z��gYv�٠O"��-^��^��s�9.�E�o�n%$���?)�v��S�
���� vx<�~'�p6���97_��Y��W]%�ӥ�D��������[��xI�+Ԩ�~0kOL��h�
��#� N�;ߛۜ��633�2��fx~q��#�Z ��U^�X���<.�=1:�x��||������ D ���2
VC����q��P6��]�%z�vr��\N^��hP���pTT��<�r�:�<aOP8u9�uV��|��o~Y���l���/�b�6����j_��.rn2�^�
=�
腗�:(}���V���[NRϵ�����g���[�$�!�Y�����.����}��^i����ʨP+4��KA��1ѭ:�^�R^}��?�c���%�`吝/Q�^�m� MԨ�Q��Ԓ���@�w=qX�A���r����"k��e��$\	&�2U�����P���p>���F�_5}-�}� :;����ED�v��E ��l9'Y�R��ھTR�`|��N����daQ�ǽ��F�ؕ��rm����f�͢�3Ӎ���p��S�)rS��?��e�R-��]�2�f|��[�J��,�;Z�ޡ: X[)���^�5��RĿ��P!�f�\X�|��i"�R��ŷB��0�B(C��9��@�᱙-�x����H���:��!-n$��MkyI��u��U�� !����a'Ԁ����'v�GVq��S��U ^�K�H
Z�{���Y�M�@�:�|�2�ߴ
kq���qK~���m>���r�} D���������-\�>A_�I���W\uor�[}�M�m�tʣ��oL�ѕ���w�4����g&�k�q�M?V�VL��w�$��'�:z�^��W9��(���Q�Ѿ�����L�'$&M��[����1���#�|�t�YrW܂|G�|gT�*-�Rs8��k���X?��?=�/P%y!-m�7@CK��W�r��ㄟ��*�C쥊
���)ߓ���	#����>`���m8Um'c��B�LU擒Y����@�c��-{>'��/� ۍ� ��_>�����U�L�whI����K��7�3�-��?\��gL���������2'#)9v}tN�����������)�N����W�b'�W���"��*V��;z/\+��
��])�ɧ軜q��W߁4���������H��]�s�"�OuǮ�������awp���IQۑ�-䷰r\��Ɋ��췸"�<���K�Մ��2��ֱ�^ަ8��C�W&�ϡ&�vz7�66��O���qzrr��N�,%�ݴ���|�l�}�Ȫ�~D���0�<:jk:���E�w�Ǫ,��FSk�>�_���$����?t-�0���MD�L�dYG �rV~UXA]� ����l�^��"�+��[r��0ܢ���*��-�����y�&d	��bmݔ�j�\HݜJj�uP���5/�<� >py�ht%q�n�T�v���Zʾ�|O,�=���-�'��oG�ܕn�ӣ��+�N�8rG�Rl�������/.���	��^�]�~#�!�e�m �:�	��ͺ�����^�0���<��{PxZ�ϸ�j�'ʤ����{�C�Dg�V���| 5
���u����|�ع�����w&��}��b�5=S��[��*i=Ѣ{�c���z�B\�׶I���E�0茝 ���y?�J|���x�R+E���7htY����0p7(�v(,dă����)�L1�Hb��y��ūA��ď��j�Q�����GU��:zv�=�lNh�Sb�	ι�ʃ]5�z�|����%��]֖qu0����t�	��?1b��\	��/�˦I��^4L\��y;��O����ͩ*��
�Q�#c;=��xU	�]c��q���
�^��ޙ�Z��ǟqЀ	b���>�w�Q�d6
�@+�n(/���#�vo�I>�.�����Ξ"`�'wM�,�$Z�q�䧚�vH\�������m�hzR� F�6X�"����W#�U����a,�Q �vޙ�g"�h��-/X�<"��7Q����{����:�I��h�%o� A}���ι\1��-�;�����x�5�nt~J�`�Z����?�}?[>�޹M���`ڦ���0 6��(�ŷ�O��`����ˀ}c*�&tpF�Hz �4��Ih4���y;�����H�v|�%{}[b#s��~����׌��L/mK�a���b����������>��3TW^�C�?�BӷĶ��wU�*l���>{mݺ^4�����/j��fx�y�5��A p�~��/�_g�Oox�$=;f.\�D��z�"r���d�YJ4ŌhUx_)������9U_Q0 k����ɠ��|P�&�ٜ>��٭���\S��'�XtKw�Ūm��V���e��{�v��ȁ��	�m�[ �� %��<?��uJ˩&�6��RiK�O�F�N	z4lL����B���)g��EN�9:t�G������:]���q E-��g��1����C�^Vu4ߢ��`��6G��:�?�cr�{ī\J�?f��`r0���5���hu�P5�"��I`�8��GT�:�J�R���#���)�t��щ���u҈n��+��n��&0%ff�(�� **x#P⛚9��s�զ��7>t�O���p�x���Tys��� o�����]q������۟]a�������eXv
_S��$��ݨ��Y����x޾� �[�������<���}Y>�wTl���7�q��(ǫ��߃�=,%��U�bfy��Rwl�f���#��j�����.s�}�5?x����K�=��;2�;
R��F�Q����A�����A�G��]_	j�'��}��;���T����<ےc$O���h���"%�1lWƏ�]cw��*�{@Q��|�Mc����Z��QN�Ä����_�pTy�4�+�ޔ�BW�J�\��~+�H���sv�
j����u��њN�ha"�mM-����V
�Ƞ����i�YwqςO�7:�D���w{e�1"A7\(߳}|����nL+�n��pk5i�����o�
��6l�]�|ߣ�8��a"
{��>�
��,�L�y^���n�.�D�[�}�'(��P���6�	Z��ƛ�ы����'�}��>�L�r�ޏ"t�q����M@Z[���[p���(
,��_���y4�}r���A53�O�r��󿀡߇��g#�$""��ܕ�����q|����}!zx2U�,��!9���3Û#y�5�a�� ����Ku��8\�)��!xf�����FζRO��X|����9��V�7#� �Xm�^~�C�3���Ï
����8ϥ<=��0���W#<QR�C��ctJ�@p�`6�3��y�e���߿�X���X��y��Q֭�N�~MYH-w��'�6?��^*k'T�M��u����-M���^@U�άkE�� j-+~�H�H�x<�c����PH<��A�9M�q����hx��:%vl���ի��\���ڙ�M+�g/��0�*3�P��^+��4�-����OC(	~7I�z� �p��>b[cnPSW��K]1)?�[TXX;��۞isʛ�BG�ls�c�|뚎��l!�����J>����v�������vC�Q3�����K;;�Q^��u�E�ER��W�4���3�h�q1��+G���,qTNF����!�:g��+0����>�
Pk$N��?Ǘ@ސJPA&�� |\����"��t���/���Er�<���_XĮ�����ܳq�9h��{��������rԳhi'E�f ���������K�c�!�y0I�a��y@s�{p�@�]E"�A�z�+���>N�يvA����O�c���ۧ��	�o�@����	Њ�m�Ao���	&�&�7O@^�~�㱬�K��1�.��~��W%}M�� �J�&Xa�/T���,Twם�k,�_�0m;?�"�3��}i2��� Zi`������)=L%l����f�W�p��Bb�K$8<��Ì�H��JԨ���%��-:`��Kc�u�|(����/���;"�zC>V)��Gܼ�U�����σ�0G��.����Rή�K�3�9�&��Q�k�G�0�l���W_��!rd�!OI�3q=nGk�h�y`'B���c���>�Ѓ=�y����E�7,$c�����g$t���[�Z�Lw���;J��}�7��lFN֤|/i��e���X;��r��'�k��0��ޱs(LB�Z���=��0�p�v$�8���l�|��ۣ rc��yU>�'���>b����S��U��o8������?;�lF}�ލo�eQ�}&�� r���âQ��Å�Dx�1��H��[c�*B����JNi��.��Ww}^6�����\�ē?�X=�����2X<Th����%����!�upb[mX��$�t9�<�)3�B���.��-(���\"���4;��� wZM|崞�n�|��ʔ��Y�	��k�����V�` &�No	jm�Mh���$��.chqT	7�keL�o;�?��*�E^�{��v�uL�Ï~>r��5l����8��a�20F%:�� ��רCyhk�Q S@XL����x�~�cT����x8S�߃+Fq���r"�kA��Ќ�DCwe���a�h���S��
���a�nm��V��/ fO����
����틀 ҩ�H� "))]�!�݂��4H	Hww
�����������tɽ�L���̾g�M,#��<6���������Q-3r���⌻l�Cs#G.^\a~��*�~~a���?.��[�dA���L������)�+�օ_YR8~wr]��P�6�2.�P�s�O
�*\��u��`7)m��_4�_A�ݷ�l���p�~ �.Bc΃ U�vu[$�&6���ё��k�����Қ�H���<a���:v����BC��􆃣��q���cTD��֐\O�l~Z��Z��Q^׆-������k���)w�Z�1�&�0ڟ�?{�^��rXBGB����{���fY�my}�����Dm��	{�#I��/�\<�7������?m�����1+�&:GX5�4+� ^��z>B��^Fv�z�Gh7(��y�(,,��>���=�Ӧ��1��[��~~c-
Rx%�wD�=�@�r'p�]��>�|����t���S��e{c�|��J����L�6e1|�f8��l���b�T��u�w|���`�����.EW�{�ߒ����F����sP�"�����*�neY�SݧAS��~L�&���3B��G�`����_~�;5RBzэ�P����S���<<�0�v��}�XA�rU��S����"���[ggA�H�kǁ �=�34��[L��b<�鶑�5�U�����^� 4���D��A�_���L���u/?$�L`��x.fk�gH�5���������4��I�&ʬ�b���?J�^�3}�#Fc�á!��U��N�g�i�m8�������,h��4Cm��A"I��(���,H.l�&7s��
@v��a�sǿ7Ǎ/W��nl?Ҝ)\��)�aA2Y*����4Ǵ5����Ĵ!c��⟍�h��G\ �4����,m�b�X.����plwm��Ktj�Z�%�,��*���6�:�8�����NGJr����M��G�.j�����Dp-%��+/�N��D��Q�R�'�y���F�Ay��_|�����ī����pя��6,��;��| �3���y�4�*Ѣ���-��mjcHO�]�V�����tz6+3�%�P���㛞X恙+=Y�$��oe�<��s���A��|��g�&ud���]Qӽ[���^��X�.O�z9�mE��f�G����ywlE֓7���l��8#�Nl0�������~}�q/��c�;Y��kDx|1���p�f�ر�?����b�Q�Ao�~���r)��Z�yB�ym3=����`��7�$hm����!օ/��p\i��f��&�5���+r�[��󽛥R-����K��)�9<�Z"F�F$��<ݝ{�~��I\����rټ�b��ʤ�9n�x�������_*�ik�6m|���Ul�m�Xr����&닝LH(4=Tͻ���X�V��r�GŃ�-�-��t����=��F:��%�|������m���6J$�ι���6Y�|ު��q�o�bDyWO�G�M��{�Ɵ�T�)0��������"
!�>^���ߙ��½�x�w#C+����8D�z����Nl�5�,^8���3B;*�b�ʰ����y��~֞����E��.��۟Ӟb��U�AX���Z����G�x��$��zJU������������Fvz��~�A�����};���Q;AV�^Z;=o����A��<!�ɇ�?J�����k^�}�h�2��dC_�YL�DV�"���=��fGo%���Q��v���ȳآ#� 4�̾��4�7�i:M���d�Ey�#a�'�inoo��;A�:m+��x���D�����0�ە��sVw�g��Y�k�=LR�,2�5v���� ��)���=h�Bʠ�mD�œ8x����x��u�˵�%^�g��m�?J=�N:��u��Sb�(�VT�[��ߑ��`L�]����k����n���o�����\��������ZZ2���e�֓���r�
���S�ѣ�����e+�P��$U��y�_Y4��#ty��L.2��n[)�x���@����c:�ة��*��ޑ���y�>%�GՉ�㟻�:]Shu@��H!�[�L���Q��"��ܯ�y#"@�������_����X�ֳy\��06�Ot���?����B}RQn�shW�����!���|�C��{�Aʅw)�Ibľʎ6����9S%����A�`٧�PS[��A]RwI�
���/>��l(@�ֲY���.����^��x�k1#���N�[�?ө�cn����fфI8���y��b(�/���H����9��R����=��=�'א~��:�Y`P=ud���>�V�O�c%�_�����1�;~`Yφ"�12�Tw9����!�n�W:����mU��v������� yJO~�O�Za�,����.����!�����ܪ׻؎b�P�ތ��f ����b����Q�6a��ϲ222	7cck��kcU��WQ�����#攑k.pw:�*�0��|ԥB��
g��m���x�?����t9������>2]I���������z�h�?[F��u��_1"�Y�U1�F�b��zP�������x��yU����uU�@�Q���}䊡�����ٖ6��f5BJ���2o��m��x�f솈�N�ۋ�H|<����դS0�n�k ��x���,e�jO�_iZ7����<P�/y��쌫`��տ��kN���kg�'F�b����dú�6'+y9� ��+e�\�s������4��#
�6�5�I5��5��xc�s�Ј^ɐ�=nÕ�
��),���o*Ҍ>s�y�tѤB������`!��d���Y�,�Pv?�!���AW�Ƀ��&��f�l��ak\N��3��&6��]Ƞ��WD$Ϝ?��~�����R��֘�G5h��$T�[�S�Z7���-|�=t*�۞��Kx&2������/7v��7�T�o�'�\֏�2*�n�'�gQ�6����������6�[3/?_��A譑њJ��8�~	!@j�B)�W��4����k@� .�R"������R �7{us�ϰu}�p�͗I����c�2ࢩ��.,vW�+�S��k��.��ƌM�p��Z����F�L�}]��|����Բ)�ҏ���~�r&Sy�ګׅO��\�'ү���>�"��{������f�������ɆN��'�?�9�j�#�K8�M,���f��ז�k��c��v����(���L7~�\U�r�B^��Xt�ys}&�����)L eヨц�'q�TEI'G�x�I�B������ڦ	�jL-��b���+�\�_x��=��l�6<�&L�}��o�ߪg������_��aB���:��l�aBA�/֋�-�,Y�dL�&������Ϝ�f�������a���A�Kఔ4w�_��N�t�6��\�#�0�/�3���Y{�u��+C�H��$��K��p�J������|Рg������/*�3�S�Mz��+I������yÛx�ĕh �]T�BLl���Z�oo�s!�~�v�sOvnnFe%�������$��z�Ђ��N.���vw��}����#ix�Hja�v��_�'T����Dc�6x���w��_�����_�?��*$YL��l�-W���ֹ%�w�>9B{��m+!.������+�����F,�D"��.QKvۃ�9�"���`;��$�ZT�AJ)�yPŬ��J��e�+� �qg�S�f�Ɯs�kI}���B�����&��$G�/�-���hO�b������p�Wh:I�b�m�)?�;t�*��R�vn^�r�����y��=R��k�{sI�yY�j2�#ˍ�3}��gfhU�&d,f��F(i�3nO~�np;ӿ<\R�TT�a��ΐ�_�n�F�Ў�㳊�y�2M&��^���=ʵ~t��7~��r)��c���~���WeQ�Ҷ�D_,��"U.��4n��b�^Z��{�L��JI�ͽ�Ϝ��٫O��4��n;]�#;s���#��Z���x5�f୨�������X�tͲ�����f/�3���Y6�}��+�Nm��0f0{��.^a��YldjR���v�|ؔ�_��U���N�K=EL�侷�ZF�ؿ}ǳ�(�Kv�$p��������sr��k�����ߗ�*ԇ�Sb2�Y���h{���6��l{,_�%���f��M���rl;�u�)Kr�>������U�11�����Z���P��SG�����Ok�#���T��:�X�$٫���Du�h��4ۄ_��[�`B͏u�q�}���~������ْ#������Sh�O�*����O�p�����%��������l�ޭ�(<�y.��f1������ ,��4�ԡk*<�ʰ\���d,��Y�F�H)�t�9��)�,�۩�X�pps��3�u�y*%S��]��ѓ=�աo`�_Hj_�}'l	�~�9QD�([YSa>q<�i}��ĺ\O�.:6rONӦ4�r�LZjUVdy*�,�TS0::�I`��M�<o�3��VlU��Z���ժm�Y7��z~�Y���� "����@_����;��[��U~'���6��E蟯Y
��p;���l,������#�������&c��]����'�R<��Å��� �S�7���y��ה�(�my�d�����0��9&�9Å�9���mȍ��pņ]8�fa��$�D���RгFm_Wخ�5>�8o"���.�rrm��#�����e����j=�fɟ$��`o�U1'?UJ���å��8[���ƺ�E�0�v��ʫ�ƎX�xw��u�U�l���Uh]e	�I���fxL��>�2㾟��$|.,:���q�o̞���d��'�4ݟ1�?s��{��Nм9��}6��n��B컉�����WHBg/�&p2o� ��e�"H�8G7n:��Gi�l���@�yO���(a���U#Yg��@e�%>�z� s-�ܷ߭�@��x��J���4�YZ�9lv�K�������D��K����@��}AD�]]O4�cz�W.x��q�	����
�9�0j��-)F>4gWg6F�סƔ�6����������j��.9��
�w��g��Ǌ���3�}&�_�� nk�Ͻa��fȾ��躽q�����P�wTll�|*��D���%|���:o�ǝ���e�D��h��|����lBg �Sr|���P�8����E\�m2�:�(�@C"b�E���_4=T��Y��l����JG����_ʔ������d��*w��9�k[�U�q<���E�Ь/{"|�J����ze-��x6�&ѹ˷�'�.M�S�ܘÌ-1Ƚ��1��&�;����>W��I�}qrW*�f6��L�� �D�뭏�gcD{:����gC���6o/�ݙ���S-���	^��Y{����=,��8})��;[c_�hK��0��ۓ�NY�_D�$��rw�6c��9'_��eWv��1���?
a�L�f��8^�����_1���̂�x�����v�c��_�N�^�|γ'8x!�>�Yez=z��-�5e3´��<i�]��|�uy�g�d�k����rя{;;����R�W�Y^�`��,��o�c��~���� �z7�!+�I�g��3�G�r)P(�����1�	\Q�K�&=���潘s�����T)ݫ�H�?lEMt~���?X�v�ٲW���,�4"�BF��_���E��T��O)��`��^�� x��5�j�N* /�������[�qx�#*�l�B�
��Gs�cg�fc��Z7�ũ[ǬS�<�����вy�=D��I?��V�&H{�;*t��6D�f4�}�X�D`hJ���U
4D���<�O� �B���;�W�ΓN3��Gm�9��ٽZ�R��ֿ�B�
�{��	 �R8 ò��
놋��ˣ��rSE��9GU��rw��S�FТ_�V]�gx�� �ߍ@ �`���μ���l;���u{5�!�V��fB]؟ ̬�|�-<<<(b��C�W&2"e�G�NH��S�$&!Qs�pA.�����,����X���	��}�I����/墜��b����0<�!�Ah�1:q[�|�4)���!���\�-��
��wh�>�G�^�'�9E֝v���n�N���������%����:� ���[���ޣ�ρ����w
�/`�I ��E��������'���YIم���a� �	��-�%.�	�:S�)c|W#�2�@X�N}JIr�+�Y��ZhL���~��f�t.8�>p��d�N:�u��[�j/f���ϧ�5�jVq�lv4�'�A"w�I���i���)�5s�����a��*���-��:�33h�4�1as�A ���&A@&��>p��|�Rd�x�\]�����!d�I*2�(��>x��h���B 1�s�`���~�j��"|BV߭���U.
����t�ز׏xXQ�բm]sۯ�1{�i��;џ� �n� ����zpq
O����0�}�Ƴk�(��%Q������T���p9���{?M>�����Mb�EG���Y5^?��*n�0��Ԝۨ�|�tv�#g4��	�;�`��剺���SE�8�Ǉ�����~�@��Ѡ�#
��wJ1 ~�v	�{����}݁��G�)#S�z�+ɀ�_UF��<N,�z��zA
�WYiu�@J���'�M���$�~�+Af��# �	`�h�\��Z�8]�h�"���n�L��� �8�O�	O|}���K17����l|��W/{�g�[��\�n{���D;�i�]9�#���e�ZG��ehe�h��*��4O�.���+}��(�b���|��%��jg���N�{f'���޷G��|���Ή���r��֓ JJh�O!Ѿ��n�/)����~!Vl���E�>��ktll�W2i�U�IN������GGf��['|\�|��g͸{s%FRD�>�?:>��{Fs�D��@{���:���.��jѮ�	��=��ٶa��X{��0�1�b�-3�oe����ӆ�o�mA�k��uqs`���l�ĵ�-���f����O?�\�zד�P^�{������d�L-���*\7�@6p���#�k�S=ܯ;8�5�K;���m����l<�(ʈF�yH6�ɒ����o�j{�Ob��ǹ�
�;86͂�V��f�,��G�d��M7s*���I�6SM��\VB8'���\���򻝪�dIǷ�v�ؽ�'�v�ֿ9��;�AL��uգcUѨYe	!H�~���9)a'&��2�`��h�����NX�Qw�{fC'��o���Tt�^N������],4	����Ƶ�v��:��}�I7�����[�&�.bhO$����eU�����{ *j�������Q�H��v��`3s� �4<�c�z�29k�A�-��c�8�i9ϵC�L>���3�w���^�p��L�t�X&MF�&/~���_�=ف-Nڲ�\�A� �)�Qe��è��au�!2^gy:{��Z�I�>����,�Ul���C��|�I���L�oʯ��p���[�(�?���g�3#���� `c=��#���ړWIo}�(�<󌜻�{��kQZW�;�z�5��co�{r��(�@↸"�S�%��Oʙ[�##������ή�yʠ��nrq$��m�
#���*	yi���m>�uW��K;f2'�W0۠s��KV븣���-b��|W(E�S��Q?�@�*���� ����E����MF>�3F�#�:n+%�8掖 ��l����sb�c�����S��bdA!2?ٟ�:�3����(2TR^ΎF�7�:�0Q�f5W�8B.Q5o��4 �A	��o���=Nd�P92J ?4q��U��%���"��^� �33C���,��Z���a��l��%H����Y"tb�橲OR�!�=T)��@��R��ʀ �k(/>���vP�V�~O��v����P��b�2H�1i�c����x{�؅�r�mG�
���#���x.���OΘ�q|V�vWu�.�{����G�����a G��1W
�� Q��:�f�2��+[���!����F��ͪ:���	֍�yg�A�5l�q?��]ZH���v������c>7��������rr�����Aga���؜V�,��0�b��&-ZX;��@�s\��j��wpt�����e�<�Ҋ��T�� ��t�:S:^A�{2�{Prطo-�[d�� �J��m6
��[` �͉���SD�s1\F#J�@����'�~+������	OJ�f�s��5� �5�7�-�ry�ھ>��bh����C�d����)���-�*����,f����u�f�Y�&
y*�B�<A �4���V���`Y<Ua�:t�I���M�׍�2�������ff&�z��q
	1qP�r^Ph��)�Z�rOT����Z�b��t��@�
�[��?��I�b�I����6'9<T�A�<y�$����8;=66�2	���ݩ�-���G��5��|	�U���y���Y���|�A�7\��g�pg�ڥ.�N{�WW�BΧ�;;;Y��O�����fJ=<2�a��	-555�VZGUλ���}�R���C'�A�-@����N�x����8u�gҪ���'$49����6�*�؜�X�v��u��j(�%%��)�~`��.�>[�� ����sӕ���� W��-�A�9&G�A�Y��_��-֏�	d��l��Ҳ1��*�S�BU��Ҩ�b��J\�$�%�4�R���ζ�����e��	�v`h(O�R��	�3Jo0C. ������=<<���A�4��?"Z.=N�ר�B����b��PVZ��qS/p�C|;��`o����rˁ���ep��j��*S`a��l���2U���(헯_[FFp����>�-�B�H����#/�������Օq���=j���D���	�����Lފ(e�����\n����}(}�����_\��u<<��0l��!��	3��z�a�7:�L��� ��?�4r�mKlW;�I����Ƿvvv�ۃ	�C�j� H�ɤD���e``J�>��8hV�>/-�5�QS�b.m���,�;�F�B�899y�r~� 39Y��"b��Z72�؇X�5p>aaa�W��c�����#�N�Ò�lߕ/2��h226~���cVV���5	��Mלs>����+���֮%{\ґd��Pd�|U�x�
f	�3���i���u�̲u�����ż��lM��$0q]��-��� 2���>+oxY��F��D��O�655����w��*���M^dc�������]�uJ�D���:)+؏�d�m�ig�A�� ؤB�D��Wrr�y=ƋttN�?䥪��O,��{�n��PI$��7��R<�=~�`���OBCC%�>�F���Nu�/�Fɋ�<����0�M�*!:��ӆy!FQ�ҡ�����|$�V|QႸ)���p���F�Z��("""_`��r���p�h���>`J��W��7n@�>Ӱ����ϧm��5�3j�������½1�aI�-�!������L2��w�5=AC��j���i�J�M�Ȗ�LoL�����\j;g�0DKkk���#�ēSS�;9�5
����R ��F������S=�T�֌{��E9�{u�������ß�<�����%%Ϳ��ʇ���mo˙ʯ�t	`0���QL�/>v���0
�cc�
�	|~5�W59��Qʖ��"���������9~cT����z_�-_cg���2V�����BH!0���6H�{-�{����� u1�j^��<����A>Gis0�o��G�;aal�
Z�.8��)��Md�pO����gu֧%�e�jfl ׂ�"Q6"��O@w�CY]}��D�
G����k�SRD�( 5z����Q�-|��X�[ �_v`��=�OILd0g�SD�WH��(l�o�ֱg����#e'"����o(=��ž����ϟ#����m87�G� {Ti9��-��ۧ�r&�S*s/�_A�]u�]��0�[Gd1�闀�4l��J4Q��F��k���!�����½�:��C�	�gS{Kvs�`mΑ|�)�H���E��?@�'2�l��Q�ʏ�V���t������K"//o܎����v}�c�~W��j8t��؈� ��1�׽�l̐�z��ܤ�7������-����W�K6��XJJ�� ����c��������~���_�0�t$�+����m��\+�uQ�`�x:jjġ������NC7�7o�����;E�s0�G���Hoy`G��x�-d0���xs�pQV�ׯwo>?���[�}�$�3f�](C�6	��?�>�v���n��1Ul��<�]4)� =��c�z����],�K�k��b%��J`� �t |6�* aa���_ګ�|�
�ZO�FL�!fh� ��t9lΟ��5�W��d4]�@�2`F�J��FϡtqL?�Ѝ����@�"ϛs.��|�������'-Z|����ЃPP���Y�x�ūk��Q��x�+u�B>=X����b�V���&�����C~4|�V�T����J��� �r�Ţ&,Iv~2zV�P?EָC>9cڠz�a��s�l�#����{3�����ra444]xo����L���յ�������a�1�����1���@:ra��5mO-nnn��ӭ4"""�j��){�
���6^'��\���^;㌳5���{2�)�|�'U�cs��k�/}���c1Y,d��8��hT�j����ƶm*���k@���M�y����.\���\Q_�'�t �+V�V�NS����c5��OC?��`���J�6h��:���5��S�
3�8S����"/��$����ŕ!}\Z�󶎎������Cp�8�L�Sb6�5��h6f✫ED#G�,��$$ ��{H�\W2��C2`uؔ��M���������8��9��o�fӊi���8V*ff��1��i�Q��6%͍�7"��ÿ��:l���9'D�R�|c���jϷ��)�g��5J�_�
.9N���m۷G�R*���.��h�vl��Y,4�$iː�5������9�"��N5V��g�\�2$�e~��4N6�3Ӄ ��|������n�+)�+9"�ũ�H�L�����'��r�K��	��	���I٘�����Nמ7��D���VVV�O>A�732<\l1�zj۠��� 7���GYP���S�urK�Z�b�J�Q��&�i+�!��0�,N�(�d|}��r�\���	�[�Xk���9�����o��M#�ɞ�����jT��o��K�c]��O��f��Vp���SE�X;�uձl��I}�aV�x��L�A��p�ME�� /i�E��qNV�7���{�;н�	'�y���	t(ih�c\�+Z�>�	���4��'a7�W�9�v�)�vg� ]��M�]�fp����lw'K�#���b�|��Z��>5���k�u	���X�(/��s:�G��z�;��م�f5!�ZZI�e=#q7�6"b��I��:���2(�a�޿�s�x�gt,�h��Ϛ���r��_7TT�*���׌13�`ߌ9��q��S t������D�؉��_�&�^��z�����LG�Tͩ��P3HmV��^
�3V�
b�+jL
�����{b �����j+n�	�ݘ�D���ڪ��zL������q+�0I��iҎe�'uOE4 ����Ӱ�V%�A#���]��L�q�44� ���j&���2�%J����V����'�=F���Y!d}-�K93�?suu)�<�Y�ЁND/F6+�c���ޘJ��q_'�L���ٚ3EEE�6����QVZq��t���'r���Y|��犣U�@���Xw ��e#�9��ٱ�g����oh{���?��؝��M�+�1�=?^mb����I�������r�?~�VDT�hv&ը'��a�N��ASV�0av.��|�(og�C^�=�H�X�2��ᘾ v4:�r�#���w�=�z�_������p8]�X&����l8o�W���PS��R��rU��b�1���o�N$�މ��J��Do�yyy�����uh�9�iu,�%I徢s>�>������(r�������0�:'@�؀˹l��?|����r�P� �8��Q�3܁���?Q�����A����6�@�G�A�#!��A�-L`���9��`]��̅
��MW ��\m��zG��AA��]��3h_���'
�L�Ҿ�:�`�[�7�p��1��<7Gd�4�KREںd�%��Fw����v7�5�,,� ,�ֻe������Àq1 �B�P�7�0�\�H�(Y?�A Z�e?�?{����F�/O�2>+�����M�D^���q�^�Z�T��Smm"hD�f*-�&s���7�,��96� d�Gi����]$'$h�n>.}�
�娝@�C�_�@���|c[��gg5�!N|Q����[>�Qk�j��x�.��y��q���E@�����7K|�t-M�	!G1Yb��QO�K�ȳ����ǺBoc(u(-��
ü`��,����x�mȑ�����lp�5a�H��09�C|�rl�^�˼IY��p,vG�G<{�L������Y��W��ѷ�u��a�
���o@vI�[0����j�"jVY�fH.��0��I!���T�k?��Z�祼k|4^���{c��a�
����So333�����I��Q��+���8�U�rKe�-��N��ϐ%pn����#o2"oR"�0!g3"g��4�&�țTȄ��]T����l��*�@�1��L���ڥ���<�m������OmDҽҴ�Z7�m�
\�t�e0���聳���Ta$���	��:�X��l��\��ōC��U�:e(����q��7tUЪh��>���-k�#v4s?Fܥ��{}R���};za�:p�uj��-]5��hgP����2T�3T�&%����Ai
�&��..��]]�׎�TT�@̩��`w�̈́Ϭ���x����dE��A֝ն+����u���n�iii,n�&]2rR=��9�O�Q���gl223�9�h�=/��J���`�}�0<x?������X�B�����Q́;;v4?C5.0�����L��#r���4�I2)�T�^��`��Q-Z�x�9���������q��Pr����F�V@�U����U��NĆEN�IC`^����8��]Ҫ����5��Vi�^��IA�� m�� Q��S�rYC�*��" S�]��Ij�B`?w8,��C���&Sҷ7���ˁC̎��F�N�"J1GU��������k66QU�*�)�
��f3Zmm�j�3: }���B�<Ȁ.[�zb��-hr����ry\3��&�f.������r�뼯{{'�- � ��G��ޗ77/��1�[$��EdeC[���Ϣ6��	�F��rX��7�K	���G����|������<�V�xP��f7O��h�(�������^������Ғo�܋(�?&c����`�8Ѳ_|��?��*�?f��{��`}ull�CaUqE;��[��m�H۴B�T�� <3������N	h�-��q{�	��4�8��� C�U���/ұ.�*�~vn�����|%L�眾Hw����@]MM�̌f����ש���
�Q�u@NbJyc&��>oNƳ}���XX� ���".lg������ܪk�S|����DKK���j鋅#[h�_Kc���b���ޡ~'��Y<�f���=�t������JS��E jk1ژ�F����Z$���JA/��g�~�4y�0W;�M+�zD�)�Z���s���z>�]�s����"E}�$�`���}�R�y�b�G-��$()]��+J�'���Td�Y�}��9��k5[�7LJ}u2 (��oWNW�����u��ýgk�-eZi���������:�~���;��Q`������� ަ���r}(�0���������f��l��Iچ���asS�� d+ ��ζ�"�001�^k�Ě��RP`&�~r�ר0[L~�m.cT�@�Q̒��L`^���$(���f{w�����=�.7{UG�rS>7��@R�譗Wc�=������:�E=��a�cg{h%��m��80 �*͠�����)̎�4�� ���7.:��֦�q�_t��d�]�%����T��$�-e��.�������-ʣ�@��39��"P/b�����/egX�r�d-,�[6��� ,:�`-��o/�6'�R\��7=Yʯ�-bê�~
(km���o�ur,��v:�d���6HF�&2����N�=0�jeO�w��m,l41B�'9����s������&��Ʉ�^�������v Fs�����~H�A�=[��~G�N�����
�.�XX�@����u{{�EJ��bRA/������Ǐ%�C@�)�0��3h��;py�Q�'���Mw/kms����GX����/��4��gʻV�I��w�=1���]�~�:++���fo�gkE-w��q�o��D��P��� �i���@�����'�@�0-�T>�y죣#��jے tI�����` ���H�7d��t+&&&���/o���ΉϠ�a�������������-`I+ �ŀ��7����jL�C���3�c4OhX���BXq1ːm�Jp�q����L���^iR~7%�y��x�n:M:�/��<yb���Yr"�](���pJz��]����F�/�]�h�*<�S�7��\L(_���D����_h#�R��W��yv'�?�^m�	Ｏ�D���_��S?iW�0d��g@�S)(�mp;k�A�1Q� dR�q�%с�����x6�v�������l�����@��櫗I��UZjvi&pZ3]eɥ��/T�   P�y3�:�6WSl�֭�P�X�>΅@�[q#4"_˙��ļ��%�!ߛå?G�u������s7�o
��/���I^J�Q�p����N�[�'w߫�X�e�p�f�A�Vڱ0�w%+����_��훿���v��@,���>)�F@D4�N�>�������d��i*�d�n������c�E:::���~�5��jѻ݇p�����t�f���HHH�:�"`����ظ��h�)�iv�\�z�Ȕ�0hsl�6S.��f�@%ڃţ��o�%����t�L��w��j�G����-������>�誁����܌�."h0���I�Xfl�Pw����v)��<s��=�����&S�Q���+b������|�	�]�AF^is�;sI� �d_�i&��s�Ot<���ON��.�-i*2S�ZP5�cI���螮Y����0U�E��P:�qo�3�J�3��:�Z�4ȉ7�c����	p���`^�8/x������ԕ �u`90����)HB꿃&�e��Kl�s��`�]��[/P�������6/1o} B��]H<�-+䤗z_\�H������v`*��6�PT_`T�sp��z�JNAAa1Y]088xu��`>�^%�o� (���c2z�%&`�=��/����$b�����J�|A�sƸ��/2���d�A-��	��ߦ��Q%?�So�R�'�dd���߁�ݼ]� h�vii�s���0��k����ަB^w{o� �i��h-�#�d;�444�:M���䄄��]7��Wp�-�Q�>���쎚]^����;?�H����	���4���u�i���h��,��V���O����z\��^�y�� X�3|m�+��"�]@<P���%�o�$��%��'�zm�؇��LP��~��7D�ʪ��j;��T����\��Pr� p�r�ݓ�@���4����t�u�~Eճ�f�p=6�s9����9(t�*�%��Q/��?<2B�Z�0ru�Ձ}lmm���Q�l�k�,㾟�����n۴CG^�p $4�":���?$���H�����s��X�[�D�2�����`�2}W�4�t�o�(��:w3��E_�x�$��D^cE�6�����g�U<�z�C�������B6ŶU�yJt`v��2�����`@�k����: �{xx|Ȓ%��-�Ԗ�<Wm^�uW+�*��I5�����0W�W	��j����k�Z[��-�=�Z������M��
�چ
R�O��ɦ0��
똭�?�|��|���j�H91�/��=�̱�"ʽ $+44����1S��psqY�����K6a®`��r9Xq��,���@��/��~2v�a�}ª���$�󽙀O)�*Ǭ�E��@/�xޜ�x�����h�/"��9��U��;"`ʘ�C�x�<�>iV����>�'d�Fc���y�H�$���
_��l�*�+�2O��������C%`j[�����?  �y{ˀ��u��K����Jw4=$��	(�x3}��p���珞�իW,�E���׻>�H2�ٟ�����.C��{@��%U��n�Z���LH��r�T5|�N[�h�i�D �
m���>>�gϞE8�����=�vYB�<I�-���i[�p ����OV)�fft�c=}��!�{�-~���%��"J^.�v깙��Ew'I�<���3>�N)���	���V�����.�J��^�ϫX��%�>č�3�m�߽X�wU,��)'�!�b؉����͝�uw��D�����T�X��3p� ����_����"f�-��|��ݼ��X)!���g�7\���`�広��۟�p����Q����^3����ߜ�asڛ��)� ) ��0Z�9������@�3�Ҳ`GS��;WO�d��N��\�C��K�2�v��d�kY{��D��x������=��Ffff���)��h$h@���Ef4��	�|xx�7�Q���D�2��i��?Op_�fˋu��d�L���A/�Ԭ��l�;��i3�]�| �Ou�J�J=!�K�u�\X�}ի���t�խ H-T���x}�H�&������Z�%��wj��E���<I(k 	�M���LG2S����r� &`�n�*���	������W�A"��4g؝o ��a
�g�j{0���
f#�M��@�5zԴ���0�а�������?�7��D1����|h!�͉�!sd�p�jA�t�[nB��_0��9�v'?��.��8��sXLB[��:�K����-�O��:�E��ݫq��e�� �	AUU5C1E"oL�;�V����q�PU7�ۨ���- ]�!"� ��)�!!% %�tIw�tHJ�t#ߌ�{���﷖.<rΙ����ٳgO�pN���d)η�i`�\���lIIIC����vgIC��_ �9����xXRZj{yj�Q`dxs-�oB׍��g����Dt����ⶮY�^K�,�\8�O�Y37��PRކ|�����
zQQ��PD�6^>���a7�6��ר�	`���2�T�#RI���,M�s��(�`sM !}!� L{j>;�I����W�H��ߪ�`���t��B�?�MLC���˧3y�&���5gu� �C�|Js�q�i5ZJ��Fw������lNbw���~U&C������g��J;;�@�g,�>��ܸ�bѨ��>c��P���g� �(��������wq᳚k9=uR�������)7�|P]]ݛ7o������"*3hِBc����Ǐ-�����Ea�娩�������H����;`��N1Ov�$��>�ƞ���}Y8}aC�@�����\�ǉ��ú�3/`4CQx� �a
Z����Z�\�]�Fh����1ܙ*��F�R{�2'�1��8��U���W��,�fMԯ�x��g��r<,,9?[Fj�u��!��/æ��T�����f�2�b&��kȇjޭT�w���\�ש�u,�@ɦ��E���Y���XGCQ$��p��:C��̙�o˃�b�h�W( ��ٚ`�yta��(3�Y�p��6�!v�rø_K��2����'��k�qz�&������b�(���]�������4��x�f7�sf{_ �.6��|'`��62�brrg&�[m�
�(��F����_�V����)\����s����++q�����:k�4����Q���%"i+�l�?i�ڞ���^��Libr��HM��C��p��*��ｿy�_Q�!RP1S���䓄��W8�q�}	1�ɡG�C��K7�QbCG�E��.���*b��':���
W���>��¤�>�$#O~�����I�N�����>2��,��_}�?��M�N�K����$�8=@��~*�����8������p��
M���`�����8��Bƪa8������y�JCU����9/��N�f�4d��1���C�O�랁q��n�i)I�h����S�+�ċÏ�3q���g��㹕Կ*����k���ո4���(ǘ���F|��:��w/�����rZ#	o�Ȅ�r���zPR՗wCݩ=\I��IX�i��=��L�?�����H������uWO8�)��_�u��w`��"�[�ѸK�˂-E0��V�~��mRh4���Wd[�\:�����o_�E����g�L��(2�UrֹӒ
��,��Y7�U�ߺ5������k��n�XC%��VZ�BdF��&A{�-�m�u^�,����DQ�Uwz׆���a!��
�,T#,7WYyd�����f<nz��tu����5n�H�ԯ=��[���6��++}ShIH��M0ʓ���� �;�a20\�O��s�+Dۙ��?��ki���Iʄ溴<G��O���i��x~x����!�;{|�o���&o���3����3%e��:�"##���n!������[Y^~�>����Ύ�#�?m��F�$�m>������b� o!���˽y��2TL
��E��?
P�xx��l`"jg��.�	�{GG��/�E��Ջ� ��z�M�9*
�5ѼQ�����W-��^0W1�@̝���4��g����*B��䝹�1��뫋�RR-��\�.//��w���������3ƌ�GgN���r�/L&�S ���"��˟���}9΢��Ǵ���^?
�?�ק�ML��	K\\<�����H���x��?�@���xhzA��w��R����}��(��3"���M缲��yVj���C��4@�`8rؔ00���@H��U�0+y����C�1�΀��?�T0@��� �O䱽H]{8�&9��xhE�#q�w�`�bb�ɞ��Pz��!%&&F�H����G@``s�J1�~�eƤ���q4��<j򗙎 ���He=�ML$���Aޑ,�j�؆ZqQ��T��o�������|>���#b��y*��sBb��kL����;���}�  �3`�樂!�_]��Bt���b�9Ɯ�@٪jS)�T#����6�(�|��PY�$������$~Gxha�֑��(d���N�.om}�'��n�FihhD���n��q9������m�@���S�f�;^��0#�>��;�����} B7�������s/��1��r��n�����t�r*P�6��
|�Y#44�Pj M�s�B��?�`|�!�����G��,�L��H��E��Jy66��6�?c�Z)0O?�s���뗖�3��	 ͣ{q��1�̈́7m���s��g+���2YC��NWb���=@阘�������v�9�Q�p�@IE5���HRRR����X�f��n��,�JH�v_T�'N{:�F��p�|��r��������bdeea�/�ρ�]L����L��� �,�/G����4�T����P�b�}=�F��w�qI��[Y7��K��Q�$���--=���&xk��?ͤ`���V����@��'������8:��[F�����������ŅVY�������(�WV����OOO�0����5���V<�������Էt����}�_��V)"3Hz�o�%:�#ZZ0��}�����H՝���st�_ZZ�����"��r������Xo߾�ID�<F����a��ps�7���������F�9���^+  x��a���8�j�]^��b���3/��`����ifff�!���|#�hoH�|t-h�ٿ��q4_[NN�@�點�qo��44����E ����Ɏ� >x���=���� �w?���$%-PE_!@��
Br$��5�M�q
��`Թ����88]"l�+����ҩ8z�0���l`��@3_���Z��(�̋����=]K��0�O�߆��g\\�y�!�$��8\y��;mV�q���s������WU��@j"�7�z�R#�?��T���!������#��d��^�7#�ثW���&}�F2�A�r�_��b�'�/T�M [m�
k���;�?n�1�2��#ie+�]�zbX���D�1�����8�hg�����֞,���i�2��{f�S�7���
8��J;�g��v�6����l���3Z�Z,��}eY���J�z��HV��̌���UH�V����H�MR�o�f�x7�njsY�����dN{� ���A.]��パ�:�E�|<�����<ra���������$ZZZ� �ր��˽�*5�Y�N������Ţ����G	m޵��R�a��Z)��C�o�n/R/���Q��W/P�t`tFDBZ�!�v;���{q�;>�� �?���F�ۺ��t�H��	���$�߹F�F���bmm�v������s fR7��w�=���ia"�kW����B�8MR��oŶ7�r]t�Y�n���$��KϢ\���'B��͒���))E)OͿ���j�����l��T���$�DCCc>��p�M�j�~���Z��Lm��T����\�K5�E��a`2�1����^��MCCrǧ1��`-3p�=d����jx��F	CC�m޿�zt��m�������>�{��GF�mM��p�+"�E��M�C�too}������Dr��ŏz9t �f+d�n�֣^�h�>r�߲�jj&+,���w���!��&����:����|F���e����g�T��2Bvvɬ�((��k	��3������������LW'%���T�ZU:��\n1�ps��y������MH����l)_ø%�⊈��:0�-4����UT�_W?����}|ڻFn��L)�i��0�ÿ\c���Q2���c��>�s2B�!�����Y3�Ş=��/.Wg������3��Y��<U-p���6r�z98pssܧ���CHH���V�;�R���흝=�0\��{�V8�	'яU�<�`��苌�Cx,�Y����_�� wu��4�w���
����mmY ���x:[��J=��>x�WTT$7�sN�Q� X�g����﷧��Sx��Ż�:RK��3���m)������{UTTt~u����xqi� _N����ۃ���ֆ<�W"?�������I���/�0	��dW,fw,.m��b�@�=z ��E��� <)2��ь�/%��N�`�v�;<���|��02�'pS�͒Na�
^|"�Pj<�MVK�������h��]��� �
�w@T��ܒI�;ݩ���FP��W��7�](J-�Ϗɍ:�X��K�Y�ք-�:�e��嶞󗡵Ɲmn������7��j�pa�O
Z���Jnx�P��b��X~�������ޟqm����nvS�$�~B#�梟m\��RG���˗��0o�=���d��\����B	�����zד� I�`��Ϗ�a����&E�����U.E�
5�6�X��da�h������ἃI�!}�7LOOo��b:��A�D��j�l��G�����M��*�Wd���r��q-����������}��if���,) �D�BBd�_��3_'h�(�aʷc,|��M�����p��c�O}�!�󬑥�+�*���Y.��_�����2ͦ��i^�z�jK�����,VЕ�I!I���]�?��wp�L,��c��k������t��ۊ����7��~f���-��=:a7/�)_�7�yJ��R�1�����)�8{.�-A��D^���
�?b;=����'N5sH6����3EE��O�p����Uzz4"�Ǣl�JG�l$�50��h�T��9 �ߝ��n�/�X~q`wnV��=��L�meaw���������i�$H'�0�hRx�1L=(��:\.���G�{��S����x^F�6gԬ����Đy����}�� 76���W��+uyb��&����d�gR��d}[:(�Ѩ��fy���\h�����f>�Tw4,]���z���XT�w^i�?N��T`ά�y߿c�m��j{CS�Ty�l<��Z�*���*�W�v�䌧���k/ [����ߨ�����֭�RC����a�� ���_G3�`᎗���kT?T�U�c�x��꥝���P�fR�D�\�S�3B_�q��{zzZ�IF��k�>�S*5�����V��W�6��&G!��m��u����8c�Ŀ&[��K= i�~h�I��h;b�
&&tВ�7u���Q��πW��.}�)�K������F�	=p�y#ߝ�.�7�W��fix�W	�M�\:2L��%{4���,8������/�Z�
�h;�7�x?Zfgɂ����Dku���O. ����K@���hX�V!�s=�Vq��c�&!ٺ�������:2Ta?����t����S`MPc�������qG������M4�:��*x�	 ?���k���KRN�2I|~�7�����W`r�@�sZL�9�?��|�<���^�WI|�p[�/Ha�/�� �l�Z.�0�j]�5�Fsqa�ߛ��?���^���I� ?�>8-�p �iO���񽃂�j���n%����(((�?w�˦oPo�
FR�R;}����܊V`�`!��p��*�Qh�,:`�N��O6&��;�� /��U!��A�XBC7H,�avm�����j�"��t�����c�f �ln�6���7��ʇ �-=<:<l���xq�+$y�1t��{'��gg����L�����`�b���aԞ�&H�ż�*��ackE��6���L���֏�..�N+�I��y�׊���c�^K\\<�@�����@lZ����4����ys�m1Y���@.Y��Wq��G�׃_���?99����"��j����m<����݌E@���������y%$�l_�M�4k�G0��3��D�}��n!		�K�d��Sث���)���|8j����V@���q
3>�V�GM۱�����&s[G���D�<< ���cco��ɉ'��:�����]��7O��������VVV/%%�������6� *��;����U��c�ZS`MJ�a���`Z�I�[�(�Ж�`>�H�7_��`%�:�C�Â��K�9Ҋ[�vL�Ǩ��D�V����2�b�F�В'�����S��i���\R~ ��(V��I]+�Z�ޮ��@��F��ڣu�\�/��6^/�ٱ��~CNv͔�x��2�=���t{�7�1����]*�{@y���4�h1]����IĪ�Mp8�!�
ܘm����v�>Rl�"e��ay��D�m��n�g��OmP�4M,gj�.3TUZ�L�|�	jl�9�u�ަ����'���4&;�H�C@�l9��?�۷��ՔNX��T��r�BBHx!5�8u+���p��>�N�<���߽JP;�����J!'�N#|��X������3�� %��N~�yP�?5�IW������֣vo�p���ZH}J��������|�gwK�g�R8֟�*ݧ٣�o����}3���=� �b��M��n�w`��	I
vv��6��h�<�q$G��_����N£�X3kD�D"�uC��z3C�O$��h�D��w~O����(�x�d?D��f̦�53\��g�����mU�uV�k�\*��}N~<�e^�s�1�ddf�5���ڏ;�9o���R=}x����������}	�Se�F�r�3���L7L�M�����Ph�^��]�A�8��b1�S��{�Z�&�{�V|<:z�*E����}[��I�Z�I8���emR/t�0��d��s�R88^LL���Ϗ��K�������z�ɇ-���jKK�h��܄��bϭ����`��kBsw�_�d�?M}��;�G��V0�r�V�nFU�*/r��<���m���(�3��<D�(6��_�'Z��d�A��_]���6,���
{y�O��"!���L?�B�T&	@���S0Z�H*�.^�VL��ܪ8��&��q�]��s߄[�͇�������	�ɇ$	F4�l�_�n�jl5I/v���F~�����.��I޸����L��ݡ4q=�����E��0�t�*�<�.�eTnjj��*(+�5s:��~L�г������lmx8֋P�'o!�|V��3�Su���
�s| c��ޟY�?� HV�U�0����f�l��~///�3Z[l��!�<��p��s�&���!����)*3n=}}�2�\sC��u�qph��8=@�ge���w׆�7�k�f-��h���7��Q�8�/�-.�5��G�O׋J���E�2,<!!��T@D�Z(��5�(da��0��ZP���x!)�*J����(+7�^ss��d	��l�p�}�����,��hF-?��2�b��12�W��:�|"�\nsUR�+�ƀ[���i����6K�6F��l�.J����d��Q�\&�*���m\�l�1�@RP�9v	jjj�X�2���
5�)m����:#�v��᱑.ɓz����'?�?�m�1���E�@��L��L,y�8�))Af��"�����kG{�����/1�U��i��8�hiiQP�(��i�a�8�(�h�s��ν�r���nF ي��X�Pp$ !k4�r��F���	�S%P���~�;��]���f�B����۷ī)�U��t�XO������7��M�-o�'��m?L����A�A]Y����Q���_h���L577_:X�Gs�Ʌ�����ݽ��}�:0��G������W|ɂ���a���z��sx��s�Ɔ�'ra2�d��7s����)���퉄�| �yqqq_�>�F�����Tvy%%��aĸ��'ov/^�,c.�g7K���X�&7�	.X�o���B�y�l�sdV�1�>����W�x*��|���S������N�jWO�s�OV�U��,r�z1�]�x�~
	i6*���w|�(�5^�777}}��ay�c���{��m����z����捼��������>�D*��} �l���|���i�.<2�gbBnu�2��&�b�MG���ͨ����e��訲��@��T5u�#Ce���O0�s�my��Yg�U Ԁ	<���6�]X�d�(��---�[�1$$Q��`P\�l��8j�յ�t�Mp��^qH�>X�6����]�Tum� 4�s�B��Դ�����\&��5U�ߩciɬ|?((Z}��P착\��(�<XY����Ǿ�<n�O�FSb"	��(#�����z+��n�D_X�C��qYt�1��5�톆��2]�"����Ɓ���:�����~]l���ӧ���C��G��o,Ү��?;��}`.���#�FEAR�S!黢xq���ڞ퀙~-dq�x�Vg��&�dS�Ȑ}>`Q��9ޚH�[�v�?�,96��s��j�>p�W�������۩q�LMKk�ejJ/**�0����;���W\\����++�ut� OJ�iJ��c|<�%�/��ל/2"����Y��wUu� ���;����	+lD����a�?�b|2JJ�WU_k]����Zu�&�9y.:̟(�H�+��F����T�׼>,�L�+kQ�9��x,�����;���sr�J|�K�%&���Pu�oKe�?�z쐾���଺�~��mەU|�����OJJ�تv��X�[�!ġ	g'�y�J�s�<Q\����hh>0�������dLxh���~`1����&âhQ�};�w8���Mͧ��GF�a$�y��	�4��s������>Q�Ġ�*�*�������uu���a���<�Nez����Z����h��NLP�=;;���n	;����I�����^���������]��t273���������kqqq��-marbb~4OE�rhhH �]�5N�� gpx��t���⽉��<QVMQ0>kG��1>Ϟ/��z�7 �ߚ(���,��6Q�q���&��ȅoc&��N�8��x-@�6�P|\@`���+V��!���~�����W.L�ߟ������y<�o���=_6��!��,1�(a�6�-�8x�\����W'sH���6�G�;8X�>1Y���4B*�N�tzEc$����ׁ����p9�O���1�1�&�H�$�L��֡��2��\^��'"QȒ�6�;&@�!�������l�9;;;��wI+#���MNK�d�P��I�Nuq=*!���W@�N���1��氜�������k�[ <�Tm���32.]T�~揞�W��ξ(�]��)|�ZW�b�$=����6����4
���}�"��VJςSu����h�ïJ���L�}�+��Bx��kE�M���4���~�l,���׭��	,,�7

>��,i����'�&C�ie?_\�a�q��U!eQ��ݴ�#���� <b�=��j�"ͧ��ۜ�O����G�%�:����V�������o��v� ?Lޟ���&҅a�?66v
\���>�1L�(��j�x}k��C������/�������T�tL��I������<ޝ����3ǼW
��u�%Դblη�!Ĝb�ɧ�N�mY5k������rJYc"� R'ք	�)~���BC��K���^w'#��h�2u��Uv�<)�Y����	X�^-_�/��uK�\:��?]�2�O�e����jko�
\jAA��uƻn �淶>��02�F��F����`�3��Q�������h���p*�����?����p7������4O�j��<###���%��x�y=�y� a�-�X��)YY�vO��vvfz�!ľ�b��R;�n��=�E����ǾlAK��ȭ�b�[����i��;�|�U/���>,֗Шs�۲���C%�:��$�.W2���b�Ѽ�Q%���a��]z����0b�
�uI�'��k�ۉ����g'b�ζ}�?�Ro���V"�1zwO��t����ҳw�9�'H��_�������Zd��O�^JI-���c�����|����g�3lյ �?x����l�h]�{.���rP鮆>o�6ͫ�3W##(#����Si=w`����&�A�y�h����8��i��X�𝞟/�-�
�`**���0���.薖��<��Ƒ�4�Lb  U{e�N��a4)���w���X��MsH,l�����hZXX4������]_?��a�����#�dd,�Y��[S�h����P(���j��):���77>6�L��i�ۙ]��;�F��4E�ٮ����F�Γ�'V�w�.k$r�zI��ϫ���ڬʇTlw�d��ʔ%�6w��U\��T��y�}�,,-��< �#Y���2]쭚�DD��y�혛���z�	�žԾ���Wx�U�+ܠ����Hۖ����{�'�s����X �&Y��星�j�fl`P��tƌ� 61�gQ�ُc��Ǐ-�<ZV{��E�Acs����~x�p�00��$~|���yøo�K����F�T0�yH�0��dfg���[x�=ٙ�Gi~5� �u�Ν�)�莋10s�dv��%$�%Wo���cy�i�jn�24�����x�&NW�O��V�� �[����Z�<��.!=�����s�_����?������U>�x?oOi�6��u47����M�X^����++⼓��i����l�R�1��h�k�;"�<L̬�� _�V޾-,�mcc��gs�k^��>����~ss*v�����z�0������[ޓ&2�֬U���K���k�#�'^�Io�&/�q��-�lHВ�a@�&:����M�崸;�^�l
�e<��aR�沜�_F<�!����@A�q��T���!骼��M�	�b���22�2)B!���y������,����7mO�t�6`A��[T"]A@��������e�F��v
o�K�J����;3�[�r��+&ܱ411y�w�b��8f����&0Y���Q���Q_�������� ��v6D��� S���W/�#�N*?.��˵ �U�^Rd�`8:� �G0zQ�p�V���)12'��*q��W9	���*,�l@��D$�,���--�����Q�N�D���#�����x;�G���	0G��Ǟ�@1=dn�
���*�t�W���帤�� �;
�	�޷��|�m��X�`�i��	@�`����%�} ��F�����Xe���|}}�kJ�$���� P�<����wyf�����v	x��Ғ�\{�'"��
D��WkhT��e�������:��fT)�1}A����TYY,rۭo�CH�����>u��Ɋ��q�6H!���ֶW����X�T�xs	ɫ��m��I�u*X�u�pn�cck�y`E�������\c�p{���rɪ�Y��=�"z�[��0��%���F��P��+	ʡ_T��0���K
�Lj���p�_�c���R�1E=���μ��]6��[�*1���)ɥ1CBRվ*�߳[�x���w�	��K�`?�mAl .x[��g�}����G��h�����v������(�mmb�fv��<"� ���1����+~�%Km b�˫����)3idO�Fm@���?L�������J*zT���%݁s������H���i�"#=��wu�%T���|���XqFF���h�?�oTD�>���D�r}k��z��e�G����.���?*�V�
�Z�N�@u䅺�>	ϛ|}�ٺ@�z
n������󣵤F�vP�p�LWL�/u��,W�|h��ȏ׿w���9�z��A1�P�]���\ү��22S�<׭�+���!LT�O@f�}����ɐ1�>CԜGn񦣧��x<��z� Y0O��\<Y1 ��V K_���J�I�ϼ�F�hTkWTk}F� �,�c�R�ᓠ����$��	]�ֻR���&|%q�W��&�~��!:���wMMJ�׵���k�aI�5������+�L�?G��8-չ(��@�.��yeu�_��L<_��s�rӀ�ͧ���`�-��77��M��B�0XW?� �x���iL�{�#qS�[zke�/ �n��&����ix�lz,��$įrɼ:��
��{����&�͉�:>�A�����"JO�y�d,r3p7P@����v��̂vfj�3^���Vy�V`jas�G����a��dկ��4�K��J-��E ksk�Re£�M��'
D>��n��&i�,;3���ꚝwhu���q���x����	븄��**1���r1����J�V\%Eq����k-.)�U5D<<<\��~}&�<����2NjA�N��%F��/=#�V��n��8����YR�ƤL�^�p:�!=ޙa���C��H���<�q�:_ E8PM)7�ݱ���p��oj�^��Wl�f�c������a�9����L��.���6.����uagG�9�Z�����[5��:���"�b��o�N��Thii� K��x�H��|o�Xu�{V����7 @�Fp��L�wr"�������ϧO��/;�b�����E5��}4�M2����7T� �3���uut��/-����\V6L�E�(o�5_��X8FMMM��O8���1`m��$敲��::�kE`�my��ɼ��  g;�,_�x"�VJII=������n�X%"2���������dU�0�$No�e`6�zV
����#6{)O�10cBBp_�+�����Vqv���mϓM'W�%�)cZM~U0u�E���Cv����2N|��^����SZ���=��/�\X5#cc{��=`��`<斳�U$��4��gS�

�B�ޟE��v������?Ek�<@���MA�@��${�U��n����r��B��;�È�C�;jx>���9���2�i�wE����7�o5����p��S{Y�]��`q�X�{y9��DK�(虂TE�$�+�Q����`l��|�O�M��lM;bƵG6l��$$Dutt�OOM�4������>���Oy�W/L��ޚ,Ջ&�r=aYy��������U��&��ұ�7�Nj~[�#Wǝ�����r{x�Nm���DLT�B�j������`}$�S� ��i��8p�6`��@�����zd9UqS�H��s��uc3�\���?�-�L���6grWg��?�D)�
#�N~��c�Oc��{�\�����:<����������<z��^�Ǔ�>���ZR��Xi�v�l��e�����@2n��!�����m:O0��������ߪ���c6���E�����N9��a���3��y�������|XL\V�q���c���� v7�G��h��2kpwM撕��B-3���N�/�����i,@���Z�>d5+5�I���L(��'�HÝ;wb���ڀ)"��u ~�����Ԯ�Ɲ��Ģ�y��u�ֻ:6��v�Ya�t9�E\>|��G Q�V��,�`���Yڠ\n�ٗ�L��\�3���-/���M�8��7���b��5�tY�}��07W
���9��Q���w���Q�����R&e9l���ad̒Ub��ʀ,6����"��|?U1��'��#lC��sZ���u�`Tl5xy�.`��,��B7�(���a\[[����Q ����aY�����n�����v0rNS�L�^��<5O�8Z�Ɲ�u��;�~OIy��6�{E���J�x����G=��̜�^�3=3�ka�;�%%%���T=���VKt�b��h�"c���gs��>r�L���	VH|*;�
p}ua���x��=��K��\h�M��dQ)��)-*E�-C���ε�x 9FB_K����{l��~�}����h!g�y�.Y.��B�D�q�ㅇ|O�� &
��]�c���Ȧ�NV��2~��F�j�^V6U3t0�t�t7�4Tr�URzM�Ì�՝�q��!�B�v^�4ʷ�"2
���U��G~*�鲩�\7~	,f��G���v����0�?�d���E�n��ӧO�(�n��#|�1햚}P^��|	��z���~�躺n������}��~��R[�����@m����t��O�@j�E�����t-�A�Pu����iQ��C�0xu&�^)�ͳ4\^�#��NXC�ݺ|ԗ{s@y+�ϥ��� Sl;**�f�'}��#x7�p��x`��j�Q^�tpxP����,���[InMvnnnjn.ML��O��i"t�&$�I�/�1h���:��5AA�����>xj���Po�&��è��s"-�Ӵg�����B�ڭ*��yumHaU�D���Fy��򼬼�o�:�����勴K�+���-KS��X���L�5��K(hnW����_Sr����|�9��{y��iba�Խ~�.��x�����bM/Q��wd��nLk�����3[.]�O��jfQ俭��x�*j5�t5��J�USX �s�`0|higi֯��X�5P/���O��?N,D��9�V6y����l,,yBm�0ϸ:N.F�����$]�Z��ox��;C%qz�����,����<P\IN.���V�:���n�_5﷥����s6��)����$�(3UH�:z���o�5��}�\�{4�h�����\�6#���b'�6a��턴��ϛ���Cq}z�䔔l��9F��
/LΚ��<���8�9U �o��g���q+��x�=/.���D��P�M??���`�!�>��)�����vd'ϐx��٢��c��r�"����!_������Q8��,E��ӟ=e�ʃ�\���ן�-����%���{�F�=췧�/�����)S�y�AJy��6�E�m��,6��Cf&h� �?/����T��B ��u����%�/��P�)���H"]>kk&�Ɇ�����Rl~MER����ח�mKAA�:p+P��ɺ6Y��#<"�zf��8��gg^��i�1 �Z����{����8�����h�
1@�����Ki��ff���>� O���f��H��Ҕ�/D`YN�DlSS��U�fFs��Tl��$%+<�$���q}���d5oλ��g
���\���lzACr�4+�;a,�ԝ��Q�cQ��']]/�1ד�uttt`Eط�ܡF���&k�3�?%%��Ak�3oeqsUx�X�[��<�]��o88�ɣ\o��6�h��?u�*>��>A��E׿��]yF��?9�2+�0�#QҾd˴"F�md��4���+�J`�`�? ^�����4�_Q�$��:� ��|�{�tI`��N@����R��A�+�����a����fR2�������N�>��o�=�ŝ�=���`��pW�exd��4�:7K}�8x@Q@P�?�����dtv6]q'�8`�++��0M�P(�����6!�81)	�*��7�H�9��D^{1~Sk�0�H���#�/S$�����>wP�o��"J�f|�����q�튐�D�S�E��P�Ww�,��8��<�������ps��n��?����<��Yگ�����&<l�W�r,�8:�x�Lܽu�e̫�F�ɩ��ׇ�?��u���5Q�|y�����l4���\ܨb<�;��X��rJH�s�~�݈g4��?�6ltr�����!�R������c�M7�+C7��*��p$�;^��"��
Y�{{_���.ڦ�j�~��e������u[?�sm�;�����᱂�gF�\Q�����\�`�Z��~���Sۯ�z�����`�w10V�)�o��L�؆�#���H�dcc��n�.����)���hn���θ�

;�i�=�H;�,���H��_�>5Ǜ���v�>��m�^�R�X��N��)�����	��޻w��Xh�|�[O�Ƣ�M-��ĴS�	&Ğ6[��J�Wܐ�:���߼�dU�<c4]��4�6W����:K������^����̏�I�����EEEuLTON�Z��qW+��@�2дp��'���&�]��̒���2v�kK'7����״��eC�W-�g��XC�N|]�N���&�S��4��O�=w���7��B_�L�+>��Η�l�[[���������b�mR�w�,,�*�f������u�ffHa�����w^C�@��l 1�~D �<��"��d�N��B����#�)���ٮS7�gee�ų��>�)��R`�o��Ћt�bU&x���0��qZf�
�����a�DNΏ���SO��������+�:�ճ��<x���-J�`�������+�h}8c����)<�b����!�� �����F���E�c} �L�]*�5���9q���#,�d��U����e�$�y���Βڙ^o��7'N��(��V�S%��[�a��sY���n)����c>|�5נ���R�0>�\�$IA#?J�6Mx�V=���)*�P����x�~.�,O8+��ii�>az~��b��5c�y�gg�[�]ʾ�5-��8\*�ZL|*�{ە�'V�6�y���'��"E���K��ѷ������G3���g��8��X88�`�A]�vv0>��=�@Fz{{�@���xeee�g #�E����2�k/���������=~����ɓ'^��؊��f�	II!��T�S���AŦ�i��SQa���|�<������g�>i����:=Mㆀ�o��H^���.u<�Ot�\��XNE���G�?����O���ys�0��p��]���Ow�#D �enN�.h�c痜��x���s���+���g�]c��ɀ:������f�|W>�fOHx���UXX���	��,��t8>$^D���f�L�ǥݶk썏�'>���݄>����Ͳ1��^���y�vO}e��ވ�����X�'��I/LM������.<h�m���ŧ& ����(BlPQ?����.�{�]�Cuޜ���~G���Ht� ���o#cwժ�0i�[�ؾD~�m��]��Q)>jˌ���<N���Į5+����c��rXw
�����
@J�5��
$�?���5Jİh�r��M�.=0A��1fM��� r� ������I'��~4�bO��trBp���>�A���U3��
������չClB�a����oSӳb���r��{s���"�!�===�ɛ$CK�S2<<��?4�`$X����ҹa�)�o�d8՝��	��x��ӝ��677��Z�cbb�Д���ݫ��t��o�8������!�BH��:;���(,��ݱ,͋���4��$(~<��f��Xb��x�h�R�Gss4��jU!w���Sy��z����ߦqҿ�����V9%P��J�r�*��) �ρ�m0���d��=zj��G@w^vjԻ����M`	���)�e]z�Z�V)|�qoqs�b�,�����k�\(�����&�H��}�޽����?���/��������%E߭�WU�:�����G��55�j�)		��d�'�t�a���Z�f���@x<���4��'��UK�[W�`��ߒe�����a=|�}��K!�Bn���-P3ꀂq0�_a2t{��!����2,f�t�T�����'+���6�li~��-�~�cR<�ԟ��;�g������յe����1j�9.�Rb���3yޑ�V=��#�+���(_��݃�;�����-H�����n!��[��a����zTQ���i��3}�6-��G�\�d��^����u7urn�&��*B� ��Q���-�?+�***�Z��04��������Q(4���g����k/��n��eq���PQ[]�u��O��k��4����v͍�d�|'V��Dy��gҮ�W��~�ՓӲ�IMő�x�0������*f2��V!˫��S�.v�������-�67��jj,�_���p�'���x���#��46����ā��@i��/8����P�}�?y����8��p�(+''7�7��sp6�@����������s*CT�� O��ߣ��['��XL�{m^ף`p��Lf&zz1EEp�v,�ż��`���P���9��ƒ4�T7�R�CP�4�ᣥ�v>�<?���	`�@��O��Q�2�l�9=��iZuɮ�+k닺���9Z�#�8�qWP���%UU��倀 W�$
~��BD�Z�1������g�����B�}F��-IK�f*~�5���&��t��������b/��ي>�v^�T�Et�;��ZDC��S.@rK��022�p}#@"䥈��{{��|]��d�Z(�.���EbGn�K �s���oI�~��ML]cЃeC�����������y�j QYXX�rؘ��+�fd����X^^���������Å��8� 8���	:��~����	x���|���6���%�'[�?`Z��o]�v�ۀ��sl���2\i�:pخ��xת��18=OF��o�pDKK���/--�`�N��@����Ճq�������t��$$do�b�97�~�Ox�d;{��9�x}.w�#�u~���qy��	�T��?��A�y���ؘ̩+�λQ^= /@<�NIѐ����}�f=�[���#.����k�T�If__�hR�r%77��N5g�=5����u���Y�|?1��=///q�iݾ|��g��3bL<e�й_`X��lmך�
M�.$sp�lagW�u�S��WM����>T�2Ӂ�#q΃�+�N_o;4�&C�a�����dY�#!ڎ�]�%�HL����iD����4X�~i���xgAjz�@m���K++��������J�F�`<����?~|bggϭ�Fھ�,$�366�C��2?0:
^B#�\\]_���$�{��E@D�KL�d`8*ꀇ��>8��JV�ۘ�r�*-Z�����H-�v��(@�}�ck;�4�'7�"���az5"����o��#&�/*�V� 'ư:Q*� �����8R� ��M���;����K��fg��74�[��tS�(� ��]F�݂��]� 	�2ܞ��҆��h���%��CB�7'�L�anMЧ[Z����UX��t-Q��iv���H�&�俟0b))���Wq^��Bin���ӂU:�FO�����YY����1=�`�(�X��_M�[���'&:�����!�q�>���M紋 lf�� )�YYY�յ6��+��t�	��9�����W��ooo������
$�E*�?���Ą��E��$&&{�Ƅ�C$$�7�T2p���#ᆣJ�JR#�$=��d������+�b���dee�cN��B ?���6�D�Z�;��]���VS4Ƅ���B�XH*��/�|J����H����U�Z���Q�vO����mqDUC��)��_z:���9��O� ���"P���ʔ���u~yy��̡45n�c{P)S}B_�`Z��7����ڕ����.� �c���������o��O�7#M]K�������c�����,�5ӄ�z[_�u�̰ ɂ�;G7�A�n�����k0՘���#*q��dsqq���SY� h)y��&���(�HrE���)����rn$-M�7�;<�}��1��Sq��f�Zdd��^a��b/��������t�W{Ca!$ �d�3�x��i2�n��CM}�h\6s��~SVf��P��km���f'��1����C3�GE��=���VAm��UU��hN���������O��������EJ��� ��5m�r9�Wދ?�Mkk�)�b������T��P���<��.*.�Y't��ڿCBB����� T� �ɰ0�u���*��C�����(����;\�����AIsQSSs~�N�txΎ�A���-���}U�+;Բ?���!��Q�����S'�*��k�2e�3��%����O(|HC?�~��,*M}����:bϪ9�vړ*�N%���p�����z�of�3r��g��A�{|�yw��D�O=�
�lf����(<�V�X������B����EY�TЀ��Z���>�����rO�y�)��Z>�n����n�uB���?�i���p}8�f�u��ߧ��\����(�_��ag�P7 %�^�0W-��~STRJ$a=��{�|���;�.�[Ew��b�[��Y4~����x��;�f[\888꘲�ʟ��_��H?�b�i�����׬���{�d"q��&�uI�,�B��|���'ԣ�y�D&x��Q糳9���i.���L�����A}(<�
�����W�t���3f4�8��7Z-�������d��e�J�B��tAW�T����e�(��)��^���<�<q"��,����TSKK��>�X2���	�B��r���sk�U4���������~��������J�}�Vþ��Cۍ�;+N�Tϙa�u�dEEE�ÎH� !�!�c��gG#� ��� �	</55�/?.:�z[)l�`*����M��ۡ�����}0*T��.f��4!<��gm1�z��@/��ss�NU�j��hF 4�rZEH: *�����f��6uW��}.�-� �B�|EӑK�:W�L��Y±����Ū�	��ގ��i:��ӂ-�6����ڋ\��@н��<Tccִ饹�<Ο��y��0ũii���>���m����Ǥ�-W�W
__'35�%'�C���W�7�(�����Ք?��lK!��JK�E�{#"lK����u�zl����vwՆ'�D�J||��E�mO���ѡ�>�!��Z�/KAk�[+*����D��/Ɉ�+�PR*�4�UWt���z�@A������B�C�XV�j=^��ģ�7)kiEE��V���C}I�Y�$�]���f���~P�\D=BWj��k��א�Q:%%��։Id=��ii����ڤ�c1:��Mƥ�������F�m�;�/���.R&6�񑏚�� �M�����%qFLD�%
��������/��%�_n�;2��l��vY���K_-.6�"J��v��3Q�E[~қk�K�v�]��_����YS�I��Ɲ$��]n%(���g��d�-�X($##c:���W����i��:bt�p��>�Cܝ^��0���fc�n�11Y�p%������.8��먉��Z��*����,L\iPv5ص�W��V��}10@�E��A)��D#n��ͼ� ��#W�Q:�"�/�v�k���<��?Kk>q���u棥�=z$�k ��z'&�وoZY��%���W��Z��RUU'e�#����E�!VT���CD�\^I���edZ����Q�:$ [���VPn��Q��3��`iM��X����rb弹��ľ��[r��MR�G�����%��:6*�\\��l�8�GR��M�O�MW���5�䤇�pp#�!���1��ܣ�������%
9���:�)�!���[\���<��\O�c�~�B��ߓ<A�`��4o�t�b��m����)r�W$6P�����XJ�ntqvlpGf��NuYY�͍x����8�`�UE!�Q�!�ʞ�I4eiv���W��a5沇�%	�0�[�����?wNE��95�Cō͠�3�  $�o����.�W8�i?��0�[�;�>xD��Jl�2�Pn��A6t���A]U<���f���P�#���j�D]�+'!6�<y����G�z*����#�'�[�~��'�!;w�h���tڮv��F�*n�ݵ�n���v���K�3��u�����No E����CK��2^� �A��$����o8��	�HP~P$��2�� �u	9�e��NBp�|̭_7��P�����aրљub뮮J᥋�Fr��릋ڐ����om5mSUC%�69,8"b��g�%1yA����p8�v�������+�U*��;F�I4�����ޯ��8ޓ��ٺ�y҅����'Z�S���(�
���k'�V�C;uN� x.�ml�|�U��"g�SR�c� ��w����u�K*^/��ܧ�1�#����UH\�:.�0���&#���1h�_�#"F-�~l�TE�16�w��Ǣ�59����GL���A(������{.�L�}Qb2u�rHm %��>�0����EMA���s����pV��{I��du�����c4N��̈́�ej>���K���9::����M���C��X�(��hQ�.���1��2� ���nR����䪍cc`bXv�0J
>�=$Ô^RRr�D>�� V�#�֝G��Wֈ)���[L�9\ka��mS>>�jO0[���o/�R�)���?��������d����0>��x�p. ӛg�kl�EK�]џ��d�d�Kgv���y��x磷�s�莊�Z����-�YQ�ev�/B
���2�1��jK��o�bb�1�B�fߓ~�>y�����1G��/	�T�ߑ�715��Ds����G�h��cp^�D�x��n�ι�i�I�q1d����&=��"r<�����}{��U�¢�s6��/9����$/n�:��F��������2~Ka:Z�����A�%k�:��ر�R����:�}.���W��b�$��uʄ���QZz-_����Ap�s��Ϩ(��Ū"�l
�_z�3��ww� H��+HI	Gb1/~�a.��mW�S%����2:ϣ+lE���әST9ϊ���8r�օ|�
����Flsާ��!7�q뫆����@�%T�*�� E����-$���F�|����1v�ΫX
K���Ѣ��J��3?n��$uz���$��:<~����O��j����p �M1)3>`�'��n �]�q'5�(Oa����0����)�����U5k�l}�+ݳ0
������r�A
qr���ۅ~�k��xrJ\o�e�MS IoyIg���;]���
ܫK��Xb)ך#��<YR�uu?�m�1-�_���5D���i����@Vi�0���d;�/�<�n��H���Aխ+TP �a�E���L��'Kx!D��pT�h�0b@ڷ�w4�MQX�s >��4�WS�"��>X���]�1�ж0(N�c�LZ;0_,F�O��a�"�etcI<��W`ͣS��[���v��tr�~�}*�(�<�<;&����9�SbOz�r��pzV���/kguR��hۗ	p�o��	'ddLLLy�����ֶ6 y��9J���ˮ�o�:�AFK*�����o���͋�����}��0]�z��k ��9�R,'�����B���^h�����4�<���:��X/��Jzzz6�B9����>��T��;���!�$0���_'m��s,�����TL�����)������ζ���Ƈ܉*�)����uR�4."I�#@A �5�T@^^n+�IW��у���p�\gG�I��	������Y|d����8^��	����}�pYNON��OX�\�}�ؑ�u��7�X*C���[߸&��CxWP��iʈ�vbm�W5�)��\EzŘ�Y�J��p�l�t���U+�pK�v�	���������y�f�Փs9=�q�0�(�sE|��x�=O/���Na2X|j����V�������y�屻| JxF�/��z���h�Kf���㝙�W�/��jo���3��ʊ�R�^ie�]�8+訣k7ޡ��b2���j�л���:������*
��-)IN���O:]%��?�����r:A/׎�g9ê�g�}�����iQ���1��OUU�:���&2��}��	�z���(��c�Q���Ե3�}��Bd[I+n��� �L{Q���0�P�MQR���B?1�M5k�tc�^a@fV*��}T˹r��نa[w������/Vk/�1��w�ڎ�l�n�W �R�W(Q�V�b���T�fذ�nA���"�,�KR�Pp�r��|��v[�%���Gm�s��q�GS31B0��O�&'�X��2,��j��u�M�r#~4󚧱4�"�V@���贱,��/�NJ+#����Qm!�x^MU����W�;���4��~s{$�jA�?0��������+�I]C�U����7��;����%A݃���	bI2�i������,Cx��
E��4f�^����٭������2j ###������`�x7��{�y�r.A�܌�d
���jD˹�a��I��]H��li�[���Y�-�+[b �Lӯ�ZU-� I�Cu�-�����Ijcg�
��h	]�SX/*y-ګ��80��!3��m���8Ƞ���AO���Ig��rj� oɫ.~(tI�� /�;(�������'[_]�S���HD�6�e��X��;��e^���%D��˹��F9Y�{��k=���ݛ`���Ņ���,���_l9�?a��k��͡��Hy����p;��Q��b0��[XX������`N�zz��1��~Ra`,>��C����8TTX���u��mv��<q���F���8���V��s%
%���������9#�l��}�VA��I����Ê_d�ʭ(�~(t�7�A�z�N%d�eU��pbS����Q)���#�8�lfv��wqh�Ǩ0�@d�p	Rn�5�KM�6jRq1m����|tԛv]�(�W�NY����ձ/h�t&GL7'��J��e�A4��
ښh ڮ�?�=߭�V��8�;�1ʸI֮[��M%'1���>�ޛ���;PJQ7G*�#�^��l୩�#M�(S��6�;���� �
�F[�����j�G��.�l����|� F3J�32����S%fEr�\���������7�'��;��	j:Zƪ�1�b}��X��h�|��;��ɭ�. "������c���U�j��7��s� ����^���q�]wO���cA��5d4��"��Gz����ó�;3~k�ʻqMRf ��7ͷ�v���2�rcL�sP��W]qԿL>��6�}��V����W{��a�4�na�/P/�-�AU�^ԕ��^����aQ���|\��߳P�~s��HKG�l.Å_����)��~�ձ��ƌ8'j�yY�w����|#�����3]]\�0��q���6��(���2PE3MS���R���A����Ű8l(�.��EeZ


ayy��{dbA���*��1S4�t�.,���j�ǜ���ӿ..�
f~I�K�.���+͸�x��.�B3H97M�����V���N֬��?����|�{�����h�5����G���.[��?}G�^�"u���"P����	��aۮ��� aj�EM�}`)��3��~q�RO=\��&�])�����b��~�*�6��O������ϫR2ۿYh���Z����5�~��x:/����"��q !eD�~�~0�Bq�N�JY�/�A�F�h���!Pkuؗu���h!��-�0�q����yt����	�1�u�o]�χz��_�7���*��:�s��F���+�7�]�E�x@fn˓{zzƦJ�b�!�2"1�[��"�M,��k�:n�Ή��#a������N�̏>N2��:6��!��3]�O�A&Ĕ������EJ�{w] ��z��>'��?������p��,(o�O&E'��d?n��QE���}�뼛ŋ�)���	A����:��ɽr�vyqZS��⁌��b��(:��O���F�ۭk��� � 
�ů�1C����?����]�v��5k��>�kӫKj���Jd:�^<�G�4u9��n��ǡ��;=���"��oʭlVj5���D�9�49��D�P�\os.�?�VU[�j;=W��u���� ��h��e��3�H`�=o!���f�'x
ӣ��K��>�P\jDa&�e�G�r��{��Q�!W��i-�QH�=o*��#��V��_'�@[��sxv�.�tFa��ǿ����ݿ���7�y9�E�Ɋ���n��1�#�}b��)�1k�F�3��x��%8��V;�~Q*ޤr?k���y�;��#��������-є/����~�/Q7�������菏��W9���TiC�Ӫ�Y�[�_������^)�A(F4�`��6��\j��_A����^�ٶ�ߘ�"y�/������oc�Η_2�G�����RvYjD�1z#�C]���SS��@�L�Z ���M��9��sN���}�q�o��7�ry�z��;���S�{�g�e�y�9mx��R�4OA��{��J-�"&K����a�y\o��\;h��1w��<��nbւ�cf��x�����ו��$�C�!n�,�?��00D]=��Hӂ%AM���J=�7�<��|�ߊ�\�o:��ub��$���)5���ē�Ô⠻J#
� Â�I���U����Ks�u*��m���m�v��&qy�Wȏ��7'pն)`Pi�a��}'���r��$�aE�  VO/��k��T-��Z�O� a[Y�����o�͕98p�M�1���Z::�'3y�޴)R�<�[�pyٹ'&6.�����7�g���dv�/��
�0��r���&^T`->����гm�@g��x��+m�������k��f.+��;=AhxMhL�3�p���W6�vǾ0�:S����,��_�4\t���F���'+�@��:IR���ާ/*�4k��d;�����D���G)��,�`��Q�$ �~:�3/�NhA�E��"=n��l1?J�ED2����	[����jHb�!g{��
�I��)k*�;�����n������c\�E�he6ŝ�h������ywfeR��"�luT�V����,Hg.���bk�}U:-��)#��2~��?9ٖ�E�Y������������{ ���R9l��9~���:+����Ӡ�*�Z�fʪ��������X��(i��x�l�+�� w�I�&7�A5����Y!L�������S�F�&/������鸐h�B{��;�T	���d��/%����Sr��f���0උ,4�s͏ a��v��G�%9~GW<*Zo�y����f~��G�6&c����[���P��/44�ZF�d��_v�H���O�[�.����pP#��V�|ϻL���*ŷ-|�J�ɉv���G�~�֙�JP򏫮�P��ܮ�`)�)9��
�ծ�I9�[$��c�K��o�����:���9��z�@㈈@tR
jP�*�-��?���x���xI��}.��n�M�I=",�<�����\d�Tm�����^}R�����6V,+N�	y�%�)�x�'�����s��	�q� ��9�����{A���C42ҤRr��C�	(�	�f�EEE�!�Q�|����e�/��
z�Si��+��?GLݖ!�S�����^�E4�k�n�� ;��_� **
����bҗ��$:feI�O�e���F��Y�Q7C
t��8�dp�V�'������1�\�!a�9e��/+���5���DK&p0 aM�h#NbO���#�wSN �s9�Y�QO*��Z��q\����H��v�A���0��汱�Rb����_U]ݜ�,5ե�.��yV|a��,�\�z9�ƥ��K�a'�]QWW�Q/aS>'R죔��|qu����w���V��i<D���d�:M�8gmm��c����:EUU�u}}"�"ef�(ĩc�᯷�����Ȉ�.&	��uG��C#�D�s�ci0����f��e\.<@
B�0ګ�yFG��+��'���\��F/LPA3,ܕK�������&a ?v�HQ$�a��Fi�^'������zOlL�	��Q���0�tJ%|g�4wB@:���r\6n:�R_É��@�O�5Wb�
5�����`�CM>o;T*�4�Nm��\����Oʡ��ICf��J��>릨 ���5���� �eRm���xϛ׶p�F> ����i~Jl9U�|h;w�ٚI�GW� )T��!<�c�.���<\[��Lg���ťiXWDBY�OY���V�����#M��8y�q���2&�@��i u��,(J�:�Q�˸�^���xmg1�84PBQ��X9؁�ڼxH�M��`���{ņ���cI��R����D�����M�o;��O з�������~6���:"YX� ��@T�ę�B�	ǁ����#_�g� �v5���޼p@�ꐋ�KP��?�u8���n�^��s������BIX^�6���Mz���7Tg�����<��C{�h5��g63���"� o�*��H���k�=a���F�!m�=�=+��e8���w���և'�|��^�\�v[y��e/m���t�~
��?X�H���N����Z{���ۡ��PÃ/~'�ỈC�JTf5������z��z�d8V�����d�W$��'�I�EHQS5'�v��B�Or
��R�06�ժ��؜�-��㰽�N�ڨ���Ϯ4||ٝz^�E�o�M��'���6;җ=n�g_�}���ۿτ��*Uu�8:H���p��N��'*S.%aM(R Ō~VB�Bc��w}������\�=")8��L3�� ��%�(�\$�m�涧F��_}w��~��uZ}�P���mn��끌��xHF{h�Ǒ5ߢG���<�q���8������vP@�8_���g�؏��O��/$��8ګD�m[�K5�X^�z]]�����?�?�ש`c�����D2�
N����66���4��m.��BX'�CmL�Tj��ƨ0��ǿ��rZ\܀��A2w����[��aq�6�+J*K����wY�%�ݕ'�$*�6$�7��-୞X,�&[>���zWV!x��f�i���5�U�9�Nnu޵���t�۩�3�B�o]C�$�D��΀|���DFv��/��a6�A}<=R���KØ�.e2��N�����������k1m��)f���|�QT
	Ҭ#��W��E-�$�a�Oo���!Fx�u�<� 1h1�9��g ���#�ww伏ED�U�p"t�|U�@�\=�wkBCKd�#~�o(���`�O��|C���)���/ڝ���-t5$z��:Oh��lU��n~�����HFF&��z��ׯy�
qʸnaD��zq���s�18�"���o�¢*������JZZ<{eQWWc�(P��:�zɾ�歵��)��|�6,XbdCt{B���z�g��[Z[;=���B�����8�N/g�e9y|:?�3W6S��1#�� 0X���`z#氟-�Cqxx�;�(�3��}r���🍩�-�Ӓ�J��I�rN2F<����K��8,Dl�%��6��{��ƨW� P�y=�pA��� ً5��WZmWup@�3�7vP��oX����pԛ\.�5(���P!^�F=�����'�v��M9)����Z�z��}5��~B$䧂ڂ�~n����J���aE�N�1b�%��m��S�����1,�ϳ?���6�fuT��yAw;]l=G��Yp*샜� =�<-���C�gd�eI(�n��To�C{u�'q̕&�:i)�`Eb��7���%��먩����|�Uત������v��fq���m[�k��*Ҿn��sUq�WY�|;?������p���a�g�j|*�'̓	p7�4K��4�n�2�+D76@^��!z���o�6?-N�i�r��깝C�d>
�^�^G��krJ�$�(�ʝG��ˠ�ۡ��(B�s�|�;�2��
��J�	�1j�y���(��|��&��D�����y�v�L����GN�P�Ax�ۂ�p��4=6u�ۣ��B� ����L4s�*��C}M-UA��/(���(݃�TI ˂;ڸ<��
���'}3�!hVw@�*k�ӫ�!ָ����@+j- ��dZ(���:�<����1_�Z�Hg�y6BZ�~q��e��H��L��9S�Y�� @.��.�ֆ��i��6��i��Ct�#�L<2�����x���.?����+|~Jvu^*��|a��MՎ�� �X����ֆ�`�|[-!h�;Kۣ3[˭���p�B�Ⱥ�� -�%,Ư�?��9�`zTiC�l"���-�;C�*"�)P���W�TU����xC�=#�U~��v�TT'��Th���`��oׄ��nq�NG} <{���f����}��^��!�?>���q42q#%� 7����������B�3G�a��E/����W��Y���;����u�9�=������P��$�>yi�����Nɵa�����bbD��*4�=\p�?G�I��.z?/���,�
�*���k����h;cT6����C!$ =f)-kX�ii��@~���=t|����ɲ��T��RF������zC(%��i�u�(��S�-s�����<��q����w
<_���E�5AWr���}v����ɤ��fX�<A�`������O��R���sV�ϧU����l��"H����BR-��5m"zn���}���km�an���2R/���b�\����g/f =�|!J�t0o���o}�����<J���<&�W2���4cI9�d�e���E1=J�sd1�Y�j��鷀t��e���}����|���W��>)��BJ�/�2�����Ae�^��2��!��h~l�
�ݽ�\v�l)��I*T���Ȓ'����.jbBn�:6��x|iu�[v?���KS��K���V'V�̘��j��b�C6vMD���޽Hl���.�
�Q��!�:S,T���}�sS���qt��7����{������j���\Sdj�q6��Ǧ�U���[0�O>�ާ��q��N���ܿ�n>Mg
�X�z���,%9q��M4QYĹ��Y��襪���@�t������`�%������;��4&�C�-��6<�b�VB�Y6����1��ˁ��M�	���_es\�wQ��9��u�^������R�/G��,��O�O��pS�kPx$��&՘���nZ��Ũ�d��9�bOB恄��,睮�'�ޞf,2�S|I�$;h��n���&��ޤN����_��+~Y�L���璬#W��<v���L"�J��!�����j��D��t�������h�<oJ�t�R��5�k��TB�/�0�<өF�L2#�Z�_��^��<��
=��v�شձ1�!�Z���w��x�c�}��g.���.+a!K3>�@�F~Z�.�h���t���Rs���\w~b��י�����8>A�'�O@���7@7Λ�\�O��N�5����
BO+��U?���2A�*�<|�9e���O���5���JlEO���hap~��֠�Y��B��i^�ǫk�Wăj���u����]Г��]�<�ue�kK7�a?a~��B�"�a��lqwCƛT�Hk{�m���j3:��Ė7��W���?�c�'�I�ϳ���i�XO�sL�i���'e��3���$�:��q������4
::-�m�^�=�/%,	o�,l8t���]I���g��[�B��5�o��+�Lv0E_/T��k'B�j������u��x��Dפ�g┆��� m5h�)�Mٷ����Jr�^G���rA�ǧ�c�C�B�:�Ɍ��@
�d��U�Iݓ�tL5"���N��\��	�:ޡ̯���3aY�YǍ]������jP�-\���b!�D��{w5��QN�+�����^�����������쀊�Ko$�JI���sλܻ����
�c���ƾʘ���3��T�ཫ�"��h��3\V�*���B�_R��am)b�;A�o���������	�_��F�o{�s@z���8�{�ݱ5����߾��J�T�
8!V\]]�s$�?�I7�O]Ծ��B	��B���O��Y�o�%U1�M
D����ll���Tӫ���Uݯ�T��
��V~����U�`�o~B������k�(/����:ղ^j��Dp(�Ý`)�����)5.��QA]YEKwCA}}�T�'n�m㩪�A��t�O���<XP�8^9�+�66�"-�p�8)EY~$�u�9ܘt9��Բ"�6qBׄo�.vG:�8�)���	ᦦz`���r�q���.Av������]���ߨ�b�M�����Ԙ |��;��SJNC���U��5���"l"�Ի-��X:<��u�l�wC� -\���{�����*���	�[.%9y�U�!'�R�T	/Rm�l�Qb��n��Y��c��D[kkZ�'X� \�J~F�s�Z��G���w��$��s�![N�R%e�dO2�	y�.vK�c²�لv����Ò������w��� +��o���)�&m`L/��L�2���T{�J��$�_`��\�cn:h�F%�/�
�ã�X���b�A��ހXU:����ӷ�jo�F��D�:!m]�5o�gZ�z�z��a;	NcwW-�/�*-��G�؜� �(�����"l��RB��c%;U��R��u�j��x������r�5r�>�`����k�@����7�%�g�bʹs��?�Fع�aNO���|��)��r�X����0�E�no��p��7.��:�JV,�*`�@����� �^������#hm��n_Qa�P]ZJ�>zG�}?PT��Bf7s��C�s	2�/�]Y:�y��T���'Y��d����v�d�U�vI	��:{�I9T�7A�����H���OV�1"��޼W=ő��27�D�m >>0�Q��	O���'���������;یfr���!��)��3�C����w�%�*��;g���SE׮�� h&TD�t��h5���o��\�Ӂ�p��Z9}����-k;w�k�9�Pa�Q�ѧdG���	p a8�Fk����������?_\\l�!��C	��'����IT��B� ��/���w�2��y�eZ<����nг��5�&};���_�&�()��)�Ěb�RH��(���p���@���B�&��|�_���7�6~+��b����ێsƴUU�=�w7IlΌ��w��������C�\U��;sQUb��we��1����C��7��j��1?c
H��_o�r@��VzT�z��������F�Sj8_>��ٺ�\R�ǎŦ�F��_5���+a:D����lR��{�����:S��(�'p/�z�LI�����X� V$�U��"SIEEt�T"0�Ȗ�-�\��g�w4�4D�X �H�3|q��� ����)T��}߯_��t�}r=�SQ�ZΛ7W��O�gHk���k�>�Vܣ
w�%��s����s-P��
�۫K��L"FF:.V=p��Y��4X}��=��܄�.����g8+;�/k���X���|��0١�~S����x�Ty��(�72&-A���ɓk��M�%z�9'��Q^_��dN󟼂ر���m��P;� 7�i��;_�t��b�H��k_�����ĳm)y�a������_�Ӝ\\*��g	� S�ə
MM�=�H_&�}|�e��;��Ĝ�7g�9��ԑ���LԚ�vŃ�{#F�%K֦���f�1A�d��F�3��a�I�DǷ��K�S��m?����	����ն�y�%�f�!J���'�jv�*kw��P_m�L&+&�8nO>�v�GTԡ (``Z>��$amu�}7l�۞�X�QWU�^��R؜�ܱ��CB��6�ѫ�A��]�=��oTT{���zW�msne����p�6ѿ�Li���'/��46efs�Ox�����+E����Q��&v\�E�.�5��)���\��!:���b��	�)�j==:�^f%��>치���>���z�7�6$>$R�.¬̓��3Y��T��v�sݰ��I����m�:���r�n�V}&�C���?�0J.K�Y%�L)cޘ���r�MN��tb9���"���Wы��`hg����}Qe�ې�lť��beV��޶���f���($s=+6�s�C
����Զ���tLjK�z���X���3�>���L���� t�i�ϓBӡh�R���|6��T=�6���6=�S�� �I6�%{������gn�u�!�����2������Ua�{�#!(��aH�,S��..-1�aƙ$Q���QF\������τVթ�XgD��Vg�,!zj�	 ��)������]��u�bsv�̷T�	���An��
!�l��X<:����)��1��i����="�/S���(C�^c�uy$I�0=vv��Ʃ$�zA�Qi�>� TN�N�n���u���K�Ȼc�PG�{CR)���;v�x�BȊ)�4�w�.7Q�&EfK*N�>�y�gK�S	�Þ�SP�y�G�ݹ9$EUWBm��y����)�G��򾹙s��#�%�qB|pC�¢�>�G}�e�2�BׂP�x��D3�}�ia���s�]u�w�wBo���
�"?�5�Z�c=�����j�*���W����M�@�;\T�cC@�,uC������AO�/�oD_���ͯϲ��5�Po^9c㝹�%Z���2(���vpww���$x�w�@p�Npwww�����wx�uP5�iݽ��k��t��'<����kݱ������O�Qא�}���]޽E��C�n��N�\�S�]UЯk Y�
��SS*��9��!�C ���0�{ss��QAC��oQ>3�M*���������/�xz*��4�2��ٚ��?��ܙ�M٬���,�ք�:?����������R4�n�����W�B�hg��y�{�'���ѐ[/~ E��O��C� Z��{�F:aL��UA���<1i�v\c]�A����ۺ��E��?�=e9=�*��u��/��嬨��oKĳ�(�ozͩ����-��&�p��[]�l1��v*�VV��!�����Y�g�H"3�͕�w<�� 6��{tb���k�W�Jo	N��S�ϸ��*e�������A�J����̷O�(��gU�A���V��؄�o��D���,����P�D&��xN�@|+V|u~޹kl?o.�IHHr=�%��|�5�ԉ��Qr�eh�k;��	������le�Yʉ/z����u	�J��W!�N��Ogj�j�B�3Ŕ�5v��g#�ja��ߠ�NJ'���o���k�����s�&�q�fv�O1^7�TBK�Y2F������C_ۮ�h�4������X*�
g.z_%+�r��;���򬲲�<��M:R����?o�Ƭ*�;�s5�����e@�܇�~�O�g�Gz�$���&�)�i?68]ߝz��������"�r����)$��1*�ִ�����s2���t�P��{�ccI
��cA,הr!�}���CEHw?��9UD�����MFHb_W��\1g��2@�G�Еh2���kȔ��NX !X�c����P
���� ��.��o�"��N�qJ�G���a�.؇Z���g��o�$��hީ�{$���(��1��K�?T���8g�@�i5%�޴���s�W�([Vy�
MԠ_�ޣ�r�'l`O6?�GD�V����k@�6�[U	����"����+s���!��K�(���c���{�\��h��'֜���Z ���s��뿩YU��j�	%��L��[W���l�5����
��H�>�ڤ���:�Uɥ���|V܅X�b��bE���8�c6("�>J��|�3r�q2��sD���&�S*P�!����N�{��r��c������)�	$�`G����ڇ�=�hh��l���O��>'a�Fzcg��h�`���M�;����������SFA�k�d'�C�
��B�,(����5ym�q��Nz5#���4�[!&���J�"u��ڐ�Sn{D���}?#�xRԭ��;��C����j
�_���os%�E?�%�񎲁�P�[�*�ZI~La��$��m7Ae'��A�B@�mw{���!G�*}g�Y>�1��Nf`?2f���l_߭��a:�E�����<i�p������ObJU�� �QQ邕�)"&��>jR;���Wӛ>eV}��3�ݫA�܄�6��d�䕸	>�V?s0�Lq�M�z?�b��e��9k����}1��r!�S}�g+"bd�zl���e���od�X��'!pu��[\XX�o8� $�\�ʄ�J��{Y����b��}���n��9J�Q�[
��;���_2�N�,"��Ϭ��2o4l_H.:8�`��9`�pS#J�Ʒ�w�CÑ�M����C���vx��e<D�M}&Γ^���6�W�����k���I~Z�زM��W�S ِ&�-���������D�_s�B�ǥ=,HO�2�s��D�W�m7T�����"W �Ļ���b�'xA��	\�9m��0��q�ԏ�
`��6��R\Dи��x'��"	*�{��!�36�Y{����s��^C��iPo�+d	$۩�(e�z^�p4��9�{^x�^���Ĕ��,G�V��筏���(I�!\�E�A�2��;��ߎ0�hn?�0Ka�+��,+��՗߄�a�7 ��|P�]�{�n�\2u�6�|	"���Z񼽌�#=v�Hk}8;��$���yh�4���P`�l������e�(�����'B�/�/)�=����d(	�t̓��_��C���_�Y������O�\��>�u��1gP��aF������w��ї��q�ī%@�O{����N�/�C/��s�� �:�Ea��kT��J9��Eq�9d\�gE:�v.I&"�:�`g�8���^��{3z�q8�6��D׳>�p�ӻ=#*����fw�=^�l=����F��K�� 72�=�=�r7��\N\�97�6F�!(<�`��}K�}������&�}������(���ȍJH�T�ԇ�е�Z�]ǟ���q�g���Ae�&�/�W?Ƞ�n�듵1o�}J0�A��]�VV1&�&Ő$Kз@�ƿ�bsĜ��:�O|��5�dT�;�3唫�L�%�1���̮��An�Ζ�yڈ�vG����^��Q���R�`�S],Iq`�Y�{�ل����������N�Yp��Zl���e?@�"�n��e<�&.'�X$�Fl۳��eܺp���q&���3yf	��5�x�|K���0�&f�e���#�)M�`�/�;Һ��pU�_m���rǭ��"	w�Ջ
(r������#�F]����0f5@����%[*T7��;&$3��1��v{�d����]P�)6�pW�<�]�P�N�<�G�M�-G�A�C����~���MGУ$�Z��P+�S5���v�R�,e�{Hr���(����=Z��n��(?�Uf�^H���C=��.���!���/�q��0^ی�8<.����T`F�;�{��?�>�z��|E$�x?M����	��ƶ�����򶽿�.�8��oX����@7����"M���
�#_��j��[q=I]���Q@j���K�IJb���9�{� �Q*WU�����I_�|�g����pn5�aZ	(�n*g��;�~)E�L�]��@ٟ缶�����i�TcoX"�>�ߏ] AI(% ��Jp�m�?�Eۓ�z�=n���LO}��%I�䂪uŎڸNw�� /\~W�S�Nv��v�r#��$	���H����Zo����e��?���@=��0^���z���*!��obnj���L'뚟����P5��C���7(d�y��F,0�b�&�^�]�>W!Ң���w�e4C��ѷ�B!��p�d=m*��ڰ����4q$۱��ٵ>K���mo[D��',�Z0�`D��G�м<T e�2j�&m��
z�����
J�(Q��GM�|G�1Z��6�nr����tY��> ��ͰS�\_O���F�1\3������x�@:<_����L���*g����
���B�Up?�ԥK�	����R�c���g�XKm:�w����Ĳ����{�T.�(��|���ʟ~�jr���t;5�l�N�F@����dG[uµn"���ziN}��Ƙ�h�w���V.����A�k9a3���D*���GQ�-`��/�=�t&���=t6��K@�j��T2�I6�/P�r"Ji��!ԩu}*�#�m�se�E����[��o���M ����l�6�4�0�:����������P
�L@�Ǧ���s�$x�����d�g�̈́�x7���\Gd��1����;�)��0�wһE�i�@=W%�(R_��`zcC�A�XѾ��� ƹXmT�ɁO�	�*�Z�pS񣮾�@$�}�f� �P�����6|$> ]2�4����Uw��3���iSu��T��tR��1s(}kF�=L#6��M��dݱ�y�@�!$���:f��fJ|c7�@˩z5�5蛯A<�^�?�GCq$�����S��)�%���2��?jΫTi��+�3
0���q��ڰ��UL�H�D��鱾�E	;��~�3�W	��i��M���q��D��`���7_"Ԗ����4df�v��cEҭf��hʧ��c@�Ǣ�ŏ�ם�w�IR����9�����v���w�f��y�9����Y{w�L�$I�,].��T|T�e��z��Q�7F��T=�U�V��2�����%"{0��U&�-�iI�b�c�
C�.=�u��0vH?�����`P�~�(=��-�{�"�M��W%����S���Mh1�ag 
�"�)b|�Z�Z�@uT*��t}��2��M �4i(g�wGTQ���U<f'��2ov��c�����KN��5%x�.�]����mZ������;+8���A?z.�
�4Y^�!*�we{�%��;�	�Faqu�!@FE�f���-�2��0c��m�����k��sm3����������-���@��ɣ=@�Q������R͞M�/~��Bo�d�9���$8u��,G���.���*��bF.�<��Ke�tW�2�4�KB�\O���a����k�  !�*M��	X�z�y���G�� -9�m[�EG�����½��>F(ڪȀ?���!���g�>Bt��1U��ߗ�B��"�	~�:2I`g�=\$�B)�L�2�e�g��N�_ G�#��w������*0�6HÖ��[�B0���q��ie����C���+Z�����۔��i���u����,V>���q�/���::�H�+F�����U��4��UH�����=������h��A�w5@Y�%ϻ���	���0�������K�n�0[m�ME�ǯ�'	D�_�/����k�ᥖo��d�YT�+�a8"?��"�æ�E�����8����7~]�t6Άh�͕����Y��wF�V��
u���kz�����|�A��-� �Q�JV5���p��h�������_�4L��(����H9�3&�J_; �.v�~���˓B�%�w;�y����9�z)����, �|Yh���{�e����{����Ǐ������8��=������JxE�L�Tw��8I1��Du�ć$A>;}�*�XT4�h k��q��iH{�$�2����w� ҏ�PR��t���M6�<��&I+��FR�z�dr��҈TS-�li���N�Exs�"��V����^=�qbF���!6Ǜ�08��Ͱ�WPP�#A5DF��bY��4���dI�2Hm��A��+�T�i�����w7t`�B@��SfW�q�FzC�-��h6����\���&��jH�'�e��6�_D�[i�	�Z:6������m�M�#�i��u6�ߤ|xs"�U�u���͉�4�ȯ)	����[_��Þ�8,�6+^�l.�AXFw
�O�!V�p,�ޒ�!�!����n�lz�.��M�#yDZ�E���2�&"�7�D�������)�G��u�s��v<���߿q��ZR�ZI`~��ɪX��W�N�}������d�t��P��T���͊�����\���J���(u�������g��Bbt�-䮟@>�A#��9�_/&�Lπ8��r'�����x��Ľ�2�o�[�LOΚ%1�8�h��̻��DQ����@���	L���P����!�|��Q1J��GMM=M��sW߿�W�Tj�ڿ�����8��qׄL�+��Sé���M�s���t;��o��y��\���In�/��T$�^��K�O���ٺ0`����5#N��c) �]��/L$W F�Jb
��θ�dN��Ғ����/�Ƶ"����d����N��&��&NNY��::a+����0�/�/�9h���XD���SD�f�ċZ%%�b�v�=l����HU~�L�A�ǇA�-A.ب��\Ӱ�Zk@EQ����C�Ɨ�bw`����_���N�D�/�jvk�`^���jЛ��W�1�o�u�y��5�j��)�z�ˣcU���Q��|r�ܺ�u���~�Bf
z�熕u`�Ċ�j"ȁ���UJ���^���o��b|:zN�e��
��X�CH��8�tu�]�������k�d-�:!�^�ɹ��qk
��٧�j��-��k�ܥ�	W��忪\p\W�X����Y\q��&��ߎ��hfg�ANx�_⌝l��S籭%>r*Y�?
�ۗdzҨ���P��y��I# ��$��((�7�һ�rR���֧�MZdr����};�w�65(\�Kͽ#�xxt]O�Y���mGT��(4o�EGs�)����ȳ�4P2
h�������D2Ut:d�*��(�춶�?_��z�l�xr��Ɓgo\F|d���@_-&�BR��A]��C�a�������7�����Ѧ������G_ج�)7HL��GBoU�������|�iK���rlۍ6���]���҂LB��b��
�:555t+�ȓkk
�U�����aWk��ft��,��q�rU;��%���	F�@ZM��*}�-'��$!��)/���6�6����?#
�h�8}H�Iܜ�Gra&Y��!c���;d�����FO�UC�*�]���)6�7v�ı��Y���.?�]��@x����;c��H��Ӿ��K�[W��e~�{n:�ӟ��q��8����kh��0�n��\6C�u����Ͷ���N�ձ���o!h�d 0X	��_#���d�;�XH�%�uۃ6p���`i�5$�|���9.6�#K��g$A�>rr�9�_E����P��Iljjj��>�kh`Y���ԛ�#�z�զGw�S��ǔ�\��S��ʙS�_����>N�O)=��ٰ|�������S���~��b���d����x��_��n��j	.WO��)��e�g3{��W�����б��:F�1����n�QY�Ӡl�$�@����S�L�f�A�eZ?+A^JVڃ$q)AJd���k���s���~�D됧�76.����C�'[c�-�:���蝏|��o��3w�����B���j�K�q�h��Yߖ=6D�Tees}�FX�Y~2f4�qT=�%Q8����m߮��R�W����w����ܓy�rȮ��ŕ�oJ��m�1��ؤX��z�A�K�9�w�]`@�ߐ<
��WNr����QO~�Qc��$m�F�� ���g� @�j�?B�G~�X(�(�DX�QZ��������5ȥ俅!���^
��g*5�{7 [ ���D� eil�t|c��ز�,P ���|�U���:�A�f�VL�&2b\���JX��]^+��.v�"�3a�H�
����\H��S�c)������sr�g١���!xRI������뭾��R�<ߙ�S��a��|�Q��hA$dʺ�#e�.M(�)�t�u/�T��ƅ�$�J_�K�~�̆b���a��� �T�q�j�&�#��f��d��sC�Cl����Q��É�[���8vh] ��0���������x���Z�i�p@r���� ��~���}����UЀ{E.XX���j�o����%*��<�'�b�h'{��6^�2L7�s�-�I>�ks�N���ԕ��!$ך�������P����g������+R�q�'bNUd�GA�Z�S�����Z����XK�
�۔�
 jv�
2�P?�{< ��3M���i�:n�ˠ:�1~�ϥi��b��"B	%�b���V�,c�L+����>�C��ѡީ���M��k�u��w J���3��EFS�{�^:>_�[`�F߾n^�7���F����^m�}��&MZe��u{=�ג��>;�ں!-�z�K���̸��(ٰC5��yn���OZމ��px��/�6���l777z\9w)[����j�d�g:�qr��Gk�g�����7�}r( �b�M7uj��
���e��*`����^��O��(z����d�yܺ�w�iq���ln3w8�	��EJ!K#�b��I���?�"�oi$�o��P�y����+t��+:ʬ��!mֲV�"E��M�PC�vwC��,�5�e^1�����1�-}�W���*m� A���Q�*�3�t
�0A�K���ȯ�A��(+���c�q�l�d�3g�+E��29��!Z\�_���^K����! �fAj�ZV����ֹ��B��Ģ��@�/�a��}�9���)��?�����B���-�KkL�B���*�Ϻ��jK��H\W��}{GyԐ���WҨ�-�����xkW�1C�E�,���,p�+�	�d��e�ކ��Zpm��HDEa���Χ1Xp��0c����I2�0���$��%7'44�+���0���c�òSZ����)�F�6
�O�Oppp$���G�<$��G-�}�+��wk'�;��^��S�"A���f^[�3"�S�(�؜���B;�����9�K[US6�C桙����[��)-��Կ|��c�߿/�jAh�^�*2FZ�{K3Ņ�
�qC��O2}�P�M���ɻ���U_}��EUFԹ�n+J0�k[}ͦa�����D��r*S'"= �A�?;z?�%X�IZ.93��[q�N��!�!##��sz4寁�d����A�C����ȗ}/�����*�-�h9�ȏ@���1�(P�O�Ʌƺ�~�<夯��kj�}��O���	��X3�ž"N�*:.jo"�{�
@}dԣ��γ���k��ǃd�Vv�{�����hNj�@�**�ߡ�� r7��n�u>���2+8=3#V�.�>��C�����w�Խ����[�o晧5�BK����Y�QV�"V�oVT`�Х�!^N�L�-����ᵅ��b~\���j ���2��m����69�B�����h�p���je��Wu����絶�c�R�˴��{�5?�-{f]�K����&��`>����g���Y��n�.�>VJ+5Swe�*f�:l�m_���l��{R宑������g|5�s�y����6J��x��߅���d<9aI�c�s���v�Un"9FR�
���+J���Y�$;���H��q�	���%�I���je"�<����(�V�7��t#"?�Ϻ�h��_>���%����A����xG;��T��~�y\z֤߳��������
�Ζ��A�*����M����Α������ExÓ��#���p�\쳓.�PM��|�����Ҁ���:��;�mut�T�J�ˋ��z��XA��P8�p����lm���?㋼����6Nf�ֆ"��fyq+4���d�U�Z�3��?�k�h3��)�/Q�mٶW-��=� ��~�:F��a�x(��~��?�(>��rx����N���h��X��f�!�:u�nd�0u��.�V� ]7���ڈtrARZ�^�ꖤD�����^V���jY���Y1'��ֻ/k�����Ć/�WQd�S(��l}�x�v�aT�V�����u�  Z;��x,��Qa�P���wNj�8����\��(�E���!uEiq�� r�1}ʡ�4uG
�4�o*/��kUE�f�BgG����A'�O�y�I����2U(}�L�����`WN��E�Ռ����]��^��3k��>t�k'��5N��)��?����CG��Ӟ�#  @��;�����~_O�����$��@鐢�,k����\�kJ�{��ƍd�b�ʩ��YGI�"棍��;4x����6meϰ�k�ǥ��L8�B0ғ��x���m$r���f�CRO��L�/��]ڶa�.tI�>�=ـ�sW�`y��dh�>	��OEv�W!���,�O��F�%�<��-����D6��JS[�(���&�w<v�ȣi)���
\���ڋ�y1F-���y���ya�f���m�]���^Ց��*�	��a��Ą��J*m���t��`��k!�����4FQ�`������S�'T�$5������� �;�����T�ӵA<n����*�h#�H�X^��ŝ�����A�^.���+����9��o|M\ʊ���w�{��r�U-[�_�~>d<
~DA��P�{p���V��k����xkus�t�KJ���;��iw���� sX�d�@�|Χ�L�-�ӭ]�i^{�:j>I&�X#�?�ı��;�wӡ{=:��}�l\3tWۼ=Ya���0���^0���:5�ao��7��#*�־@���z$�񃼱����I�-~��'nl<�V+�+6��lCM������25x�k���A��0��~!�j����8�+��R�D�|&��^��8���<�4�����_sT�4�aK9�%fUU韢r�3�Yߕ�H�]��;ҥ��n�1J��"9&�"y���pg��o�ի���k$�JLԭp��{'����8L*�ƌ�s3=s�5{9��eT��Q�{��#�ֈ'ȧ(�\JMr��t��YP�$��vg9x�NƔ�kW����5�Q��X�Z�
!q�p(��e��"�#�E�
��>k����A�Q��U���"�*�d�f���L�T���x^�ݭ'�c�:&l��!����.��O$��cm�x2SԋZNW<�+6,|S�Ƣ��#�Ϊ�빘�ځ�*J��ut@ԑO�N�A O{K��J[o��Ԏ��Å�3.���x��b;�֔]%Ҹ�e�'�������:�?6޹��j�a�������I6ƚ~�ҳ��x�p���JGCۧCZ������I�E��!�j/X�'��?��$��)�11!���-�P��r-A�P���j� ��a��A�Z]Y!������0�
5��Ɣs�_b����IH��4]O��R]��Z133:dd��y��	�̷{���\�Gk	��	�vш�Ϩ`W��د�C��d�w�|h��|�[���g=D�mbC��Ka"�P<��`|HP�TO��W8y�Oh���`���~��o'����~�*��/��qp�A ��Y�|"�� �~�58(�̈́��.א&�ߤZ��/%"ɄY����}wx�
����VD#�IE�s����?�%OSk()h��	���#Ä ���G��}BSZzp3=��omL�6�z7��"�*?VaҨI��ѨU�7f��9d;�`���4�aR:�����㭂zz�ZC8�E���΍��M=F>N}znl� rL�>�l�M����:��&H�Ǘ`27�`��<���tm�\+���#�R��YUcV�yi����T�Q���k7��,繟x[?�馲o&
��k��|�M=�.��an�Τ�W���cP-��n���2��䔱��~�ixJ�S:�#\�y;Y���R�O�����A ��y(�o{_��A��b\�
V�&��e��뢕��1u�S�l�6F<�k(9y;g��ڂ�v/��2I��+�g�a�Ä�)�B:�OYS�^*�*1_V�d�4�����R_H����c�w���_ܜ��\�ų%K~�Pw�٘��N;� ���!�sc�:��8��P�k��˗*6@}4Q�0.=PM2𩌉���׺M��e�E����t�߁�ɡ��ڐS�|��M���jfQ�>ku�ݪ6	�G[ڛCŽ��֖E�/5���z�2q2@�*0��l�~А"�cs:������.n6�p��-1jU-�\|�����W�[Ҷ�i��b�_���
�x�8��kv���n��Qd$�"������l�n�;�W���E%�E���w%Ş��6�8��9�rr����㢈��@��}-�3>�&��f��=�~	U�Qe.%�499��t7W���vm�pF[H�Q��e8�m�~���͹A$��^���N����D)i�E�\�Wrȩ���������N���������	�%�=#������ X�PWN�'h�s.�
P?�:�ǣB���i��Tq� ��!S�3�yr	�X�Fr��[����X�jp�á�U)+�U�ͪ����\�VO.��~w��;ӏ֡C�<����©�3�v���f?rgб���a�?_�EXJ�~�����l������ə%��-���>x�����#8b�R�<�Y�q-l"a�75/���r������E�����\^^{��8�l=!��-@�w�����̶0�a�l��d�|N�g8�=��Hy�g؊�H���q���l���j'?��J�7�=AKK�7��|�|�X<���(e���Nt�`�o���&��]1Gt��&�ḔO����s���aG�Ps�����Ws�8?�b����`_ѯ�Pb�;�Gi�����gd�S�SE]ǯ=(�(��Mý���yX�1 6�(��G��>F�������j����F�ʞ���#  ����v�?O��=˿5���}mm�]�ˇf#Q�K��&�
{//�^��ҋ�y@������J�/�EM�׌��8Z%u�
Z�rff����>��
�dˌ:сYy+���]�O�4gȭ�
NL�ȹ".��J����
�ag�~�m����TB���}��̇��y��ZLLԘ���jQTV1ؠ�GW�3��X�-�I!W(��Ē���Z�
�`%�J<[���"LKra�c �
Q.��0d��J���Ϲ���q4����Gʞ�׮w�Q��5|���x�kV�S����5B�S����^��4�-\y��gR��T�d�tS{��,=�w�	g���X����:��N�S#�o�x��Dʻf��l8��i4+����_*EOW�ՠ�E�Q9]ca��� $�DY�VHDg&��ZI�Ƭ�K'�7ViY[��.wnK�QCX;=�����O`�|`�e��	s7VA=%-n</��Wj!T�u/eC����2T٩�c�2F��n�FϢ�qCv5�Df4�i�>��lL�i��|�ӭn�a��J|�N���-�ewG#��9�ؔ�*̭�v�	�Yyʌ��'ZWGFFb���n�?�����7(*�} ��nj�#���#I�o�e.,i
�(:�o�.��+�,��{�M^���m"T ;L�-[���޳���ڎ��[�)���y�����j(�{�r�amN۟�.�s���r��2k@�6��	p�T�^��%���b�D�*�cߡ��5+�����2��!�_[�ê�D�v��B���:y2ݛ�z�lYK��{Wܕ�~������b��d�;X�퍘'ٞD��x8��ius~ޕj۱����ܶ��}�3��i@���~ym'4���+���(U�wUg>3���r:��r��5�h�+������e�ġ1�*�����?�+*t�o�+}V=��L���{��[lzaJ�'kv�^l`L�=eE�_l�N��OQ�T��,8��F�+��a�Ay����-�o<��톋�r=���L�z�-i�b�}�5�p��!���=�y��׶�W�/�H���ޏ�sF,�'��?�+�-�5շc+�{�]���vӉ�91��iw���$�헊B��܋�����;ہ�W�i<@]�/�����55	Y�2��x�X����_㟢*//oB���B ����r��F�l�>yB���^B�� �'��`��-@�^TT֟�B��< �=��>C�B��7+qΨ�5u��T�J���������
cd��/U��Ҏ(�*T�!�^+�n���QW���z��O�"TK���]y+�w���Yo+����,-�����_ӝ'�x��v���[PS�7�oDZ��Ȓ�ouL����c;̈� �L��ZsL��X;� �N	6ka��-99U��냙/obt�gh��Aq/sE5���N��@��{X���3ldr[�e,_��� 7 oG����L�v�����U�!�Fgq,�܄�o}�R�O���&�R޴����?��\;�_]Q�m�����\�ubw��OU�{�9�;��o� ���S��������r@<��exn;�GeXD�F����/�97t���RM2S:\��8w���?��``r(����X>�[�X����T�D����z�-_��
������@����(���ۃ���cş�l촑��X����P��₦*�ɶ�lǆ����癊�𛜮6[L�b#�L	����KQ����S��|nIv�,9r���"-&x�l�+�o��nA�T�ܦ�pC�*K���[��<�>ۚW�ˌ�����݄�=�����aF�j�m�!�bKk�G/��Z*��'ǱZ�p������{����;_��H1��o!�@��z�n�J�֪���[oiS�������ey�GQ��w����7rw4��Ǘk�B�f���dv��WB:��LOXT�������vw�3�D����:��eNNNT��	iymw �p���^��I�WX�ܥ��sn9�2���}��~O���T�(l�[Ĳ�����ޱ9RRE��\g� Hډ�����"~�����TS��.���$����ria��Ϙ�1��@}ծ ]A���)�|�&�m��(_M���d3�x�]X&�{��y(&�5�����qa�y�Y��Ԫ}}��Ԁ��v�XlsT3C}�#W_D���or�ϧ�)�5�Υ�Fd7�$����)�����s:�~m������B]oA�l�� vz�Z-�F*lDʩ�F�������70�0T�A�����so<����H�Z���.A��a#��=�������Ͽ���֒DÁ�_��nd��}�7<��6�Z�8"VH��X��.�x$��Yp���=k�= I�	���^66��w�p`Ć�����~�mچ�3�9�ը?f������M��{P�	_�#��Y����;�O���N�>�g�k@����������������-k�M����XK��mݭm5�q����ANL$��p�D�@rp�髧�����Ew�F@���Qc�I�����ů������n28�m-#bn�����?^����U�u�r��J*Jo�-�����5����ަ�622�5A�`?uM���d  �G��p�+����xu0G�
jON�$@8�'���N^c}��E�J��*�����Ylv(d����e
�?��p���V@���qz����Q�H7���1��$՟��Q�h���2�ݶ���y&:j ,~�>�;��+_ku��l=U�\zZZ�ÞbRj�s�-�p�0\�l��	s�eF�jf2땦�������b5
����x9�}I1����F$ �P�M��6{j�
41�� ��vy��֞���hЉO �/̂,��N$�,�`UT�U�]�	���;OPF�*����JXS�US�bo�Z�-����D@U�k���W��u�M��XI�^�2�g|| `�{��3�ll詼��j�Je�T|�K9�DN,q�eл_p��ns�j"��Y��5���{!|WZS[��;�fT�K�8xێ�q�;��x���� �}F?���(�m�Q^7��o����
�ֿw޶����DDH@8䐯�Ѭ������f붢A������H:��{ad������w9��W������h?�vǚ\T���Ih5TV�Օ@������@����L�6�q�$����='�t��Rp���3Uyu��w�ܣe���Y��[�Ut� ��5�?��^�gE�RAP�S����RTf!�zeT���L/�0��6��{lLhΙ���#����F�o�1�~,�^��]���r��,�/�,S���{ĭ�y���VAy	 ��Lk
��͊F��Dӵ�A��v�jٖ������AF���4]C�L��Po/�2~k�&D�� �f[�	�?�i���k�gEO��u9(r1���ɹ��B�~�Lr�[�zl,&�V�$:�����8�P�;Z�o���RI
� T��|��<Ծ|�  �2Į�8̞ԯ}��Cǯ��e�rc���j��`�z�|��S����:f\
�-:��^�w�� ��!^�Z���PM]���O�2���ݙS��5W�&;H�TTVb(��^�r��7��jDjZ��X/e���V��BǜKK~],P��m/[�hW�� `�����ԳǪ�rr�?yPL�X�~X��W
�?�栓�^���	�_D-A�j9�D.4��j�	Dw�Ф{�U������<zx�l�h��\�Ў�V�b?�S��,�P��UTU}�/�����`e^�����tMw�^��XwW�y�s����eq���b h�Y��:�1Zo�b4�nP���A��n�N����Q"0AH��v��j��-XHY�"x���̒ꪩA����P)��%_���˷��<Ʀ�������D�-��M��EJ�Ԡ^f�%A��~W�]���ϙL�jPrq���Wj5���P����
��k��m�Z]mbU<<�l�M��K�9e#.��Tӿ��9�+@�I��K��Pb�F�?SUm}�y�0�u���J�0z�&��Ҟ�п.ur�ʚ��~�_���9�� �Z3t��_WNR�Yx�܌g�R�ٽ�u���S^p��D�?I���f3\H�k����v}S�~'>�!#�Վ�_H1? �o*��{����歐P��nq��+��!�7A��S��7ǢEpbrM������ �۝>g�aa�v����z)//bb���b�����w��s �V6���;�Ky��g� a``��\9V���m--��҈W;�;��`�񅪐J�/����څ�I0cIy���L�}�nEN��YƏ���~2K�� �����4{��bԨ���e��(��CpĈ2^i$���6XS�U��L�	&����*q�Xrja2�LAmv��N�c��$8��aUy�Ȍ�SgVU�v�Hw#)(! )���%�ݍ������� Hwwl������>��\��k�Zs>���k��/|��ABn�K?-����e<�y�L7e��X$�L���
>��d0���|�f����]\��|ϖ���*�-�����B���u8-�v����>Ax�
x/R��~P�Ma>4_��pI��އʱH��/*)1|���G�u^�{��3���ZW���4���jo����r��ty�:�{��E��K��/�ť��2�3�.�W�l�������2�5��o�ո5�MQ��~\�N�Bg�l�p\����8�s�;�E)!M³�z{3U��� Qm��q���X�Gm��=�n*CJ֋	�)u��ׇ�$���Tn�|K��Tu��.��%��р�eVs�6E��/���l����R�����'(���0��o�ϛ� ��~ �t�ꌋ�UHo����NC9���;#fk�J�fS�ɻ��p��723&�P<�ͷ�"'�]E)
��Șy~�!awJ�~ח-9+޷��$��?$}~V�Ղ��%��K�������I��2�G�j�@��DkY��M�(
��9�A�ki����M��8��2÷?�,��ztx�J�O)ʫ�%(S��Y8M���5��\��>����f�I8��6��:l[l^"�Jm0]�sK5�2��)�W�p�����nja��J����%rZn����yB�zR2rS�u!H[.pA��ssz�޿�\'
��Z�uQ��&k8�;XE�p��~�Vq��7E��u\"��������H��)�2M�8�(/�nqӹ��㐲�m7�"�I��5�������}bk����b����a�mb��3����^`|���k�#��J㿡)&.,b>�7xkF�Q��9!=��7����Z��w�.9`l�}���'�?o��o_�f������Vh$����*P̂��ٳ=��l o��Q��9���%����}^;v�'�g[a�o�Q��Fnϕ��P��!Jy~�Ŧ&P�.O�0��)5y�E�'��<�0�z�Ԝ��P���R�q��&�������֖%9��z�}S�rp�Y� �����5���gC�W� .�τ�x�n�����P(y�մ�G�؟2?AF&3V�}	����c=�VBv���7��[$OH������ѣ{k�%{���.�A�6�I�A=N�;s����ù-��[�Y�o�W�oTͼr�/�<�����_��d���S5w�#����aF���_>؀xh"G�����j�D�L)�V���1�ڦu�q�{�M���.��Tm���sQ�l�]��|����Μː�#�[���k����y�9�::�a�22��-!�
(;SH��� �q�H�#s^�\ԝ�Ր<�F�ԑ��E��"�?���C�	�U��Ъ��܆�.���@�U4�����aUvB򚔩���p4]���r�h�$���t�،4&ķ��ܛ/����CA;]�<�IF����{*'X
;4��s	�W�<��r���&����v7d�
��pS��7����xUuuwG�8�&����b������Q���ؑzȰ������fG��}� jU�O;���O<�w���m��pz89���ɼ���侨����a��r��kA�.K_,L�ݚ��K�{�FI����Ŭ�V�oK�s�g>G�����������?c�ρm|�#�_���A�2�[u7�O���4��ȓ��~����&\��K<|b��K�.<��xᆼ�ֻ)��r:TXȎΕ��.]bG�C�A��2�x�x/I�hq�D4�I�Tt����Ɯ�#_�t@ �!"$|h�?6.#Ȓd����IA��M#�S
~
9��Mm_�H)�l�WW���u�˂� ��倧�ln�P�N�G��
Γ/o�t�~�FGf��Xr�%F���`�-+W!�먵���h]{9�/��l�+����
�\����Y
�g7�y���[�	YMFr�;y��C��zWk���C�i��d�R�]�x�����1E�!m���v�b/Foݼ	!��8l�!�'G���ӵN�a�⪱Q�	"bfYٶ��:��ۦ�z2h��gL*c��sd�7q�[j��(5�'m��%��PxH2_�]��8U����Z�Y��[�>gd��y����P�tj���_�D�۱VL����ȓV��\wu�؄��z�۱�*#��=;c*��z�-��ẳ�0K�^�D����GM���1�����uC���xB�� $�1�Iδ�b�!��!�z���V���`܇|���
�Â����:E*�]�q��b*�ɽ�g�&z7;�'yܞ��%5��U��>pMS1����.[|��*vvvN+��S33�����zӑ����Իw��g[m[���~7F���yF�� 5�ȃG�A�Yۍ� �2萌�
����JFC�b�8+?П�[���" ���_�s��+��5�f=��ښ�eCN|�9"�Q����5A�s���O�>��� ��<�0B����,)�K�6�WjF�v��I�}�VTƜ����BO�#�X�U���{�HQd_�I�J���	�X�7�HbR��ߗ���śPnwU龜���'� �3Z�Q�)uOa#�<�8J��`��2ւ��b��:5���YNI	��ՠ�ra��3>i��9�ǡ��<�O4��H�ʚ0D�|wlfj�h��:#4\�\x��S|���)r�w�(F�P-ŷ����u!�����d�ޫ���%�-ax�<g90�e����Seuu�<����coǽ)vI����=����Z�7R����촒�-\C�_�V�br��PQ��FBd�n_�:G?���e�ƨ�g�?Se�9	��	�v������qWU|cr�w��;>_VV�mg��G�+��2���b�I��Q)?~A�G�C�q֣E��vsL�_N�hS~����7L72޵�������m�g�T^0�r�)Z���CgttteC���!8H�r�~ò�*�jw�l�"�zc�'��ֳ\�������1�rO����A?�2'�-kd���L�Fd�FQ
�fKŚ�>�ifF�NLUS(P��֟)��{m��ՏZ[ ��5�x���T;,bQ���CSI��Á����B���&}�0�-�lY�+55��q��O)���"fD�qjAF�:��}��T"�qt�Ư� )ii��[�O���\�yG؁�t�9�)(��%�=�?��r�Ѹ t�͒,�>	]��s�����́����KY�3&�1�9*>���n��ratT�j�;�_��y�4�1lX"F�K��S�)��/zRRR
��5����Yhg>Eϣ~�@��Q�XX�]*/O��3��=u����97�w��?��v�R6�����$�|������7�Apo<���o��\yN�����(�WJzz���k�G׾U�.���p<B�&\{b����v���d�Cs�$�{�@�ӂg�I���wv��j���qdL�A��񨊏U^'DC�K��~����yw4���~�!<:z�NЭ���,t%:M9͈�͈-���`�`�����rym��;2V�rG�:7SIPt��L�.�\ڲs9����|}����[U�����g�e�I%w�>��N՜����ƨvB� C�W'��#��q��t}"�����^����[��P㠰Y?��urr
�c�%L!��tX���c��������g+���+�iT[�
�w�+w��۠��!�`�b�|s�I��aLi)[Rr~F���L������?�Ҟ5PY�F��17tñ�a��W���5�S�O����Ib'j����W�|6dY��^�����W_������Fzg��f��)�cr^�����Z��A�lž������vhG��	�tLHH���O`II�T����8z~�oYh��O�\y�v�ޙj�|��q9ƃ�3���)b�`"�!��7���`�����jX' ��{�'H�]VV�5���]��Mi�3���׸;ƽ�Q�;�R��YY��)� Z��I��3���`��c@������ld_\ @�?े����8\ȿ�o���-�&)	�y��n���]Ӄ���)��h��j��5 zz���'�s���2�{����]��S&�����q���~���K(`���ck{�F����L�Px�eG���������JE	���s��wHt(�������de{��b��z�_#Sy�c˰�1��Rn��L�*̣���q1�|�_M����B��!b�eJ��B8�ē���#$h/fl�eeU��u7ݵ���6.#ל)�X�����-���{NU[.�N/��|���۟�y?׈W8�	ϑ�c����$ �]7����Og�O���;�w'��ɲJ2��W��Nl��}�-Wߒ��������!w3��}���|���ܝ�4x�2Y{jlS�*v!>��l�0���~�(Udo����ť
SU?�����U�q��^)�3B�,Nd�vR_"��������vp��xU���y�U��:�`�O�'R���^Z�xxΕ����cu�R�v�v�3	�Z)�����-���U;Tc��N'k�$]x^��a3Y���D����3MLE�	|��� ���b��y�S�S�A��M�U)N�dj�+���5�j�>o�/��BM,�z��^a�.m�)<c<ag���C*^�����������jy��r�W�Y2A'H7
qE�����+��o^����>j1��8!����h�謬tE2B̈́�?�&��G/n�ª�G3�����Q���ˎ�F�7�!��gv=we�ð��>%�2�n�B�=~-Egr��૓�ZS������̬���*k�%�n�r���_�x���J�OUX`K�(ǭ*�U╜c�����c-m�����֨��MO���a�D�u���C<�_�v9;���v�/�	�z���6M�SԸl*����<\��չd*�0?6��|D����(F����ɒEx�GL��yy�T329x���X�i��S������/�+1ǌ:��iX[Έ���j�W�m�WG��02����J���%�<nhehKo�6��<��k�}��tN�}mbl��$*����E>ڋ��]��/���:�t`��񐣉@����6	K-Z%%�����c�ݚԙnw���U~������MRZ:G��R�. I�J��Mo�!�aT����)�tq����J��a*W�}����ﮟ�	B0����H�o��KB���g:,6�U�잁7��#��۫BY2u�K'��C��~��5{u� �����md��4��H�[����3�ߍ��8k���<?�nu��܎{�?JI+1�k�#�c����g*��mm⹖� ��?v����>�����>:�ק��(h&@)�Nevt.�>�����J�S�d:�Y]�u;\��qX4�2H��*3����m�g�RQj�/IF�F^r�"��8^jC���b�g��{
Ѝ��Z̩�G�'3U#;�L����|�O��zax6v~��q�8Ɗ+x�7�r/�����LPm�w�|H=~�Yj�\��#z��X\�0���?tY#L�E��['�~������ȫ�����ݦD>��K�Z/}��4Wfü�/�ǐ��|>Z�V�G���=���A����
�8�߿w���M�lsY����WVW�7��G���t��;���F"��?�<�ם��MVp{��`�X�W��inv�M��=��G�8���ٓ��9��Gʅ�`'�6GݣSe{�G��ȭm����ʕS+�P�ec��2a�AAʒ���]�}m�M_��ܑ�A�VT��pu}��I�ċ3V��P��<�u�Ī����o*/��9k�㸿��A��d�Nn����o�ߺ�oEEg�o�����-6��[&���_���9oX&ͬ�ǝ��Z���Z��"l$[�3Ő1�x�5��粘�=�h-5��;W1��~�\G�BR����]���#	������fF���^`���֕o:��S����,�,y68]o��k6�����KZ�&�x��Z�Vl'��G���#�z��B��w�ל��jS��p��;jM���1A���R����3����p���`։�����jBP��/r&���D_|ؒ���3��$/���X7���E蝯�y2�I�_���5�!�MinT�<ȱ	�wjb�$-v���b�+�1X=��9�Ay}d����կ�V�Ƴ�C04�̑���l����^�&Ck>�ЃG�Z�3kB?:e��M�h�RV}nsf��A��O�i�f>�f����>�o���Ѳ��]�L�;7A��p%���rZ*��#sB��+>��E=P>ӂ:�������A��W�y����9��Z���_����ӡ2�{�n�[II�Z'�G�Pm����.���I�1�h�`%��Ŭ8f�:�_8:-��<( �l��Ɠ�л�;�W�5��1k�2��LH�3BF�q@����u���e�F���S<��|��a�
R	�ku����
�ޟ�E��M�:벥%�N(��>jxj*�fџ蟵��!�'F��.T���Ϻs�ҋ/��r���f~(1����u�;��ж.Cdh�ll��Lm�(��9z�|Uđ���~���/��I��8���o��Ӓ��G��.�1����܉�\��.[2��w/�B�Ԩ�9T[�h�~u�9-���Z����7�*�Jtq�9*uIAk�wh�P�
�U��k_&tttYYᡨY~���_�T�������,:ݜYu��211�4�xX��ҹC,;:��#�C/ ��B��`�g�ZٌZ!����ܭ���Q6�\���z���}~��!I�ښ���0��{\��f������>����6���Y���ɟv�o�# ^��{���R�:��H�\�F�+XN���W�C�\h��1���(�%(E!�<NtU>���= ���GWW�Ǉ��ff���+ �&�

��l��,Z[��tњ?wU|a�1�5g4]nv�p{��DYS3��䏼<��M�$����+,:��RG��ð޾{�
[=&��0�%���سV���
��&�ʮ���7.�g� �,�����=�<cf��é*���Il��\����/���<��Ǜ��b}I���4l�,���VEC��5���a��wF���'�ɰK��z͡,�$d<���U�;��r:�n�ˋ���^���E���ʥ&�8�c!�@c����w���B�.D>DVP�6�U�&Vu�k5\|�Uw��144�k�&����`&b5 �s-�%�Y1���������f�ї��>�(e*=$����F�m�����&M�������P����V2����9�<^b/b�����#C�����ǁ���[c?�L�_	I`S
��!��sIBA�D��`=}�TZ^^�O#S���5.���"YQ)2����U�)w$u.́��������M�g�ޞ-��i�J9��f[ouo�-60�?�~��>g\�����s ���˧�@�n<:�Oz,�K�b�7��P�=q��d��/���
���ub�@0�X�|�΂�6�sp�#c��Jд��tz���na%�j�!�,�|���[p齲�y���Y�z_".9y�g�Ύ5	���*%$?�	�A�=��w�/��Z� t-0�շ=9YَY��"�y[��ȗ��A5ag�/�F��4���;�	�T��C��p51����F�?���_�����@�tk�sd���29*��|�R���6�P���e����J@��+�]�U��W77+�9�(((F�	j�]I�&�ۣ��4�2|�
�VŇ`�*vU�'Fߨ�z{����$c�{��455��D()fH�����w�zz����m��^ᗔM\�j8������kocH��Pvk׊��U(	�-��߿I�d���V����ē��G��)�YY+s�=q��?~��N9�()k�5�j]��d����C���6����2'=���ھ��q������.�"	{	�����K`\%�Z;;����P	O�v������-��bM+)[��l	��������.¿���b�ZY싾�����<���`L@��30`���o.�X���k�N��SQ]\\$��uz���+<2���7[��ԕ�˓��c�#�x�hŸ�*,;5{�#Ի��5S�l@%�W��v��H��'�!8�o�
�ϰZ�lG�-�ĬY��,��^Ύ����-��y�JKK��aX���Pa�6�w��j��wƈ�8�w#T�k}ON~�1p��4 ���w�k�����_Z��������\?�K�H��ib�t�@�;E�×��_˭� WgZÿJRA�m����Qܬ\d������Z���*����q��2O��`6������Ϻ+�����v���9HPPPTlMuu7�������Ls$��.7+;�~�	tl���^8��kĝ��r�
@��m�T��頔�];�����_ ������N�0C[�) i����AH9Ynb��a��ϡ�vsK{�����u;�ٛ�<�T�6�s�X:Z�(������WX��	���|��cZt�.�L�Q�(d�.O�
��p��d�� %�j�\XG[���_�+'ڕC��I(᠂{�䋏��g_���#D��@=��a��n���i�+�ځI��O�7M�?++_�mn�����ƫ���Ǉ�;�Š(���_�7�zHkh��3>A}f�t�k���n�?�#�+���3�� :*���j�Y��ı�2|H�{���U��K�qV[�H���v'W���"heD��
��;�nZ�B<�C��C�w��{��B��j���s�o�;�L�K���#)�1]6�`Kj#��fE7��G��	+__,ˣ��L�b�/\�/�~���� Ԡ\���[S����7�/��7�9�����Z�mt!�ҏ��]��3��i��i��Y;^�� �Ù����E#�M��;�p�>�H!=�� $��͂?�P}t�8j��E%��$Lq�3s�Gi��C�	}�0쎞w��2[��F��L��6E@F��E:�fq�й0������d���d�I,����G�Ghl[U�4���ź��ŗ�R�}x\B�Pj񏖍�8�޷?�JOF@쁌Ni5reRԗ���qU������uK)z3//��l{��k��R�d�g��[.��
c|��P��j�{l� ����<&�^�%���g��-�u��:RW'謭��`;��,�	�v-M2G4�܎�nrv0�f�-�Ps�(���o�V��j�{�����Þ�GG�r���!V�*�8K�u��4�O-i�_�2��Pc��K:D��w|��
�
�cѼ���dA����jr������F��΋��w��R���UOI	���T���j-j�b���?+�$�����9��*%%e�џ�����5�Pף��Z���>S)*����\����W�J���be��M ��9-�h�X
�%d�a��ʌ\M|�;�Ǉ<�
"�<��%�u��n�N�8X
������W��$�8�*] �&!d����&Lt|Y��V�wП.DC�ZYnJ�l�pq�0��g�$٨�t0��AyB:���	��,��aV�U�������]��?��͜muἯQ���&��%!��K؝�r��:p�dC;5�?�D#;�A��ZPƆZ0~���PUU�$^y4�-����l�'C�EV]��f,؁m���V}� %���镚@��Ry�Hz��؝V$$��l�e_�ͼ���o>ӱ�e����xNNNn`U����-���������O��2��[R㙎����Of�ҥ�G��+v �yר�C��-��$��l�{�����mmp���8h�����ݹ����ԛ��n	��@�g�w��ʓMMO��̐������-��`�)����x�i�㒨����I��� 4j���q�8:y�m.���X`����M��7n Q�`iѴf6����ice���]Sy:��P��p�hr><��4w3����X0����	#N����BPV%�C��6�6��l��� C��E\�y�n�������O���]�mQǗF��H���t�*%�9N6QA
MA�5ߠh��(Ax���o�8	�9�4�!�1$���O!,�
�v�j�'�4�]?ٽ+��^��8:>(���6��E<:�*,��>\o�S>���b���
d0p��U@��o�LNOOGr�'�:�)��|b�=�3�@��ǔ��p�
UG�#��k]���v��O����֓���)*v{�4�� �W�ڂ�dz�M��|��]|�y��ݛ��"
&&lɘ�'b�ލI��l,рL�_�7ԒR�O��������6+ ���{<;�'���w�z��W��\~m���eK΁��/Z$��}�.�m�6dV6� ����,�(�X��F6�3���;?��V����B��b�j��jIb�1��AP�e�>�,Z�ܷ�U���:���/0z �&j��t�9Б��z3��K����wnL %Z�Fp�k�c_��|p���q���4��eb`��'�c�:�kp��6�XC)�	�U�mlttW ��4���z�r�d���<��@2�f����LNbU��'
::B���Svs��o54�`T����]�u��)�z��O����[��Q$m�V�����?�4�����cL��Ϥ='�BM�u���s��Μ$KX�0e���߶����Y�⿌D��Sm�e'�~S>Gh�� �> �NM-t+o�̄�������r}V��}� 6��&0/�}�d`P<.���5��'���5��pj?M_��t���������Y��q|�X���:���fC?v������t:ם��ŀv����5L��hff�34�5���g,,9������sO��Q��ȓh��w˭����<�3QD�O�o���M�7S�^]]^]��[x7����
x8ͨ�Δ��rtz�q}��xbE)&�w>�i����@�>pvS���zc����֌ I�
.���ta���*YQMxD.�嫂�/q5�+TK���~[JM���������S4���84_�F$��6����N��2���8]$KQ�K6TT�a��� ���Ϝ����v��>!���G�B���̑x�x�T�ß�)rT�u3?��>���KT,Eo�f�29�D7��%nr�u�L�ŝ@j���[�g�v�#����%��׷8����΄ݢ��s�����YMG���ts�i�w�xHHDjiIm�;����͑|||�D��V�[���`@��h�5(*`��W���=�ђ -[
������nI`Q�CC���Ht�)O|n}]���.fJ+*ĥ�Q��P��#���҅��d�p�©A����h�#j�������B��w�T��Υ����� ��WU��|���{E#-�R�À�g�-_�r��Z��W35
��� tb4��v�R1��a�m�d�w�B��'L[�Q�v� J�$�gh���o��������P8���x��j9����Լ��0^�v�3��)�m�p�&�-Ք��k��/>9�����KJji�����*ԩB��=
�8��P�B�������қ�M���X
��.?SMǺ3;(�D�����>�����,-�sT�ӓ���*C/!20��	���G�5��*,
�p���o��w�Ͱ�O������FAEm;�oP֜<�_�p7:^��*7E�-�5�M�A��"@�V���ԝ���ȫ�͜�\#""���O��4�)��� Z��D���&C��N.�����nn��]zl@D�P+S��>H��q��+�}ds�H����\�D�J��EM�|���1w��y��+ �:�͕0*#=������������1&2.m
�'W�W�7�V[A&��2�(Dt��8E������T
[(�Ȏ�K�I,����,?�\�J����:~5h"KM�K�1��Yz7˶�牸�#�����^�A�Ąb���{`�[�����bvv� �^���<6N��^1a*a������Vs��Y-7�B���j<� x4cS���>@7d��B̢dH�.��� �⨇>#�b���7h�¢��&�Is��D�v�V�h�U�R�x�fv��#���������cA0�or�P�_� �)1�`)D��P��srr�C˽ƪ3-Z(�
���B䕱�?6��]yxW!�ǹL���*9���c�Ǧ���.U�F����G���.��q����W)�8JA�@��m � �˴�]�Zgc�$_����-o�cq�*����#l�Կ)=�$ͥ�4���o�m.��h�����:4r��ۛ�˚ ����aI��pN�*Um]�z�q^+	$�/M����`�fx�r^c�'���8Y�A#�|��F)>���?,ְ��q:F�t�C�G!��cTy�cMX�������H�S����4+:�u�n
��� �.����ƯH��Q���5w��{B��	|:��;Z}檟������)aK�T%�	��1 �'4�Alg�1#�Y� �ݬT������b�D�C�~��?lI���^��\dnnN�!#�56V�m&���7j���.�c��RWǗ�������x0��k�C�x>sgWK6N�2�`�����j����p/%,���A�u����'�S�~�G��-_�:>b�{z򊉉7���y_���m�  K���YB]
�{����*WB)2���D{G�H��f�AS��+����_�1T"1 j��Β�+����M֮Ci�E^N<|�	}75;�C�/�r���wh��_�Z�۷ok���xP��{����<M��]imo���$���:�NHE+�@"K9>�Z�ni�`����(��~�tA��ZUc�� �q'JtYxx�̐�F~~>i�&��������Tjq	±Lqd-mm�(��zBl*�£�� �IWwv��o�LX�F�<??��}���B`��M��ԁ^�?�����.�XQ��I_"����k�&�p�|5k�ؙ�X�->>�D%��+��+�� 3ͳg�'E4�EE˫����ۡPd��b �׬'�j�ʸƔ/�m����Ď��k9�KT���f7a`�0������"�+���\�C\��h)=߯ͼ�cc���Kn�i�[y�6O�q0p�!��\����c�r,��@`{r�?ajaa��f'���mll��wwvЀ�¶yh�t'��e���S�"zv�DbQ��,n������}a�}��h��z���,�՝/�
U�3naT���hE���'kĖ������anoo_ZZ:�3�s������o�~�{�0Q?��
��cl�����c�?Y�~��O�.�\6� .��1������W'R����d�w���Ag��\����
s�(��ҥ�Yb��&���2�o^:��0���x������d�%(�N.)$5o��:|||�� �K6��� ��t��PF�KN���*b <8$$^�j��d<ݿ�`��S�p����joYmO�R��ov8�A�������R�;��i��lmUYR�:%���5����]&'�8\?���3E֦�!��TC���46a)�S(k���V10����$�pBL�!��N�X���Nl�ݟO�9�Jz��tLNI�ʎ��E�ۖ���2�er�����I�EK7�cf�\#����:
)��������EzF���;ey�˗��0��/rL��Ԧ�y�,-���o�B_���SN���$v�Jg�=���`�h��3�g�}��X)�-Z��6�Y?�Hnl��azI#��0�W���-�$7���c*�i䇨�DWߦ�H�8���>2ccc�h9:�s`LÆ�1�h
t�8��d	���_E����l�l��]&777  ?_�\�4��n���*��ģ9�L�x��_+��p��1`���}��\D���>uE�>�k2��i�{g�UX;hlo�	S��yTZ��;&��i`����4�/ʳa��y�����]�lkk{��+�&��w��;�j۠�0)7�$���Lí��CD�K��}�q�Ș\�YYm��a�fmmo�ԧ��If��{��I.-� �6,�q��h��՛�JF�@��ϣ����dܶ�
i���8(��������L�z�,�({�)=C7]\]	�����T���.�~��Kw888�ꆄA��=���ϵ���t�U����t�����Zv.vD�����FOutt>a_�bP
j�n�����E�ǏSI,�,I����um�@��Ⱦ$99��� ��J�d���{}s���
�N��=��|(�-���|�ݟ��h����������z�'Aɽp��i��15}����(sj3�����X���H:1����H��s횱�aѿ%��I�'Y��_�T�Li��1����
�3lIg���ʥ*F��E����	�ʸ�Z^v�5��K��4��5�$/�u�'�{+��@�hE�>EE��%���(wppCG@@8��u� 17��&����[��څ/w��^8())�n�6z��
kjNr|P�	[1�K����r�`�$�����5 �O�0@�*X��k�X�g��ҥA#K�J}G�g�%��T�x�3���^e�6k�$�7/hi�=T[ʚ��j5�mM�d�v�6i��)��M������Pc�?:?'�$}���G6�I����j?$�Ý�軳�E�Eou���!8YyyҩB>�I��S33��Ρ��͞ _v���������������XN�f���붷��vvuY�m�5M�loG��1D�eee��j�W�@B�����sT^z�m)o�yS�`Hv�.$�T�uw:���>~�����55u�!��S��0� �+�<�����sCO�����my�ޛ�<�(1d������Fr�L�'���z��������"�p���-,,�k�]!�����@��<�g�������vc��
F�?C�!b�
�D�k�ҍ���7�+@��[�P����G XM�4qK������im}�����	��M=Cm�G�\��f�Ld�s�ʫ+�2p�#5�~T��0�444�5;��iT��;�Ғ�M �W��wҍ����v^:�9����
�}�no��o��@�D��&�����v�n+pٷ&�4�����>ЛF�j��Ϗ�W��(H�o��>þf	��o~Tj���ނ�麻>}ki����\X��u�!�j2}��.�����KP=^�Y�6�㳀E�#z�p�����ɀ볽�PY������ɑ�ك��g��̵�$3���sp��$������յ�sZ�s�*q�����ٸU��AH@.�x�ڟ&�	��A�gVQ�l$W���j�E�2F>�|Нe���;3�V�HF�́mH;��f��>�����[YY�����/Gww������XⷑD�:�k�l ���X��Mn5���TO9D�X���v�;���0�t�	Q���#�]]���Y[Z۰?��AI~��JK|r)��U�#S�4͝��z~�����[�d�c�L�c�XY�:);7��$0���Ҟ#��izzp)f�a��_p����_�p���?��t|,��f���)���i}�*ێ/���3ȉ�C�/~�(�������qX$-�FƠ���������^�`n9]���������a4
�z�=M�l�f֗m�0M:����K��n�e�}�9B�е�
�Ú^б���|CK�v'^-��2�ٯr�����q�����ؙ��fmMU���L��"��j	 ����~�_��d}f5`?�"��;S�l:m�X�d��.()��)C��!˂ϡP��
��.��mCCCi�+��e.�9:�����0~��@T��JI������v�ֻnE'6�����u�X���� �~�{��),N�v�tvJ���'���g)//��Ƙ�����8��װ�@@ dcc����{ikEWW��D-��P�T,l�v'��/i���iZ���̟��wG�wG�f:+��"Ю���Lq��2�O�>��◐�h��/�l>���ɾџ���]�mlc�;lk"l3s�%�:n�5�Ѱ;�`�Oa�6Ufª���V����%!A�x."򌟟�es04##��
��1�U��LRB��(L����a�h�a����@aPA� �h�/#�y	���+zAGG��&�<mmmH`�<���%T�|RJ
���.7B222-]ݎ�n��� �~�z���\6 
?��P9p5�D\2��j�>����'�n�s�k�s���]��
�ۉ2��݄��3����y��#��o�y�������l��eI��I�ۢ�lk�L�p8$ ��u�O�����fm�RUU���T� ���~Hq�#��CB,*a溌�<	7	R@ޢfHA����;��;2�=��������r��ګ���J�VQ�;g�eeep�!������$%1xȸ�g<Dd���R,p�����s/ǽ �%F��r��+�ʋ��K��D����W�cy����2[��v���iT5$���B�Nt����F���+��u���7��Կ�����2�t���0���w�f�A�	}V�,JP��/�n&� ���]��qq{���P�y�fk8C���e��/5�N(tT݇�&!�A����T#� zpw,.�jhDs%l�&�\���r�u���#�^.QD��`��J�x`"O�<�J����E����<��j8A��uvf0Ga}wuL*B%�M FQgH�L�Vi��N�K�7B\!V::$888�æ����y���#Y�[Ӆ|����'�@Fߛ���싅�h��WV��9�P�&�m*����lM	�Sp�yy(@:a��]� TTT@ ��4�R�w �ϰ� *`�M�1����@	�������c�)�!^S��~�9wG5��ZW�Yxrz
22�k�W:������-�:\	8��߿R,^a>����1<�n,K�	����ou&W`�}�wB��g���]���QP`�����z�:3)�Oli���
v�1@`�_&�s(��<<����<hM�G�4K��\�ޮ-w���������{��p}drʹ<������7E�[���"��T��bC� ��P�H��M ��?i�^B@�����Ђ��o�/�n�wa�Sc�ILL&��N�4���n�w����xץ�t�ǡA�Z�< �r�,��		.q����M>& �i)�@�OU�un���^�ߝ(��=�y<��ǿc߆B�dKHeO�2�ڵ6֐���KDF����%���VB�De��Ȓm,���"[���{����̼��|�<�yޟ�<�d����lu��Fo�=a jѺ u899ͷ$��1����i����)�I����7����/-�ѳ��ًg�|�S��p��h"�ј�R�R���'�qsT }�������՛�*�d����{�Ƕ�ݢ�Q���Q��������F־PF�����y�)Z�W��:[kL��l���H�P^^��3�����˛�}��Ͼ�����N:�D^�u�1ۗ�b{mL��Ii��iyX �������Ht��ӛ�.I���YgF�A�:et�fv��|�_�5a+��QhW����S�9|;�Ọ�m��/#p�{}GI��'?�okll��Q�w�|jR�1��o�p��B���z�j���8����m�$��::��ɨk7i�A����1��Z[�(v��S��P��7aS�k�c�I�nn���@Һ�����&�����.|�	�D��Ykk{�a��|||�`'�q�178��cE��w�w�fRa��j��n/^��lPW;߿���k��} 6SV�a�	ֻ�S����\��d/���1z�� 8])))b1Y�"dn���R�s��������%-��<0�9F}�|��P��#L�Z
;7wy�:��@�K����3\�{sB��>I���*��@�c�kx�p|�`C�ה�`m���ud��xy����di����C�qϰ��;�s�n�H�+�h��w�E4}��ВS^ϼ���{٭�t��՚��-��I��_������5|�!�u����ؤu_���H�������Dmkk���PJ�@��'Ԋ��k���������#e8s	��Ѫ���g.J"�Ɯk-:��:2���ʊC4@=���uh�}����&�m���v&���G�>�E�r#
F�|Q}��$�������h%AZ���ks_��us�)�ߝn]�
7>pVI�@`RU��/Z�� �Tc�������okee���C��۫�qw�}v����6�E�0��=�fj��Y�O4~�yAŸ��������<��={F�kh���<��ѓ'%M��G��1a߾��\]]].�RT?	�y��j��NA�
��z�	X3��(#��RS�A�C�9R�M5�X�yD����Da����ٟ`4��#F����س���{�;YYYA��Wx���������`u��8����gr�QJ��򟜙�a����𖖑a�P5F���K��k�꭭� *��ع0^���x�MU��k5�uv0hXi#���M�fj��I����I�E&Ѡb�����gQ��lhqe)�%!��A'I[Ql+aU�#X���qx��N	�Z�0 qT
0�K�5J������ --�-��ܹ]��+�GW���Cx��(1X��+7=���G��H�iF<��5@IY��J ���T�%��;{{�Լ�DM��"
e���Ԟ�������UW�ci�'NHhii��)BGg�P��W��~~*�733D! R�_�=��t#-�v|�R��VT'�<���qq.�	��@�^���.�&ߋّwn���ʊ�#t�#�1.T���5����)���u�F�U֣��N�����߅Ls��tUUU��v�8 ��B?�c�aK��;��?N��QE����L��s9Ck�K�F��'*&���ѭ��ؚ����O[9�T>|H���OH8y��������5��6�"��:�����@w��8�Bq���*XԌm����Smu��y�陻�}�^�>�=��j��sDu9	�J��o߾���w��>��+��)0T�5�r���.����	�����ݜ=���J�Z����c��;G��d���?G�T^C�F��*���OBO�w��AC^m)n!����[~��g�Jd
�4��~�u�z8����6S����׾pxy����Un�R������FdKP������g�(؞�������]��@��|Q�f�=���-���S�[�Y��l���	包m�w0[�ՀT=p�|N�J�H
5��t�R��:T�,$d1	l[���M
�>r�I�{�LYVN�����9@x�;)���(E��85�W�[�[�ʠ�م�8�D�3��*S_����M�Ϟ���ϲ�~~~�ȕʛ����ii�����E>�X�_�ZAAA�	��7�Ʃ�fS���nWW��g��SjMlו'�j�.��8��y)/�)��H[��`�������6�3E��������o��R-W��o^�o�8���^������`�M������$,Zvvv��+`����5�C��RE�7��r¬O��LMM���xp�	�YY�@;z������b�Etu�����_�����.-UDw��-����CE��]��;�4D̒��3J��IT�������K?�9m����Ua�"�dqu[���R���Ǻ��}����+��W_�CU�e<�z��D�1�|�]����ϑ������>8<�Z�� �[[��˷������L�)l���S��):�P�!�[Tds�^�\/��(.>Փ��]b��H�j^��Z|9�2��T�|���g�a(P��e{��#,��]aC1ű�PM��nWp�.�[�Č����Ma�W�LM9Y��ˣ�H��\Gy8 X�T� Q<l��i��n�O���.���������>�k�㥤J6����OD�2s��G	Ǆ9������ A�r�a��0��� 3�x+iDd0Q����h�Q'�[�D����� SS�а����f�kJ-�dedF�k��?<��O\�)Okaa�fA"�O��~!Y�D"��#$�:(��7��١8����Ail{(A��zZ���j��_�^]IMM�;�pSڠ����5r�g+��*�]�*JE�q�C�~8u�������s<��AQZ�)�/2�ا��bhH��l��H.S� ���TTT��;7�W��j�aqtcx\'P��G� r�e9�l���^~��f��;�&o��WX�o�0IMK��c��3����T�В�3��Z_�y ���-A��=��8U+3�q�6y*8�Z�6��Y��*D��&%oD�4�fNJ��z>�BV~3"`��B��na���moߦ��A B�ׯ������o��������Ҩ�%a��#�X���;2��)yU,��qX������d�2w���r;��N�de��q�nX���(���I0[`� /f6 ý����i�����C�LN��&���~�8������l�S�ϛ&��y�nVJ\^�!�}�:>H!qہf|�{D��;�4��f0R[&g�v�NO'��@��Y����J�k��������J�)fL���w���[���<v�st�\|ϥ%�Z�)W�+j)�I-YS��]Z�n��;�v���edU_�u�ðu��5pf��p��`��4�(�l��-�ӭ!pΑ��/J��H`�L����i
��fq>\�z^�Pd�/Q�\!�z3Mr�-_2��"�6�#"�N��,p�q�V��D9��ü�nl� ����������Y�3_:ɋ�!�O��1�6���rH��ن�����˔2c��@U.ﶪ|>��z�R~�&���V���T��3u�h?�[ʎ1,�M?W<k�S��,2���*fmv�q�¯����ָI^�O�8Wb���@R����C�){�L�9/�2�tc���Js��>�h��_�5ă�]4#=SR���� PK   �X�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   ���X̜l�T~ �} /   images/9a4dac29-fc17-4e8f-bf63-f97779143c33.png @翉PNG

   IHDR  y  �   _�]   gAMA  ���a   	pHYs  �  ��+  ��IDATx���i�$�q&�q�utWs5q �Œ�5�(��X��e�>H_e��L&횉�%�K� A3LO�u�w�����̬��:�c5U]���{�?���{��ٳV�s�q|��eY�ԍ4m���}��j6?�L&���H�^����$�ܲ��ldv�����o-�}���g�k�V�0�~�/�~_�(�o/}v�z��qm�H�4�\EQH�Z�w^!��Ϲ4޶� �2e:�b��7�?������jW����I��ZB��|7������Ja��u��gߝO���g�x���}[s�Q�4>~f�=SV�ԭ��J��۷���K%�Z�n|҆�ھ��آ0¸�sn[-�^�3�G�|��������_�+��I`�{��Zw�v�[Wv�{�^��{`�y���l��J�TϤ����W�s���*��8#|������ޚ��-Ʒ�t��y�K��Q���a��L��-�gs�g��M�d#+������}[m��:�
qV=_>���G=���m����!7����?x"���Uyʋ�;;Q\�<'�����S�=� ϴ][�Z������5T����z���}*Ⱦ��+�N�sxp���O��K����po��s���k�Y�l���Ɲ'�-�~���k��o�2����z,�2Y�W�����;yq,�a�5�tO	��/?:�n���+��Yú�oT���h�ֿ9�1����+���b&��z.��?�����?��x�����������Iqp��ol��}fp��k�W�y�72�۳�V�zr��4�w�~��j����m}d�uu���f�g��������co�K�:\���h���~5���y��Q��BnF.>� A�G�����McJA�Y.k�!��~�Q ���Q��R��䅇�ER6�$QhC潨��o�'�$C �e����w��릱��Ao};����U	�E���{��t7e:</�N �n3�m�@��R⹼���{se�U �*X{Á}��d�3!K�%���P�xz�6��G�ےB��)���bs�M���dx��y�`�@5��{c�
�)��?P�[���x8���^���q���ëMh�%��� �
|�w�G���������%���N�{vHo�w��3���u��� ���k�m؝��>�);�����#(����;�O ��{��h��=����r�plܦ��*toQ,��[& c���dJΔǧ
�;��[S�;��"���r�q>"���ٹq��=<�0�3�c9� j�֗���@������l�h {�M��u�\w��<=�U�d�3�y����]��@��4�īi
<� |�X�Cp��WN��L����6u��u�Ga��lY�[��������ˠ�Sp�������g�F������}��:��� ����b!i�^{�|���Όm�9�5�vYez߲(����:?
d��m�dp�sZ8O��ǘ�����Qs�}�tM���\�>G �|m��U�&<�8|�
��"I�9'�ǒ�#Sr�r%	��Z~��a�}���7�3�q>e�۳���n*4���itӀ��-�jݾ�v�N��=���kB���-����lwd$��`➅6��̜�h{�A������"�x�8�>��������*[KNgu-�4�Ab{%��0'��F1�/��C��I��s�R����*X��w����3��3a피N
n@�7T�oʁ��������$=L16�
����a�m$q� (�!�#�����]φ�T%��6f!�,��Y�@�>��|�z̋T'u�a�⍅u���W����^���m�|z�v�V�~��t_���k��a�gQ������~��}|_�6�;�(qرX\�߻�ҽzq���9j�zN1?i�S!V��s�:aƯ�*�p��N@O�Y�"�||�e�@�]�J���PYqOe6wb��og�o���k�GP��2�wQXp��k�N��C��v�y���#]c��:?�j�P�=���Y❣��t뵸�=l?	�(�#=g�x�벇�Wc���z����C?ۙ���|'���R��'�*P�O�kG0��	΍<���>�y�v66r �.PCb�:U����Ջ��i��[e咂M[�����2�u^�z���v�b��\��sM�4w<H�I��w�uH%�Q��B6�3C���}5����t,�,t 4�
A�tYX�W�sH Sԥ;7���# �.�B���ӿۜSA�.��y���Y�4\/Y>q�&j���.R CpNEڝ~�V+��P�����������?���<�|�_����7�6�1S&E��QNP9��b.�,�����:�d0����C�Ι0����%�E i4^��|���[�+)�N�8d�e �9�awR �\g���'�u����"hY-��PA����U�Q��ԁ�ε���:Q�́\�0ߪ�𻠋*5��H�aM )�߰�I����E���Fu�99j5b;�Q��z�5��d4�5�	���m_���r}�`�+�'�9�a-t������0¨�8Y��Ɓ^�|����c ���[�ҔЋ�c,��2~�)t���]AÆq�d+�� ��h��J2�4]���z�i��#3;�P ć��oZ��=8<�s?N�����6l¯�B�6EI �iX�B�]�� 	�5�7�X#��N�s�s�"��CoZTt�s
z�M�@�g M�N�o^{)��`�2��o�c���" LSMc��}���W��Z�Th16Tϓc�F��<��.�"tU�	���W2�a��jm���`,�ʵ��l��9���5|��n���98���y7{�}5���3|v�	�-��MXC���\w�����]�'�K�M�j:ݗ$��V����p��^����{��z]��s��[� ��1����s�q�<p}��/�}�/(
�v��z��Q!����0z�WP�����<c����U4�Pp�ٺP��w�u\*<1]�ڿ�q�1(�l-�:��6��#p�JA@����uW?I���}��p��C�P��FW��fǉz�*�PNkX����p>�^�`�r�d�����<��Ae���j@~��'��z���r`�
���v�Y����Mg2���	��=R������H��x_�&�c��T*�������s��
�面�P��*+9/��4�8���Y�yO�zQ ��Lu��:�g^��*�����j�[c^?�w<� ��|�Ե�/���Mz���XA���:#�_
��|�S
}�����M~����>�g� Z�����t���L�cO����*c4�]]���Zh{����ӧ_����uѐw/Q�!�
G{� .I���'�k�X��v��Q8��.�b�-�Ξ.lT݂�p���$����B�߈�{i�y�������@��:���:��\b�7�X���J��H�@u����ʸȻ�l���Bkq$��N]+�b:��֒,��PY�<��D����FJ����M�(�nl��w�c��aP5c\�|���;^G'Ye,��{�H�'�|z ���|26�Օ+T��aȾ*ܝH0��ie,�s��J|hg�Y{��C�9�B)��X=5= P/���}�b���)iC�)�� ����aP��>yը��S�%�5 �`9�;%�Y�Qu��t �w���ps0�Mr�iR�E�)���+�z}*e�9�}�����
q�5�����)*8P�wP�;�@�k��y�=�boO�чs�t�P�>�}~,a���ʤ|�ZB���cWWj��]��`��F�%Dn�2� � ���a��SLD�A �ʊ����)�����+���0���j(��y�kg��w!�w���(&(#��i�{ ��wp��tSB�+�z�n�	�*D�G8���c�}���S�����
F}o�)��4�o�#���bl%�&��umU�a=
)���O���qO���Zf��r�򥤋���X�^�ֳ�=a��"�?�tF�h�^�X&��e|����S�1�z OP���vv���o�ID����\CN�3r��س/����)�s�n8�e"��=�並�H���X�_,d%�7�������WI�'��y�!f���@�g�T�h,p��H�X��'r)%c[�9��A�k�@4e�� �{W��F����5\���a�5����,��G���l*ЫZU��r��z�`�߫�!du(
p��E�B��+�z�x��g�0��:ŀ�0Jh��<����&ċ@O�vǽs�ˡc
��ۧ-�@����^ 
�0O4/R����I �Y-�'���gmJ��c\x
�%�<w�|A����ʑ�u!�2v��?OuRkku@��:�ֹ �M�JG� PZ��ޓ��$�y�������	��c�N6�ƃH��kN�r��I��d�}O�<<�h,�+2Ԍ9;>�:��͹\<;6��1Wt��/�d,�A"�u���Z�e�A��L�߾��'��ଓCo�. ��M"���%��ń^�N\y�F������5ڔ�Y\
��;l�_ |��-�!��|�؄:����p�M�v����t��.4��!S�:���}��w�y4��O_(�q���}H�$���I3@;����V6$�@q����\�x>�x�7���������+�������kZ<t�MS>�/����}X]�7R|�Jl�1,���X�^Krz`3'��;�'��G� ֊�Ћ�a��"�Z]�q �c�=�p��Pژ�ׯ^�b�G t�,��;�/��*�.� �H�6� 79i� ���,��Wk���񻺴�=���u��1�N�5�����kt�<Od0��h<U@�P�����=X�kY�+�1�kh���(j��	F��?� �ݠ�;%9�m��� ���Z^�x!�ݗGO��k��/�Y������X�jX.=rj�Y�� ���`�"�UA��%��T�я�3���.L�<�#{}.����������}ك���_�	ð��̻*Frׄ��x(�!�3����y��U�y���?�Jq���$WÂ� ',�xk����y�W��<�p@_��y����z���=��b=��al # L��D��!,�V�e*+��
�G�g�?J�nQ��Xa	zɵ�.��I��aʯ�ￗ���x�S�p���,K�W�/R`�i�d٤*�F�D���ȵ���Ƥ'�����R���w��,�l����]w*S�&hby�_������!~]a�^�.`�*����:h�qu�����x��� �Xo�����/*F��ڃ�p��Y��_Z�0Kd��ϥ>y%ɐF[�ʂ(���7�J %��U�-zx�]YT��g?�<����;?�9bKa��x��o��)�R�ofr���d���:�{ 1 ̘�B�,|;��/3Y�c���D�@&���� �rq�OԃU� &^�:#Gg��O�ټ>
���ٙ)2ry�k
C0�1���fX���x�DF�O�\ȋ5�U(� w?���;�to(�R��ֈ�<z]��&�~�<�WU=?}9���|Hb�S|�WC̫���W�k��PFG{2��~�LO_��^@)f8�d�4�=9�I��'�8�Cz}(ߝg�K\R�#\�sGj�G�!�V~��I�X�!�{�E�Q"�U�����J�_?-�� �KY}���Ԑ��ײ,��/<w0�q=��'��u���8��_t ����S����L�d��Ȫ�V����ޟ�DZ���X��P�`
�z���H!'�)�n赃�:2��Sz� n��������1���D��Z����y�5��}����6�y�S����Um^v��Im�0�}��³>�3���h8�����7D��n��t,��!Z���E�d�Ӻ�I".Ҥ��H�t�" ��	z�k���l��g/�)�.#�/R��d?Wc.�F
G�u��fH+����Q��@ |S��x-�x4��q+���Fc��?i'� �{�E?t}q!�_}-˿��O�����3� �̣\���Odż>I���@ !$���L`Hd�CA)6�3 �Zo`�t���d8�hY�<]Ih[-n;�yK�nd�ȠHbzYp����3�^�b�
�X�A(y��	b�-L+�nc<@̈́
 ��ê jf,�J��j�D�1��
�:�������޼R!ȍ��K������Grr�4⹡����AQb<�G�J./��_'/�߿�p�����㗧�:9��Y.R���?��G��f0�:�8FR���x�B *d�p� ��xԟH���C�G�8�Ӑv��������r��[������*��D�HH�m�N���ݻ%�kbL��_��JP`�{�Wd���g2�'je�7x�H�@	<4<왳�Z��O��� @2��>���u��R&�L$��Y�Sc�&9k^��\Bx���a�/`�������ُ%"��"�K^t�P7��)���˧�����9��|�IB��Nad����@;�פ�h"�`"���̖׌�`�`�ihD����L⃑<� n<�׍��9@�tp %³������S��z��TP�P����+�s��n�!ϼh6!n���=�cm���K��f��O�w���K(��K���� �U�0)����A�C�)i
2=f� YmJS�M�����X�O~��*ɽɝ<f*��(������0�r�Ȥ�2��"5|�\`N*(�W��q���0h�����f(�~�s)�-�lȧ
�<f��3������������$ ���i1?ʓȳ��U�E���'2cX�ܤ��m�#�����e�Ɂm)�GNu͝D�ZǱ���L�s3_�o1��~�RuNKc*�C�zK�%ù�^��������9��WO�:���\+,`2`g�7~ �����P�Qx������xvr&���Frȍ>֧j�_�r����?��\@n�\ �c훙�'s9�a0�J����|����@����۽hHib
ޛ���\��?ɃƗ|�p:�','����<���@a��^/��\j���\��
��фے�v@���c���A>�s�3����Bܾ󬆾��)M=��s>Y���v��2u�c�5|��jȹ0�������.�f��Τ���M=����ό�U�a@0��o�g��%+z�
ˤ&��hj���ŕIi�1Q$`��U�>��1�R�Ѱ��^���#%�k��b��L��z���[ �3�-���A��;���<�wX�P���?��^)lf�P�� /q#�$  �b�e��C[�7S&��a����c�a" ����f��dlB�<�������]���5��q�4[%�1>��J&���ߢ`R�>=5�&��U�ʇ�&�r)��(��� �龺s`=���Z�9&u�ɤ �kUD{G�����
 �`,	�e����2�3�?}"���';�$8�ǃ=�J\�g|��j�R�3��'�P���%�B1A�D�{%}���B��߇���)'KY��+jI�=�ؤ��O��k��&��r��
�r����#ٟ`�*���|����Q��~-��D���?)��(堹C9����'��܉��#Y��5<� ]6��"� ���ci�o$}����U�����ٳgz���]y������#I�O�م����2�j��3 �/�Υ~| KXp=������bebh����|��3y�3�d�;8�#�{���շ�7rA�:���~��P�S�ۿ�[ �T~��'r0����+�7��rᾶ�-%Cp�F729�р�e�8����O�{?�����:�"�z�f�z:Up�p^JޖZվz {�%�\@�6�>bv�`����p�#��yu���>��Ɯ3�iBNx*|i�Vb!}z��xJTx9J�p����:W�ۃ�'K<K�^��%i����CH�e�� 	;������3ǑP�ɴ�����z�B�Ʃ����K I8���Z�hԑyN�"=h��c2dZ������T⦐�1�B�KԣE�H��<d��@^\I��l���	�:��ˋ:���a-,����u`�y>#5T:J4�#�����XF�`��C�k�'f�+�8ad� 0��2ƹ�V2�������+H^��i�Yѓ�� �~xN�7;!���!���t����txvBN�JO����� }�ۧr c�>�v��S��@�]�4�֯`HB��LC�ݕ��&&�`����X�?�\�c/]��y>���X�Y|��@��`��Q�!�p0��x�z-�8u[�9���>u)}qn�t]W�V ��~��i��z�|��[�m3l���q�d����ϒ8�'�ݐ���\s�ݪ��\h���S`�)�O�kk4/RO41{�<�D�7�o�~__E�IUܛz�aV+7�j����IǑ�"�rBr�yOr1��y+K�ʌ��w�$`��9�m��z�Կ�	n�o
�������pO�мzq,��� ��c������ ����+��w���%Y�,k�"��L���=J/��BI/�W�Z���B�v5S���dJxTY�<*��w^8ա$���x���WX�$'���鱀u�;2=����#D��O�j	!�Y(��X,% �"M��x.�Ά�	����e�� ��r!>���x��`�HP�K�Ć����3�s1�"(F����2���&v�C/ �'���䇞��WX�1��

9��?��q�ܓjГ�h�yø�y����S%y2�
�ϛ #>��������ѽ�x0���|�@)�Y |�˕T /�ӡ܃2��|�|E�r� �I����4F�*W2k�͋��� k������6�)`�z)��@_���k����j��u�/�o��3���Gr�'?�����{\��d�=�n��kh�ao x<ʰ^PV����PV2�.P�{I �P��O r��`� A��?�1���!�9��:�*}�4��Y;���Ut�d��
��e*?x��ׂC��:W����#�8[,4k�@����%`
�ʓ�"����b��\�$M��(5y�������	��DKc�]KU���Z�����D��.��g� c�w ��TN �	~�H#���}�}]M�ۏk������?�����3���k(�8t]ݛ�I�O ^�#kvN�PR%�SI��~ϒ0�<ޓF��V�|VA#��Mb����'ʱ��kI.5<�Y���Ki��� b��K`A3qq����#�=��;���d�t��[+<A��]T ͨg2U���΃���	����Cy�P��'�[�:��Si� �P�_�+�9=Y7ҫ�l ����3�(��V=_NV	�3��� ����7��!��S��|��NWx?CǞ�G���@�I�5�S���HoUɸ��,�E�¶�Y�|��2@)�Z}�8�3�vD�u�z�d�3�h�/�Ǎ<�3*U�W�^�ų�0Z��q�a���B'- N�a%����ǒՕ+	C:&��~dV�^�d��n����Z��uUԨ�yv��цڀ���=�i��Zå;e�U��-��P��[-��Z(cp���;k�̐UZٖ�a�X�^gYE���D-{�y݌���e�@#5�I�a���#�CM�|z�bi��7�h!`�E&����	w@��7�R�+�%���W-�f���re���X)�3�AR�1�|1����Z;�Yn�}�ʱ�kI��EW59ga�fe�
��1�S/1�YῊ2���a B"�!Cx���˺:$�1�:m���l�ذL�m�-���"'y|ĉn�z�I�� �Z� ����҈Zߕy�����!5��h�h�=(�l`a�2����0�4T�}�s��[�����E�	v������ ј�d��� �7�p??`�e<�C�������ЅN��\�N�O?�)-��7��&�2\��%xu%��u�0�~s�=r���q���ϳ!&��}u�fqQH�J��3(�����A�ͥ�q�ܭU�3���_�1 ܣ���sY�|�JMH*Ǿ��0�z%�W����E��&n�7�f�c��(���������� @t���cy�eu�RW�˼��֣Ǣy�Z��F���Z��az\���d`��d-G z��_~�=|��EZV'{}���Slhf�K�<��^��Ȫ����r�7� ы�0�,+yc}{��g�B�7����q2}#[��H��.�2;��'�g�&���D��� "��z�� �Gd'���I>'Y�8Ƕ�*0�����9�94o�����~���1#q�{�����.��%^hi-x��=�j�=*� �
S���b�@@x6�3L��X]���$e�7bIRȱ����Ld��\��g���Q\Ô�����N��D���R�8����A(V�7a�
�� 3��Fz�r6���Yǎg��+��!�cd��1����%�(�x�\%f�n2ra�7��� �zx
#+����\�Mh��vIpx�c��N�BV~��v*Rz?G��-� �9y�����]��7?���<H��;��_,%��5�)�	@�W�do_N�Υ���3iazE��f�s���q�^$��@������T�{�Ӄ�r�����9�������B����/_'0 Ɖz���i�V�|�#�s��Rr:4&S�Wv� ��Њ
���cdI��V��0ty�Z��6%��lj��ٶz;����i����J�X) �
CC�i��~�����Aq`�#`rM[o
k3DJo��Ы���������+����BU���K����[7��=��B2o29w����TV�My�4���Τ��V}�Ȕ�~��V# ��F>6�D'�Y���T���d�5,�������TJX��P�f��m��7U�İ��wZ�W!��x�ׂmd��0-éR��A��d��2d1�;��JҦ����Y��R�m��5Ǔ��x[�����������Gm��0�p�h�C���^��*i�ue�[߹�K{&�n�)�����v���ar��k�?�A���\vq!��� ����/�A�2�>��a��^���@U!�Wq��fg�O�'�-�\���)|v��#���K�8�,�l�)�(��LS)�s�LIW���K�ή�����ͭ��%*���EM�z%잁F�~�g���ǥ�%t9y,)�b�֘
+�"�Q)�bɴ�X���@�c����e�����yj��@�����!�#k���
l����Ӊlfk�/�Q��P�ept_���7gjd�{�,�r	���h���]x�𐯵ZU ���2��b�		x�z)��i�bo5�:k2�5}ء�j��8��J3N��
����ЩП�z%ɳ�8���K|�P�ғ�R�&��c�;>)�< �L��C(��T^��%=8�`o {���U��������q %�d��-�k]���0�o @�ETO��&�=XC��	�M$���>��X��֒�O� 7J?�Y�����7ϱ�0"R��^��:�%m�'����0 �f��7K�`߲x,d�*�I�v!/ǳk��쮂�Je)��J-6�����R�A��/�����L��k�T; ,�\�X=�(����=,s��Ĺ���h0��o4S�@3�/u���5/G+K�z#�����r���D�3����}i^��r��h�F�4Y�P6�-� !��|���l�w�  }u*�׿�~�j
S�`D_H���$g�(����5�F�\���>�ye�)��?��yX+��%.l���NK���fV�W;&��b�J~��ݪ�ad����4�#��-3e��g�+M�ڔO�*xަ���JOB��$��^i�m��8�s�kv�fW���B�z]!���T��H��E�6ָ[^v>Z�S���Ս,��$L,b������]���)�ճ$pɗ�>�J�S)B��@�ȋpe|�ٺ^i�SpB	6�irv�z�#�x����J�ШϿA��y+�\�)�N�1���F�ԌV��J�����\w	�h�]�$��W!X7��a]��5|X��uqz��� �7��W�ϕ�	]fi�ր/�֊P�m�͟J�7.��Vq^��}���S�e��9�w"��4u?Yy2��mlj��L�a&�g��8_y�dP	� ��9����(���\� ����O<����
�P�$�Ă�5��9J�B�x	� ���Te��@X���n�3=S΍�K�4�������� ��r?,G��Ӭ�	�[J�j�iR ���9ޟ#r  ��{?�)��lhe��Ѱ�u�*�	�e6���_�!kla=����Ve�&-��u5a��2�"<�$]&��\����x�$IN H*�Y�%r٫��Nf��KO ۾��%Ґ���g��ro�^\��Ƌ�,3A�O� ��������_�|'�=��`�MD>c�֥���w�_��
s'}֕J�|��1�^OC���g�I�� �����iX��)B�U_�pk�]oZ����5��w��Ŗӻ�Y�syI� y�<АA���}җ3�g�s�Ho4�A4�J2���}�-�4c����k��[NW�����$��p$�M[��m��"�c�߱v�1T���K��R�Z?˥�b�T>+l|&̵�n���k� ��t�Γ��uX������ҌUz*�k��5�H0��ٺ��g�嬘i���'~�h���˂��9T�G{<V��V
K����I��ک�I=`�`�S��S?�ga����y�i$g �'Q�:2�اA"�
븜AI�\B�u()}��Z��a��%yQv�qޏ�$��� �Z�e�� _~v�%<�km=W�U�=P(�c�
�?�Y�kc ����o�A@^�2Cԇt|ԭkF��X��λ��;��F+���I���ɦ��o��LN2��!��v{�j�m�u���Y�V3z]�	^�2qV������eڪ�#��+�
�CIA�'�c���jr�Ы��h!�D�'l��T�٫���=ZO�w ��JFr�I����;A^�ʪ�8t ��56
P��Do��)(b�*p����������Bh͖��E��V`�p�+XoKC��U��v��LeA"e��p[�ɹB���t��<��ҁ:c���绝����@�cE�-j�#'+�4����
�]:��yi����#���3oͪ=�V=T������"���Kc���ȁb�Y~v&k��xŐ�A@�h$�ϲ�8�_�%'Xچ�0��7^Ww��0C0��k�ܟk�M:��:k�u�[!-Lm �kd��)9����m����N��t�Wˌd�	X*�r����L�Lf�j!�����	�FY���O2����2~<����4
=C���`w�	8�w��߲�8=��B�0�ǐ�Y��K�a!�M� �}�֭�����A(�����s�jCѓ�E�#��P	�����`o�7:*a��\� -��F�ն�;��]{��0�<0���^����v�ن��ns��	k��S�Kpo�ɰ=��믟a?�Rt�pw��e*��9@ޚ��0�,wĢ� 5,w��e:~�?��t�6P�3��{V��&�xz$�e�$.�~�wO��W�S\f�F.X�,� Nή/���%�k�4Ky�}���oYb}��P�g'�kؚ�,W %��Y�n?���~,�jE����*������x�X�������;��Y҇���˹�г;��9���Ӏ�g9 �D}��|.��ѥ.�#	���]��"z�a���*#��)�K�]ԩz�zfG����4�����^�y��&��_7ֹ�%�[�q����)��>�F��D�ìг���X���sE�˾e:�J�)d�Z�xo����r�%ǿ3q��:��1�7����e�DD���5��*C�Z�}���/���ż��E;���=� ;d�c�W�bt��
ء�w&CT��+V�4n��S
��0�ZfŌ���x��hh��y���5�P7.:��s6��0!�v�Qk�z[#���h~�F�αC�yӺ@a��Bap����uE���i�[ܗ-AF,��SL�\���R�ū��Ö}���G� ��y7&��z�k�6U�=C��=d�l�+�d1���D����� p��G>�Y�T2Y��D�����ƙKzʝM�Y���57#'sL%�9���F��Cބ.Ac�Ԯ��z�00xm�	����Բ�%���\w�N%�78�L���iu��y#K�*J�c8!�$��3��`��7�+A�:9$�8Њ/�e���-[[-1`�n���5H�?��K��L)x�F�@-.f2a=��d�	<qd5��k�JA���)�jr.kk?�w���Cϭ�]��R�)/MZ(�,�_i�
5�� w�,aM��s�CtY�~Y��P���9[��� u�8����ѫK��t.��+�J+'x�i�t&�|.G����8)�b&M���y�Ҟ���4�n�2�-��V�A=�Y#�Q!�zx]��{QU֞��.\kҌ��W}�D��R�����SRX����3=TR<)�u%=�-�� 5,,�m3 �e�R ƽdS��ow��5c�k��k�Y<�
ʙ�q5l���0����E�qČ��H��lWy컁�'���hϠxGP�#(���﬍o�8�`��ƳD�x��R'�#�Иu�*��/�.��i�rngQ{�b���Z� �l�X$P��@j(:ݶ
�X�f~4��I'���g!oj����t��_bG��>� �X�5i� J���2"�#|��+�S D������<��+�=�2���J�\�#����G�X���7b��81z �c�r�4a�;�2�bްM_��eGz�#�f.҃�z��녻�pV���y2����<K�{�4SJ�Se�L�!��Ӆf�
���er��K�����L<�̐��G⡩����һ{��·E�Hc��W�����7�']ʬ����|�n�jG&<+ *;�T,e�i���"߸X�yw�4��ky��a���_.Q���]�;��d��g|��J1b��h�mJ�7���3�@���bi1^��a|��9��~��Qw~�����}|���z�{�Vt"5����u��te�Z�4�v�]w�N�G]g��u}���R�f}�}M4cA����[t���Y*��#���=��T�+զq>A�WAZQ��u[a��P�e�f�W�^8�������� �	�Y���@=w�3Z��"��R,�kr�����귮��b�Jf�q�����p��mk��y����D�@`��>����j�VBD˄�V	�q�֞tˡ�|/ԛ�攵;c�<��u7����g$ZW���߷0-]�~n8C
�\�~�Ic���f|�6i��P7w'�1�a�>���`8A����|�����8�;�{��-S��=�>�k��#��?�a��3Z[xB���>��C�r]d{S!����ֶ�v�"7�k��^`0u���hn�X��C�5���Qӵ�k����L1��׺o����D��5���,]?�%�ck٦#����w�c���ㄲ~���Ŋqs�V��@M��)�P���S疼��A����w�V�ס����A��V
H�#%甠��U����9l���CH@��S�ЗR�.���q��BЛYXqZ(X������kY�0�E*�.��h��%�&��V%+�:��<��ZW�Hq�mλe�ݰ��S�g�%b�C��!���k�뗍N�=�� V�k�l��!ø��X�=K�;��{s��y	sq�1уU�����њpt_���w֮�{���X9<�he���I%�1Vs���׹�LK��+��R=X�Z����y��o��i��2��VK�w������;��f@_0Q�i!u���2��]̶�\�q6	�����}h�ZV50���e{T��%�嬏cgҟ�yz�jÅUؚM�<�����Yty��y�;~SHRi�yt��]�ZH��e��,�43���o��d9�N�,�E�ʝ}u����0΃a|��u�K#���ظ�y�h���^߹����{j�Rvߠ��ukzhY���at������+i!(��Р �4��k���ҁ @���k�iX���v�T�r�|g�ilk�&b4�����r�<�]M=_3g�~��V����R5]�׎�LC�
>C�;�f<�_��2A�>g7V������������*p^M=y]R�z}�j"�o5���b��H�%�෻2�7�gku_6nG��j�%��,l��8���O(m����Lc3�2oGٱ�����8�Y��kok5�ݡ�0�^�"�Լ������k�$�f<��:(x;.V�����u��Ik9�,-�Ⱥ7i�����շV9��G2R��YH�\�>�2�G�փ�='�J�I$9y4 !C�Ό���+"�8FQ貙|�m�A䬙c=X,,[�ъ�V����R4�]:�r��T=Le`�%�a���e2�M{�4x�ޅ���!.I�Z;I;@�ϗR�S-^K�ĐO�$��H�]$zC���~�Loc2���	.6c�:�Hx������AU\��,�>�l�R�MaKca-z]��2{)�8z/4a�q7"�3_���$j��8T�1Tn��j<Q���b84�7a�e�x4`�P2�>Z#��?��� ��U��b�<�>ϔuUo���/�͍�餁ᄯ;��l-��'�UGu`��}�4^[X��5K1'+<��y[�\j���g�}f���D�:�BN�
���^�����
� ���{	+4ֺ�U���Yb���!��j�?k���
 F-�j�����
�Ι��s��f$)g�T��ֺ�wj��e� �M�P0V���+��E�[�`Ĺ����֣�}�ߏ���`�1L���o#��Z;R�2 ���R�������r��y'ӕ;%��zk����v�G�Yz,��c~�H@��������
+����9 4 ն�E`�����{���CmY��X�����D,��S�Z�	��Λaݢj~a��y�i'����b��m��\�W�2�G��QmG��^�cؙ��cs~�K^t5N������(���E�i�[ߪ��A�X�􁂥B��4�6���Жq��잍�n�+GH�ђ�d���3�����7c�ۄp�0s�j��LD����`)X�&1�+��o�V�m".���%TT�n�dӹf��L��^lK�qi��l�:�,G��3zk\�I��0��ckv��k��.r�ֱpe}lZ� =��������h��<�E� f=W�Q;����]���k7�[�s�W��e�p�zwl3�.��sz���ru7ssiQQ�ihdn
���wtO��B��e�Z�YB@'|d�P�k��1�xk.�RI<�����_��?{$�y"�����O �F��*���G��|�&�.��x�!�<�Z�N�]�5Ĭ�F��ْ��
J�|��Ž�k-^[���Tvߵ�i-���+�R���V�e��R=V
"]�&Z[M�n��_s5ݘ����������Z�X���eMj-��g�S�|���̮$݌</g�L��R�L\Q�6N�m��6�z�|����\�2��xJ�:fX�I�7�4T�r9��0H� ��=CA��ڐy7���Ǖu����9W�˴�cz9kS��5$��g���T�k���D�6vm+~U.�D��7L��B㊡�})�@�̬���e�FU�'"��t��%��m�(�'�Q<��J�q�{�k)����ʵ*BmJ�m�z#��ٳ6�	˥$!�X)����ï#�h3uy>��
����z�g{�^��Ϥ=�
zQ��Bn��p�8��s r�ӽ�,��)-%\e�L��{����s���ݱ�-��Hy�>�� h!�K�r����ҌH:�]�.�I����m���h�Z�%�>R�jlQ4r&]�����?����.��|���p�6gB�c�8P]O���H��=M�Yg�qe��(�@y�md�:+-R��t�p[�����wo�ʯh9���d�y6��mG�v�3*�Bɕ���/���%�(�i�����b�K�<����s�w���J��=��d.�����U����W�������bǅs�Xa�$���P?0k\���6��MxD�.r
��/z�Tٹ6c���#�5D�X��.��Ō=I������snR�D�U���Q�K4�M,�[����wV�؝rP���p/Ќ+%��|Z`-��1ڙ@7i� ��!�U�gC��^���f-7�}$Xv<
m�L��%T��:L��?�"�*-@u����Cy����ɯ~)��S9�,.2%ÓkR���Wh!�M�����u��r�{@I�X�
�j9���������%=��~��rO���j-��@{�6�OY�jf��I`B�B��Vx����*����nzغ�vV��H�t��X��n!��Қ�,�r�"q��OdN\�h3$<W��V@(V[b^��X�9��OW�.;�{˗_~)��g��
��D��R B�25Y�s�d�FX)`���]��ķ㚝n���Ęлflʗ��y�"�ψ�|&4���+ľ�%)�}�;O������ʄ�K�k�r֬I�p��5���NUۤ��(kf��yY��k�|V��F��Z��i6\�|+fO�����2��������4��̔�VI:_�;�=[CSd�vYl4I�酖d���.��E>3����6�`�rW9�_d�B���T��-�^��ϻ�&��X4)�Yڵu��g�t�=Vl<H/\��R'���@[��q����2�p����+K��u���KX:^g��]���`���3}=��Q_��sU|�1�i�T_�d9�����H��|�!/_�m{������g��Q'n��YHߡ�C%}�"ԅE X����*I���И�Eyd�Nx�&��nl�H*�[Ť������ͦ
ĭ/������l���.J4�Xb��g}��<P�O� U��N����R/�qz�nT�~�� ����P����)��r�V=:�]	�d��m�ҽ�T��ԚF��9j6!�?ۊ�׳&���y����B����aXF�\%F��oi���7f�a�R�cg�(J6X��Ȋ%�O}Wǲ3\U^f��Q����K٭!vKȴ������1�����@̷-��B����=Q��|>W�GA��9Q��M��5�2am2dYiȁŎ�M�񰱼Ic�Q7V�Yl�u�`��X�Z�X������]]Ҭt��$�2������,�8	�pa@K����ʚws�Ҵu��Y������2����yk��)p�j���bf��.����Tc$�����2��I�cМ��w^���R��ߦ��ǻ��'��q ���� T&}�i��n�o�Ѝ�c�nf�Оy<͘R ��89?�~r���&��Ձ��D�P~0�<�_�����㙑�V[�_��+�к�-�L�9�e��G�h*1w�]��v�������1�~�Tb���LI���sF=5��m�4{z��Ʀ?#&���L�㫽7��^��&V��s����CW��u�H⧵��qe�rm����s���]��|ӧRy/�R6�_Q��k�bT`G3��܀�u9�v
�|��I	���/I �r�g�>V���,c���<P�0�M?�5�~a���	*(�S�$�L�MQ�](�3ŝ��R�T���R���~�Uh��D����el� �Am�\����G]�\���t63o`x{��%�K;L��ˠ{`a��Md�1�Ox��P�A"�?3�:$P@�	p.��v�
Ta��d�u	�1�.�3)e K�K����z�!3�[� dgǘ;#�Ӌ� Q,k��'9�[,���D��G^K����=2!]��¶�h��Qt��l�N(5�3=il	J�m���A$�?��� �R<d����A�[G)����}���M�Ul?l�;�y��:]$�O[��e۬q	�*��t¿	s��n�O#,/ց��d�����9�q�d0q���>��MOt�?�d �50�
i�A�U����XU'�����b�^�m�[ɼ���l��j���>����z�iiT�
ٻS6��9�.�b�pSxbJH��E�� �k���p�t�׺���r�w����ŉ[廴e��G�����������P�+9�m��td�����.$��U�V��B�Y�b�O(�a6w���*-��%hR���f��,��8�4��-�O%kv�-�n3$�c�"�`�k��� ��g��|�ʙ8Md�,��	k��z�q�����6B,?PS��cBƵ�� y�d��M딪g�`,�?���Kt�5��� B�4D��g*e���/����7��(��'�>W.����/����O~,�O2{�\�S��o
LAhk!SZ�Vb�$��^'�p.Rp!F.��`�����n%ʝ~��n�H�Դ�Q�;ߕw!�/�~�rr}�v�
���&�tcYk�m��ɻ�o�;��ZҸĂK��Q�����P#�f8�dʞ������(�"z+o(�s��k6/�t��ls�&Y�.���k7k������� ;�uM��-�O%���	�6����H�X�(Oh�b��B�W�0w��\5�k�\���ۆ�U,M6{���u���X��+{��7Ț &�>�	� wK�ZP���\Wv��; �y����<��z�� ���g�<&���oS*���ė���չq�N�<0
=ƌL�󤓢�g�@���9��i��3��no�RY�Nu���>�҇i���,��Yv�*MB�z�D+���={�ם3�,��g�ql������Q��T�Jʌ_ϸ�ԉ�Tgyf&_=�]�7"��wъM�}����q����۲���¾��ob?U��J]�`\E�R�H����-�L^��¼
畧�!P�͹EP�$=}�4KU��������6��l��/׆\T�Z�r�~_��D$��K�b;>�]5C��DJ�w]y��2U��4M��Z)��q���Eb���`�)��VpQ
,	A��i6�>�nЄ&�+�NO=�Z�B���̭]�FB4��,��s�fe�z�\�x�����"��Os哄�'#��aY3q\
N~�i�(-8ش�p�o��v��
��7�>m��o�5�4�6�2�|M��Yst'+��)[%1�� �����_$��X �VF�Xw�$�c݅�]��;0�v����;.�\��;�Cy<����r����Ç�H��ߘ v�)��Y̴0hB�ŷ9o,/N�"����x��H�	9>{�����g?���U;D���`|<M�
v���5r�����\AV��pQohƅ�đD�s�8��S�N�Dڇ�|y!i7�͎TnSc���h ��ՠR��ROZ�>�R;�+4�w���5Őy13��뗌������5�-ˌ�ʕ3j�Ѡ�{G�mB0��4��ڝ王sW�j֒�Z-m�WxSwˍ%4Z���$WW��b& `�A�piש�a"Af-�zB/o&�c2�Ⲹ�f����iI�Y� ��8�tG����y��D9�Li"�v��ڷ�
��o_z��H�Ik\io�v�_�v����:ֲ4R�PAe���u�ٙ,�̢����.1�Q�py�Nn.��� �?�zu_E�ƍe&V�uc� S��/�?ŭWL�1��g��-�Cl-�i!s+�ywy�uM�˘}���ylt��}]�{�IG�����ɩ�AX�lˮv$�Q�]�F
�����}{��/HY�9�z�טѫ�-�Z��t��W�ִc��IF��D�cǪ϶��S����%��4�XF��hLE����Ka�g�fS�D�VF��dc�(@���%��f�gWZ!�P++[� �hb�ϵ9|ǟ5)P+�x�j�>�j��/�#C�{L���L&ʅ��u��LK��6�:�������O˴֒S��25�D�!�ڻ�{1�K�1�2��a���Z����r)y�VWr���t#�!�xO�j"|��P���*�d���N��Kd��vH��^{�/����i�Pj�p%hb�s�eOjk���5����a��o��J+�QCМ��p��L� ̜eK%y��@��w%d�FH�G����6Xܲ��D�FSy�������F��_�􀳞�T{^�)��M�`�m�^|R;*���KG����H�7�%j<���+?�hL>��:cc��$]A z	��B����M���_7�Zъ\㴭s�G�D��O�9]��Rݛ�����������Sb]��io:�2?��xa� �s���s��W�Cn����o��MZ�ez�>�`ON��sV�?�WO0���Ζ�R�*����~����p*/~�Z�_�]�TM���+�}��A�z뎁�t�9 (��Y���Y����O*I7i��
��i;3�:�i��Z{+3l�A�{�B0�ݭ]^��"��9+�3���-����Q�Ɋ����44K�!��O�7P��
��b��ҡ붡�i��)k�Q`W�Yǡ�>���l&�#�h�A
�/����̝��sos�@&�c�P����;c�u�-����9z��`_��\����}IbW��=+p�[��k;^^����z/l5������W�eUX؛`^���'d18��5CA��%��'#�i�Hw����b)�/��w��(�Y��e4i���:�P񳍚�r��i`�H\�h=c"= �������`�%��Ӿ�AL5l
�^�$�;�Q��xg��s⮷(��b�K���Ҕ�B��{�ɦJ�!d��E�FÀN�A����}jfSWڤ��f�K˕�hc�!o|d #WAxC�w]P�VZJR��S0����bq���xv��U�7,���X]5_�J��3a<����#�#^ӳ��l�.�p�9��F3��e�3��|M��#:j��hO�p-�9��4�4"�8jV�֧s9~�\����]6��9�d��7]�s�lt	p�@�{,aU��E���}Q��iln�(�teK�$_�{q��=NÑ�cG.�2p�ے��!�i@q)�3�9L|����/�:B�j�2с���$J|I]�;Pp�*'���nd�!͘�+����}���39��d���ށ������G�+e���bU`���$&$}98:�񽙟H��D�?�|Q���k�(�#��x�lg�._ag�ѻ�bH�c+�����]i�=���2s߳{�\�3g;�z�v���E����s_v�z|����He��� ��ܛ 0�L�O���L~7?�c�loغk��R�)��Gj�[4L�t0�o02�Xz>�a^��O�%������C����"�fv�m����Aw������z�|<$���>z������ZD�,:2�#5O ���S De[a��%�xh�|�_��J�yZ���N��!P4�3V��bfˏx��u�������@]�9ˀ�.��W[�VA÷,[�u�++jYO�dr��ǚg�s�e�N	'�s�\X~��t���p�Æ����g+��J�Ŭs�t<G� ��HdW���M!]�s���3_�`La�˭8y���"�q�֧r���D'� ]&��5��]f�e���>�\��Q]�m���L:�i�Ֆ�9 ڸyS���﹟Yܕ©λ;�qH/�y�T�=�g�l�(�n��R)H�<�w�����O����d��H�υ5{�wc�g�6I��B�eC2#�_*g�߆jE�������ʅw�|�2�=���w�R��Lr�jM,���ۄ��'2���e��)�k{����z��\�䢀vmX��wz�y�B�<�1��4��p"�����,��3��|�
VJ&��3iWk���H�}5���
2PY� OFP�)A;��4���T>Ź�uO�Ɖ��Z�@�`������=�E��f}�Z]b�Q�T��=uIQB���r1���,�> w��}�o�w��,e�Ve�X��MD\��\+F�z�2\�'�ܞ�J:=_��ͱ�����r�o7,K�� 2]y$u�X/u�5��4Zl�V H
BH�X%��u���j�V� �> "�P��9���16�D#/y�w�D�hGG�r�B��y�v��E�8v�E5!�{�v5���3�(N4��CG�=�D�l3pɫ���<�1���U:C%�I��R��h�1��3�&���f��2��J����Z�ne��=�\��������6}��	�A�g}^�S&B�,[�q�:��on�4��/���BN�f,�Ik\v���`��F��H�o�F+Pj]�t���`�l��wk�j���&�i�S�Is��B�H�X�����'j����_�y&3 �9��$cFкK�&��0Qk�n�b�t���	 p���v;�a~aPA���7��d�/?�{,��oX0H~�Q@�WK�2�Fk�~݌�\�/�ڭ��W�������S�"�{��"�gYk�W��z��X3���H�u���ʜ*,5;Ʌ~j�ҡ"d�u�~���eu`�.�e�˲�g+�c��Jϲ��.弪uO������������Vh7�CwRU��� �?a{ K���z��%�|��sі�lO^4|��Z#��KU� ˙f�V ���,��F�ㆪ�@Y_����	_����i�d�u%vޒ{fe-]K�4 h� @B�n"�E%QR�%͌H���#�a�P��?��8�	َ�	K�4�diD�D��$� �A �����k_r�|���{YU�V���"���2_~���z�9�Q���Ђ��3>:��bkj3q� u�F7�ʹQ9��8u�.0ba�1%�f��������E~� ��JLL�p!�nIVs�O�oʕn'��d(J�7qp/.����JL$܂�8S��kq�ˢ�b�@�%@
y?6[�`��	�l��T�'v�ef��%��M=s_+�V:���pv֦��@�뀛��}�M��ҹ,K���i���n�(a�Ö|p�����=s�?��=���&D��9��4�.�R��ы�K����+�M�Ҕ]	�"9E	�:�=�M�Y���o
������^KF�b��w���]#9��j33��<G�a/�(�^\� ��D���#�Z��=	ueI�=:��qSj�e��J���@�\�o�Fmf�[������Bw��Z�1���.��5PMw���B_�=��%�0��V�̙6?Ҏ�����8�!��piL���x���a�M��lcG����w�I��J>]�8�8�z�Ȃ��z(J�B}g}_h�BO�=Џl�k�6��U*��'�t%b�:=	��i��or���3�E�b+%�}���5��H�^Q������*
$^g�3��8	��N fD��3\�A(g���l�Pl#���Q����@��AQ�S��d�iLbe8��2���[lNzD�� �>�Ʉ-7�vg�X9��h4�;3uJ})Rc�N6�4�t7�z�(�����,bE���Q/K�}ju�֗�-P��#��J�F,����T���j�QTj5X��r�EY̢l��|�g���ɓ�����~���D��ZE�,���z�.a�,���w�.F��e����arzבH��R���� ����5C��Ls��C#��ب����hwצ�b��I��ֻ�I˕�+. v��_���g� ��lv�Z��[����`8�ݦ�w��Zb@���+:r\��2�tSu�F�����q�Y/נ2�~i.�Nͣ����6
g�D�nY�6�4�dp�w��e�+A��8HRs�=����F	tg�.��Dn~�4�Æ�P�N�#�f��!iR7Ȱ�2�o��w�ƚ%ÐЂy�%8��$%�de���! �NՉl�oH�Î��skc�Z�f��g�LŃ�|u��A��U �.�i��3ܔ�a#�L�a]�%)�À��-�i2�A�(+;e1�*�$�"{AcK�J;�H^�� +9>�S�:Q+���+�N�㡳%L���P���LoŊ�R8S�'���*��1y�:���mv�?K(�O�����J���Gs�R9c�9}�\sI(��~��U�T�Q�ۂI�!%�����������tb�/�R��j{F�ZR<lv���mZ4�$!��~)��v}�:ܒ�:�I^:�(u�� nÂ���G�`��1�v�Ê'F����0z1r������u
t��׶��-tO&�A�m_���3G�Pĳ���ӎI^֌�&8AވV�J��Œ��tBbIvZ(s8�wq/h0���@����YE�0J��&t5�F��x)��]&����K��I���LudT�&E��#��gGk.�7��kl���6�-�I�N�H�m���k�2r��@۫`=7�n'1�<C<%{�~��]R٬&s�)�H�P�E�%G�΋����d��g��U���:JՒ=�y$c����n�}�����_�1��z)sw<̐W�}h�HU���!4��+e+P2eA�bz��~�h�:��湌R��H�G�(�G/RZ%V-L��C�[]�+��X�XvU�EyP��p��
wއ�wă�>���)�����c��7��l�h����W����ԛ��ԫ/`AW���`n3�	�+�6���N��;je�}� �,��r:�����sՑt��޼IMv+�Z0��j�k�q�o������Uo�+��{�k����%�~�T�J�0��%΋��2U� 0C	r�n�t`��U^4Z�����6�f,�>��Ũl��8�+�a��c����9#gc9��/O�)"j��nl�xW��ٛ���G�Y��Qc@�JYۈ�Kȣ�Ri}kY�s���g����p���?��c�lLsn�
a	YM����x���j�&^[�>�tft����m� ��%u�*R�����S�v/�wyt��5�t���k�5Rc?5쏢t�L:[s��Զ2��4��q�'qeG$A	�Xe��� lHC������ۀb�є o:g���c�W*'�Ϭ��h�ht�E.�*�-��*g��5˽����f�o���Cǫ���FbCZ
O�s�����X%RUO��S��#-I!0޼ȴ05��M+�s�s�����!&/k��@��V�v9�xǴ�#Ό-�̮ha�<�yq��a5B*1g���F�1�f�;����*=m]!4�EU�)���fX�U��Cyl���^���%	HH��O�%��L9h���TZl��BB9�_��el�rQ+�Z)c�����Q)Ø+��O����٩�b_��[�m��y�/�/�L따&H�+y ���c��]Ww%nYqW�����7�u���CL^Fʺ_8ɫ���R@����Q�d7�P�u�oʾ���"��E�O)��&$�V�x%�������ϛ�R��p��Ϙ����U��H���aY�͊<���"�����K|p{Bi���l婅Mb�9d����r���]4/I�q�"�^?f]��*ُ�rQ�u�q��5!L����~�$c�=�9�g������A|��3�$�U:-� QZ:���\��Jt!_���Ϝ+VQ�Օ��F�MSe�|�*�����*�MA�7C
�`����;P7��J:˶!o��E/ux�TǇDjT�v
�g�7�HM֧!���Wp9�3��	���/ft�^��ȃx��?���]ȏNHP�E{�
�^;��ښF�ğ�2����K���N����ã�|J��c�W�Ƴ?��o=��o��`�CĸN	:~�n�˳h�&���KP~������ߘ��̥I���RmV��n������iqҍ#3������sh��t���}|a����F����8嗈�b�fm�ېuʜ2i"R��)n~�}��>�Si6t��PM��^ޘ��+�g�F�U�1�6�
6vkG��JK�^C>�|�R�^���⼂�A��IV��WV���$�fq)\��U�r�ކN�׉9al%����$_�2��[��m���� I��lņ���{.�Bv���^Zg��8q}aI�UC�����*�V�S<,��{���rjL5Y$NI1%N�ҳ�wr�u�ǏD}mR���U���L�w-}7�7Q��
:��� �ߓ���jےo�����A7�p��K����b�d�]|��+�Nn��sz�����Py�S������fsU���8�(���bV�S�MT�Y��@m�R���5<p	=)x4��|���O0!L�r���	�g�;I�DEVkyOY�vK%���ր�϶��s"jI������h��2��gQ<l{�K�;`,i�hV+��1oܺ��]�)eGI�3[~^ױv��Z&��j!D	�mG�3����F>���kxYX�,��&o7��� ����ܱ�8>�Pq���!C�=�-�eyr v#M,��U?�}�q\��d,���zN�<�6�zWU�6kӪ_Hݘ��1V���c��ib;�{��#�`�C���w���sp������&��SF��)�w܍}����F�c�q�ŗ�r�4Σ���U��o1Ij*���d-4�/�k��q��թI�!$�i�Lщ,n�rE�-�.&k��*�v�r��U=&+Qw��w��c�ބg��A^�Z�Q�he�*$�U`,#�Ԉv�46NܢolN�e�y��C��9ՀO5#C��SQ`2%mR4�`,vZ�'�Jo�j^���}�P9t w��1���#���{��&pj��Wq��1�4��W�5��µ�b�J&��#u��L�{�1L��(��x���7�o~���װ��)���Q`�P�پ���+��}D�ݹP�Q�rEm��u+�-U�y�)ݞ��_��S���0�	D���1FBy?_s�\�]@�9�r%�KtS�Փ�A�U�o��]砡UC/�En>~�|��v��ʍ���o���aY?]l7p��Z�ֆw���\�]9W]�6�$,�����Q��(��Pn�Pl�#�9G�O�����v-�Ċ��ڞ��(���o/p����wG�Уb�|�%���YCųAF�g�>��\V�W,GU�����|҅DjT���o��*���+���.�ք��q�UW}O���t��S����5T�Pm�ʾe�0h4�5�@��[��5 S,��QĞĸI�l��Rp<�;JӐ�.Smk��,��N>�a#mS��3�kV(l�X�nj�	�����9:&V��~Q�YZqN�;;�z�ifn�&�1	b�6T���S��T;��Ij�9ʪ�ME�D��m����$Ϸ݉ĦxFW噜'`���t`��BUu=}���m!zv]]��l*�!ol{�8*��+��^�����S�����nM��B��Q���z�Z}yyeY�ꛛƹop�:<�ʪn�ʸ1r#�������R�XB��Y���zL�0b}M��6�)��UL� �7�S���z�s��VQ��hG8X@�P*���R
Ѥ>���ow(�]ڔ�$�UCO��R���cl�eS�W���_˿�W8�XJ�����;�;��N��S�D��4�Ò�o�̭ :�ss��&�w3�uu btt�S�Q��"�?���=������q��7p��/`��������g�Rmr�s�Tt�Fl�tG��ɍI{��N��'��k��ɮ��ǉ��a#��-��K���m����ɯ�ّ��-Ao '������������!��E኏�MqiED�7��7{��݀ө�1�Ua���J�Ѽ��}c�/��=S\lp����H���܏�o����G��]����/b�ￍ�ɳ�|�$Z���G_KV�$��WU��h=֏Oq��/���_I�vh/��܁��	��=?��?�y<��������=
S2��XBܒmXĐ�0NEq�:�m��`xD�ڔ{+�[01�� �v0?\Wb�
%�e��3�����Ө�*�D��ß� ��7�,5m:ڵ�hxt�<2�Մ����o���>���bB8Y���_��ݱl���ӰT:�nc˅|F>�
D��`�a�f�EӃ���B�Sy�Zbd�R9��8�Ke��Ч��PM��I7Qb��U���A�P��M%f�'����������4:�4�k��U\�_�H����msed�Z5V�T�Ir6)�N�[x��J�u��K
$I��3U2�:Z��M�g���z1�i8pt)�$��u��ZZB�� O$�&2]͝\J倌"���ĩ�X�Ά�SS���<G	��إ��@�2�ʁvz1��gB�I(K\��x�`�p�n:��f�Pp�E9�{���?���k+��C�-����9g�]��R+>^Aij��u��ʿ��X'V��G+QF��VG�#:-�o��W-�S"vg�h��,/g]�J[����b�VOmz=�]���9�}KF�O	MNͪ����UL���~�y��ʣ:ZW��z;<��%��p���v�����gR[֭Q�d�8�2I��8�V�+I��d��Є�^�i�ÀV'bC�y�PRŪ�s�!�J��3��'�	M<��riWD����2r_�M��л� ��\�=�c,(�
��B;X�ǽ�>�����Q�CbX���	�o�A�4[�okkH�HZm��M-&�+�1h�Z�j��Kb�ğL��~�!L>x?�<��{Sw݃���v����^A�n�o5�Rw�JRXP�rOb���Q�Z�=�귵��8��u��F�e���T��=����,hg�ZZ�K�vbR��*�5ɷ�e�9yժd;��5,s�1��B��ʮL8p�΃W�ok]��R�>5��%�ʴE�"͋8���@�u�Z=�|�2�qqX1۽�i����_�,��/|�ａ������,w�U�4_��U�dS]2�]��h4��y�N�3Y*.`�0���X<�f��&N��W��3���O�<����F�_���O\��K:�g�..^���9S��3�Q$���,[��8B�ݥ���k���[��3�EU��F ��]x��!1�=/��JZ��S���ߓl��wE�x�m����".��:�r�B�٠�Z��6�\A��j��eVW�nBs��FuJ�[�̱ݑ�5d�]��|�Z��A�d�}k�k�ǀd�[��b$�c�0�W1���<�gL'I�m��l��;��Ƨ&�ޝ�����7q�DuYǑN5q�����<�9��7�L%�����|tŘ�:�t��1$*��@#��GY��j��I�!�%?�o�#�����B;^<�'��@��<IS�l��i���cz쏿���U�z�N�,�pd�W��u���Mp8Ÿ=�
c30�>,un[��bM}�onD����J��7bq�E�z[n���	�3k{ў��9�������;}tW᭷Pa�*��N�z}�Q�d�L�	���d�B�Iʁ��]����0��K�?g�˦8>+jn���3D��*[^[���P9�xCNl88'Ϝ���求�˙���hڦ~R�k��u����ÁV9F$ �J��M_�G�PU�p*��w~ߩ$�*����$��tD�fQY�����R,_l�U���Nڕ�P>_��ϡK�3�/v��A]Yl.[��n�k+[�&tҟ8��N�B���e=+��eEl��Gd�D����CM�;Tӷ�M={�Ol�\��F���A�Fz©�����-W�t�Z�7�k�QvKL�6>N�����FͰ��ʊ�</�OAQ�j�.�[|h�IlˮRM��������J����Sɏ�;c��U�{� ��:�Zt�GⱖCn�rm��\��J�6=3���W092����d�n��{?�a��/|8tx�(��x�G_Ù�Gu�g�73cנ�ݳ�U�)[O��`��|c	i#B9'�tqO���w��щ<�ػq�G~
��:��|�+������h~Nֽ�g�V*�k���-I<É���$�r���e70�&�����V,9}1`"@�tV�e�"�f_���7�O�_���Ňng�O�Y�k��1x�)@�P)#lK�� �l��r6��6�b�R##�K�6�饙D��.���5��m/��R�bi����:��$�1�3���_�E���wKM���������h�r��*Zb�eY$�0#9T-��=-y��~z���'��0V��l�1��7İ������D��=�<>��~�~�q��$���/��W�&�JLK�����,���S�eA��L��W+���{tb%_�7)����@��s�Y<�3�9���ts���x�܈<KYWf�^-�j^�� �aq�2&�FD�A����e�Đ��;I*7_��qSs�<V�WI1H�79�>��Ub3l��M��.а�@+Qċ��^Y�̬��T+h���Y�*�����B�R@~bD�Y^��":g%K[i�.���k�f3#�:l�b:]6akpox�K)TT�<��d�9�KZ�|u�����S˛���Z�9��p��Mө�1������RٯAiD�yU:(����^��a��Ǫ
�<)IX�"�֋F�UI�|�58�N� @����~^����
������Ze�Afe����6�4�yc�W������HK�J �	���(;��ﯡ��nz�g��]䰔*�ζr`D�4�:���4�V�B�LMYiATQ��+�@8�Oj�\���ͷ�c�ĭ�G��Bߔ@L��W�����3=K`"�_S�,��qnj͝�*򴳣�n��I���
$�rN}`��D�$6�P-�; �Y���&zZ����xQ����*i��O�����jJ9ܰ�q��W������X�]��H��<� HUr�~U�b8lϭ�@1��(��U���>���K��^����� G�c�Ե�s��Z��(�R�B����{	��R���u�=H�}�JP,>��sm�ۿ�@k=c�vy.�H��&o[��Z�F�5��_�����Ï?�/}�����?�g�#��%���x�_F��Y�f��^@//ϧ^V���D���}ÄO��f9D�DQ5���x}��~�Փ8�⋸�����3x��?�A򙵿�������#�5,T+H;��1P�Er��d�2������oÆ�����@#x2��,JC��/(�&�px���mHk���AcI��_2��q�6=+x�z�� ��@yX%Ȉ8�����\����d�}G���?�;?�Q�z��~�_�.��*.�%��� �J�Aȭ"ie�^`�D����B��J0�̻ �D�sa������"���q�W>�g&>����������T�k�E̵���.��RE	��PI�ʙ��/��kOߔ ��J�T��۹�A,�����O��^�:so,�%�S����P�W�C���dr��b'���i��*��Ū/1��]?0
o�n�����e��p��(/h�{��y��8�)f,g\G�6�����C'��w��,�+�Kbj���v� o��H���\G�ې}-Ɋ�E�Q�lSQ*!<7	��܍V²0G����o|�[k-Y���s�$�H$�I0嵻׬��w]�*��+���MqHT��C\_vm�>%�q��rg"8���t1�-�y�0sTspF��9�)��P5ac؎�����n�� 𚿜Y.�^�=�k;��kb��>|lm_��3;g��}?�ioS��~�te�� �
:n�7��j7v����#�E�7�H�J��R����C[+��_�,�kI����Q�l�FӨ ���|;.;��b�M��S�JU�Hi����6��fF���}~ψbo�ha���f��c|B�r�=�ĆI���D�^#��T�+�ې�2I��&��{�CRӐ;��AYU�۾M�}��j�&~�Ĺ+�A�n0J����=�0>�a2j��X���v9a:\p�b��r�A�I�;J�+�;%���m;'v�Ck���α�j[0U�]Y�(7#&F�ĽM=&[Eq�&����t!� �O�a� A�|��Fe���0�G��O<�!������9$�8���`Q�u�ܹAQ%5��7��Q؃�k�=++N�A��J�cD�иP�nMRJ�<w�?ZG��<��_��?��(�K����GL��Q�@t�C��@}"ꠓ��ÛqW1��W�Z{���&�L���(Տ��x:���a�Q���>4.���5{%5��Ǡ(�#�KLp��`q�h/�i�F��5�����!�V��-/~ն�b�|mU��
�7xma	��qD�
��s7>��O�������^�������π�9jɟ@\.��abe�Xe��lڏ�F��h+з�?�D�m����:m����c�:�-�c����cKg�s��~�_��M�?�C��h#�83/�]Fnb�����{���N�d����s��&�2�C:���x5{��K��(��_�G�bl�(��.S��GJ�0����j	���r��{����0y��(���ON!w�006��x�5�e���ߢ~!a̵��ķt�0�W%��qT�&�F�\�aU�#��, �Υ�gH2 m��#�
����l�đ�sKĈKp�g��C�kk�C�a��*k�v���\�/J�h�R2ʘJ�y�S�Pi�#�m��9�3L�t�;���7 ת����\��7��*����~/݊��ځX�S"Ӗ�MO�*+<�$��-�\Omc˽��s��%g�d[����WWsƌX�����Ma���>a.m����'�=<X��{�J�)5�*"����AY%��5pPڛ@9���~A���|���C�u��N��KB4F8F���A�r�ukAJ<�&3�� �mψqup�Ϟ����M=7�ikߪ|��)�z��:�A��֐�֔:KU�g�|����$����tp'�0��%��('i�Bc;c`�D�B�@\)Y<Y&��Ӂ-~���`CWt�D��7IW���c������a�l��v���w������hK���F^��x�����P�+���(���|/Q������+��;���Q(���3��jF�3����L0��>�Fe��1�v�j�Q��tQ|�������'އ�K_ñ/|^�.\DX
�O��kS����`�N[�z��dO�w��k��ɑ���Y'�(�*i}��Q�Oz�-|�Ͼ��N������������̟�%��/���hw���J0Y�F[Sf+W��#��$f�Rlڎ��_jj%\#nj��bX`�����Bl�k x�u��%�@S��'_51y�"]0��(�ݧ�}*oKւ��>���:�Tj��6�^�P�ڲ /\��I"�$����N������8~g��K8�w_�Zs�1V}Tr*C�).N��@C�K$�z�j�	VV �њq� ˠ��vT�(H�WBD�o��_q�,�?����?���8���?�O���?��?b��iL���=Jq����F�r(�H����S�8qd�P�� ue��r�6uao}��Tػ���Gq~z�<*��p��4�uC��8w��Im
gw���^z���=������"!�=�����yW�eY��tT���]С���!%��GU�Ƞ��d3/I��U�E��w�ꌒv��S���T!a;�u�]�k�<�=�W����8�����u� w��m�Z��#�����ڣ�+}K��$��*��r�
 ~ݏѕ@8�*���5L˾ͻ��0�F8����e�ҢSZ������@>O_)tRqG��x-Yl

y���mI`��+l��ޏ�[b� �R)?�)�ۻ����|�q]������#�B<d4P�s��EǴ�̌C��P[�W!�ze�I�Y!+ ���-jQ��ݲϲ���i��60��B�"�^A3y_����|rl��@��\�/cS�u��h�\(������1̯/�����ɻz��;��U�:��
N$�C�/I���V]US�Z����uHEQty�V�د���%�̕�5�Q�z|�R�g ���q�lbX�$>�jU5?#�<��G��D��Ԏ���ʺ�y�j�|���~x�l��(�$����3��t��J;�#E 2f`ڱ�*}�DFq�V'�u.K�E�h����00��{�:�H?0�y*R�u�����s��t��T�8��'���{�[]ěo���'��ve�ӻq��� ����� J��_�J��lS'��Awn͋�Q�_W_�m7p{,�v����n�g�چ�3Z��z{���UI��S�8O���.�ү}SO>|�9�.������9���$�J��w�J����ـ���=[�4�
�s�16�V�	Xk���ɟŷ�d��z
_�����q�g~F�/�՗0�n#|h�K$�Ŗ��Z��vK℞��+��ʅ��$wȕG��b�#w�7�g��x�]H�.������%�pl} 6z%��)؁D�͈�K�$�4���٥�Φ�L2���ױb��Jx���K;�''�M�������������?����ט]^@0ZU�d���, K�+�_b�������&"�*=׺%��5�����b� ŉJ���x*|_��#-�_������^<�O����o�������g0-Yт��Y1���P�$wx���]�A���i��)�����J�+����~7�}�+x����o�$�%���cXYY�cX*Nb��'�������qz����]\YF}Y��ϻj8ph?��̌��z�!GZ��5l���y�_�--b�5�����1�"@�f�*C�k�~�L�+ѪB��H�9�nb�7�E6ݧ~�>h�.w�x���`�bm���F	�n���T�I��s��t�߳��F�w�NzV꺗�5lF�e�b���E=]��$��6�QbWA̰?W'�6S�fH@ �f]|Q��b\l�2"� (jA^�n�4�	9`/�~����	����ɤ��*Z
]�7[[������Db���F�2���Yi#d�+� *��07_\�(q��}��q�1#���Φk���i�+�KG�h/:.���B�Kr�.��^R{Dg/va@u��-�_O��65�B�c议jb����+A�Z���n*�a]m��!����@��+��hCS#��$��mf�yz��]X��g�|y~9�m��4FS�~f�D˾ n���I��dT^ͷ*l�W����ڡd�L�u
��t�FT�}�7%�w���,H�)�$��پ�t�yv�Pe�����fa�L��l�Q+5��5	\&d�迩O������2Jz�'k��9�Çj��|�K,���X;2'�p,��n�@�xuS�
�U�įV�+8xpr+]<�$�/� ��۾x�������F3�s;C�Eis�ՠ{�]XD�^ǧ~�Wq�G~��~/������ϣ�K]	�uxj@�4M�C�$p@o��u�>�. +���ّ��l ��J��$�%�K�'�������S�z��~aj�|���t���+WP�IeOg�	�X6��!����f��gM�ﴀ�}X��8U��h�t����&�i������E.K7ڊ�0�V6�?�`x'*���0,��.�hxJ�m[cZ.��q����;shˇ/������᧞T��/~�}��4+]PU�X��&Y�c��mX�3%6Ԑ��1�X����<�dm�t�ы����(!}[4f�u��fϟ�7��Oq��!���g���o����Tɸ6����(/�P���D<�q �Iz�bko�� NC�v�y:�%���Sg�Ʊ�K�,A����0v�A��E�.���e���Xx�X,Wq�Ss�gQY�K��T�([Q�������*��$v�R.:L:u�@S�H�tN���@�4*�=P�Z����51����RF�b9��=*E�o�FW��U�V�O��e���$���(�m7v�]�����L��L7z�Q��x�������X��ƵA�����0�&� _	�����K��F6��U��#J\ ���_��溩hи���/Q][/���Y5<�� ۷F��w 櫯���%Y�P1m%"v �)���9~��	�Z�jQ6-��ZYjc�>�b;�r�jy;�R���=��ò�s�ɬ^����'��}k�hR��+u�@��(��L9���pR�b�!t��%�R���&E�Gؓ}ا�����?q@��o#���Q�*���Yo���u�{V2�WMB�D򼱱���=U0ټ[~/�/&m��"d��po0���k���m��T'wơ	�+�[��{l$2����#�`��Ŭ�(�"Y��J�4�ԓ�sxz��^2�z�����`���A2E'��ΙXkb�8�·B;Q@�A%Մln����J��Jg`���97�}�ۻ�-�� p��E\<{E��J�c���U"�^.�f��(&��b���hV�-�BHVh��DM#+�G~�js�/�K� =c/U.FdD����[uY���v��Cx�O��z寿��+�Ҿ��^Fq��m-u#ɞ�m�Ȼ���i�8v�^�^�y��B&�A���LY�u	���*��y幭��#��g_ģ�ދG�������/}E	����Ǩr�i� ���RYlrZ��?���2��%�����EPmP�������+����~��A�0�Sx�������Uȕt�+��x��2�C�M�x��hsJ��?����o��~>ı�"��b�'FQ����|3�������=�ΝG���żr#I8�.���eV�e6�K��y}m'� �� �tlZ�e�(F��,�-%��B�e9� ��!���Q��?�����~�_��x�'>���Sx��ߐ ���|�y���KUA�|�6$3>$`�S>@Ae;���Ū��������h����$>�s?��ď��k��]�3�]�݃}�(F������w���ӓ��ژ_��*�ȹJ��ݵ�b}�wm����<��r�8IE�e��j�ϴSS����ݜ��:A�#���5��'&�['f�d�Y�q̸����j��HWz�ǘ�H�t�p@�4t!��1���=�8���-�U����v�cu$�ї�f��7Q^:�1��	����J�U�(Nm�f��U��V,�P�I�W��#w�e$;�+��4�(�N��Q��	�|@\	����݂�P��~�h2a8-	�y4V���&��������eS�������
���p�=Q�<�vaE��>N�^������Ef��&aL~;l���KO���+��"��V�Xsټb��+��m��M��٩����V�Ղ�zl��*2��I=9�ž$bM���H	��FXi�S[��=O�\ &��H�� ��ؙP�=�m9�N�{9�� K�x�ܳ�v�a��}�Ք@9��W"��\�@ �ӽ3`�n<&�$ac�\��q-����3
`�>�tʗ l�ӧi���3t��oH4���Ȼ
�����I�ÚJq�=oh�9�ݞ��b���fui+�D�{��OXW��;�ժ�%�cM|iڬ�r����Ț�=���T���]If3��L)�Z��yu�'�T0,ЋuM�6rf���>|�3�L�`�O�.��*N�x�{wa�UUV�c�����/g��l,�x��$&v ��t3ܳ��*���,��E����¤����ʊ.����!
TuYm��7�����p����v}�H/��(Ư��%x�tOrr����t�AK��N�۠��9�82�����j�i�+l��4��T�nZ�e�F[	WY)i����j�na� )��J��qz���V>��T���&�YK����*�v��K�K�Kxe�":{g�̥����x��'�8{g���h�<�st�#EIΑG�3��6��b�o��xi��� ��ti̫5�:��>�f����c�1+��nf����}R:��!���:fr��T+��%��5q�;�ķ��(>���]�^>�
ҵդ�1;ve���(ʑb�D~0��=2[�=���y=-���S����[9�@�������=#k����:���Q�ُ��VVtܿ33�f/�$���_"��$2����AO^gS�;�����c
�|�A/�2yDb��&�O�7=˵N#�_�3�u�KlI����*�ʸ��}�pTҢb�:d(��V�^p�rI�����8���AQ��qK��@�bO��rSL`�EgE�"�`T4R�+$y��_W�N3�ۛ�TCa%�s�$��ay&��5Wf���q�Qp(��?[~�tLf=��t!RA�}�Dʺq��WU�9��&3��
%-��|���F>�Z�򼚒aW��\JޮI0�5[�d{���bX�&�qAޣ�e��fr����)K���ɦJ��m��Y`OX@-�+�l���Ӛ�r ��xq�&$ݞ�zFE
�RG$�`e��e����� �&X-� ���;�Ml]�/��H��%�H�J�3�H��\�)^��Z�l���n�T0��(TdͻʯV�T���9��0��<��w����eO��#hϮboiL�͚���}vA=cy�q��X�H]}�:a9�Px9q\$��� �"6��?�b`F)@��V+R�79>5<�vLF��)�'?tm��wV�(,��)L _*i���!���ڑr 򹱺i4`y����K��bq�G%ir���nm=4Ha�d@5���mԋ����Z�y�3��������rh
!A������y�mB9��=�}���O'��mL�om�~���:��S��ش:����"��T��vC��DmY5������_�6:��.qa�:����/��܏�g��������8��}��@�����1v�C�Ih	�Zr^�z~�#��{߅Η��+����΋(`Y>;5�	����V�.��V�D;�D�-Iޒ��X~g]�	��-�}Ԓ�/���s���%[�cD��޴v*������*J�ku���kWE�Wq��o�g?���x��I\��/J�dtfb�K��P�0�=�;��LN�}mqY�P�O��C{�A&��&�5��a ܑ=����y�`.׳N!@�����X�X�` $h�U-ϵ`�����e�ZW�3��+'��<���=���Jf�,b���zu�VO���;���+�WrB��)g�lb5Zd�o�pN2�9y(����;r?>��Gq����O`tf(z?}��sǏc��Y�y�(~���ʟ_C����S*=�bÉ?P��pP�
��W��ݿ�*y���s�.�����5h����:�$��h����V��fS�bD��
�.i;�@l-5��Y�c�#����
��=� H���<���N��a��۰,���܂�����Q:+x�+�b ��T�t8�ܥ�8z�<fg0�o?�۾�wv�b4ܑ�O#�(&����U�.Y�C�����n�S��-R�؎��@Ni:=�(��J��������������b�Vd=:�����15�Pn��uI����v�Zs�Ά�r�*xz6n�J�8���K�2r#U$�<ZRlZ�|��bH`Sctt�U���d��I񨛦�3�P�O�+
������>	sCkI�� �k���ɲό�P��L8 s��o2p^��v�&9�J��U-HoHB���k�7�,���A����\�w#k��� 4)�=�~'urO|?⎃�V�4�s|cJ��k��s5a.��(X:��=�`.�U�Bpd�PX�׷���/Ηθ+�c��И�&n<W�5�mv7k1	�]p��2�}��׌�*ѐ�]�`�ⓡ�B{�������qZ�ɣ�gƉVJ����%�Jr�
�Niƍ�j4�;0�^��ҶZFR�y�B*A��﬒�ki��!�^��%jEtઔ<����	��<}��J�[+��V�b�&�H�!RE��^#Vj�����[[p]�U�#�(��+�Î���zYG¦P6������Jb����g��^ժ'[���0kkk���{�F*(�� �sB|��1M�V�u��!E��Q�׽�����$&��q��{`�@+��>ZM��v�uL�A[��އp�SO��x��Ϣu���[�H�],V^5�I�He��Z����4��O�q ����b|���\A��g/���cx�o�9;��q�~�ګ�R��Z����cn}݆�R���z����׿�<qߝ���Ǳ��W%H��Q\�#��3�L����T�	�k�3Y<�Y۷��1O�Y��&Uߐ����~��l�>���h�N5��@GY��Bf��C5.5���ʷ�RIA%#��9+sP��/c|�A�q�]:I�p�?}J޿�`|T'�8��kӒ��2YS���S�����k� ������ǟP{1�9�qQ�Ξs	wK y����������_���җp�'�]�Ҁ%5��lra�;������p��+x�G���G��~ A�
��܏d�o6�03F�<�a� ����!���J�����d��Z��W���uq�
��'�K�#�ߍ}�'5���36���?��˳��z�"N��&VWVq��Y�^9�ؼKWZ����}�������ὥ�g�3(x���y�TC"�P.iC��{d�h5�?���j�ELPHoA/�t�A^毆�Y9�Ĉ�Vg�U9mK�4ق�!e�<�R"�s�b}�\�]u>�ko�+p�U�I7���"HQ�"�L(&'4�*�ѥ�����bxy&<��C��[��V�<U+`%P����0�"����
���s�������b[t�@�`�2OCp��LcP!}���(�iQ�G�~Ʃi5���o$۽�ʤ:���%[6��t-�>�_`�[E��x��20p�Q�d�dvƋ��OH_��� ���$YvQ�c0ѧ��r��jw5X`š'v1CTQ�xO��"N�"�]�Da&c�+�v�����l���kx��0�$Nv0=���<&�By�������~��Jj�6<R�R��<�����%�����t�U��uӮ�_����y����4.K�<�a�3�0O�����$�"�M���-��)�\��h�{d6�#�Z~��+��v�2���5���IR)G G��e,I��S0�Y;���t\����@�W��|�G�{��ա�g;xY�@Ni_B4��6��}Ɂ���/af�&��X�q��Ê<�LZ�v.=W���,ĸIV��=�)HL�u�~�*��ޯ"���m(�s��������,�5�BY�7mg�h�����V��'$x��'�����;?�~L�C֛�4_��L�=4W���~_���_��_�����#�����쟦�[�t�G�g���ޕR	{$ȿ���\���{Q���I�wH�m�Rŕ�%tZm�ǔ�˹�>�#��0�m���kKY��p���S�@�7���GC@l��*�U( ���,��� ��ɐ����J�-`if�:������L�%�X�}���O��=�<��(k�>����@WFN�%N�)���l(�5W���+�c�0-��W������o(�R�w��<A���[���=ˤ���|�C���a��>|�w�P���8X�!�|�0t�@���ZL�������W^��?�N�}�!�4�/i�ëWq�#��z�iQ6b��U1H9᪁rE�?}k�g���.�wy~��N��$k[��lw�C�kO�<�I���}�%�k��~��g������ŉ3g�`�(z!�K�H4ʥ�6'5E�v�U*�͚g��L��R��0s��c�I����7砎O[*V��^3k��~*J`H�J��r��sR�k�[.U�^���"k����b:����A$:g:1R�[}b��k�ڑ�yX�aC=��?=���z;&���������2�@�}s՝�D������s�F��55��*�q�mnA�L4�C#�]�tE�]K���r@zC�8��/R��~��;M��`[�bs��j9�e����9�͖,�63xV�	�g�U�-z�2J����X���9�JJ�I������$�(!,�����+�<��l��K��&ԆA�f�Sj�����X>CW>K�����?b��pTPڢ���ye�j�}�Z�_�ܘ�o���+ʿ籫C|21yL>b���V�T�L�5�������J��ֱ�`Wlmhb���^o8$+L�c�=qˮ8?r��%X��So�Vl�۾��,5���Ėр��nh��-��
�Ð3��?�A3�%�C�9�=V���V�,h0W�Ò�Zb�7s
5�=k;=�uRx����Ԕi��$A��8u�eLO����S�m*�LMM���}�Qr+��cedDy��b맧jh�3���e��_�!��/j�7��Sj/�3+���y:peÝ�R܄*����r>��/G��Z�h��07��3P;� �$�kԏ�4�r� ��˟�ӟ�Y�&�:�Sуq.��>�pt�K����_����{��ß����O"�xsg΋�1"1G+�`bbTu�I�6!��س�a���»�}{��+�=��`�^���Ә�<��ZC}!�ut��)P��<�.V�&��4i��*��b��0yܐ�校fДD���DM�wf��U��z�Iϵ�v�~�f������*d����3��T�\�G����U��:?���&V�8���e�l5a�~ ޓV�X��{Ztpja�3{�/�����~棊ɖ#�8 3f�&��J��>���D^7�?�w����fB1����᯷�r�y	v#�~-�p���8~�4�<�$��u7N�����r�PX]�bd��b>jđ�v �w���فl��,kQ�S+��S�8ɵs��	80���+x��1��?!�{�\���|�^<�s'O��S����'���W_�첯�/�R�D�z�˴
w������&Gaxv����Rgғ@�*���.��˯ɣ��%6�8���7�r�S���$:)�tr�j��Vҍm��풽��"��������se���eʋ@�تTy7ؠ�7���N����O�؂�>�~�ųr.#'7�S*����߮��It9�E���h晤Y��w���z���L������M�B9��R�������W�l���\�XRB �s�C��� �)Y{��|�N�w�'���o�7VY��ڒ��$=R�����V����u�J� U�g<�� ��n�7�ʝ,HU:(�*;��7�s5@��jU�.���p�6S8�΍_I-a ��3���#�%�a���3�T� ��k�n�b�ԝg�"֫M�;RG�6���l5s##_ל+{���0YG�^F���ZV���XĖڈ=U�<m�g�O��#bE"'Ae������GL`��b�x����#��6�6��a|�7�ߎ<+���<����o�J{���\�]�
/�G���T�8H�ȋ�mZ�f��[�
�����G0�Tt�$[W};?�N2ȉ~��ML��.�O��y��^�uʩD�@	�#U#�.��x�싒�-���˧�u''wᎃņ%�oi��gfw�u�bª�
�qՕ���ۊ�ԧ1y�"~\WE��y�-��"�y����t0����b�<�4�1�tG!�	���>�8:W�p鍓(1!�ѐ@���c����(L��X����0>�k�����?�a!&�.h-$�J֎d��;䟓s����2J��ÿ���_��z�1���ђϐKBTj%M$ ��=]�_.�ݿr��hc�]w��w��f1��@i׸V�Y9-�/a��v%rpB[��)a�PQ\��[S����.�P��J�|��P*��ή��b�2c��2Bk���S����n�RApz��B�ZGi�(W̰xnZ�2Vk�z�&ר��	��	L�>�Ru\qes'N�;?��(!b�f�©ihҼUFjXO�8s�2V�u�������}JU�V�P�Fj���z6E�X�d`Fp�]�p�����گa��,����%K��a��+I�nu�\Z���q�ɟ��{��Ȯ]��K�r���fi<LP�F惨�:�)�#�O_�`�����S�[��r��#���|���ĳ���:���5�>~�ldYօ���ǎ��Nk�ƪ������k��8X�qw�X��`Q>r������qZ����T�z*`��t�'�(!��	��1|&no%�jl�
��4���E�Z�!�j�����dxͳ��ci�Q���u���= ���s��Lt#p�+pZ����]�N��*/��a	RG�̆��S��IT�)�R��,�����>��.ܐ����ӝz��ŭ�؞iD���If��ᄈ��s�;=��]��z[h2�ȘvD�3q�J�'��7�{�����%ZX�1�F<���<u�*��I�E%@/��|yN�CRf�┋��U0oqe�nl��$���Z�2!v���'�jj2�覀!m�5B�␆�"�*���n��_?�d���b�aBr��dx7ς�D�o�@�z���t(:hr��	�}=�I��)��C�6�ɪ�c��!YG�FǂI��$]���|O��~C���j��/]�w5�Km%H�� �H%��g�w%�����[\�����M�+wf`\�6�n(�l^k�b�:ɺv��v��sw(��W�Lvj̴��s&[�T-"�*���èU����nG'D�lB�ɍ�.��5�L��o&5�gиc��\|�My/����S;^���Y9�J��]�9<�Ѓ�����������w%p�_���bLHB��M97s��q|���+<��_P?C����o:͙�����do��xx��?����~/�:���uKr�֛k(H_��3,��!k���$۫ǎc��A�"F�����XY]E�VA��]�/�PG�~xN#R�e�DD��uBK�I�N��ď���T0�{^��?��%�iTY�Ss�a'v�|g��o�Y�����Se�H0R�K�������ǖC�N���8�rQ�gv��b��Oc��%٘	��JTȖ3VVx8����mH�����O���*9�VKJr<4���W������f�d�������3��i�P��3?�>�L����D�%\هﳽH��Ξ�M����}GP� o���텶�߹��S�3{G��Җ�]6l�d�<�%٤�>�.���I��91�/���G��8�s�O`naElGk���t
�ScX\\���9����gU���'�����~S��5{�X���\Np����̮:�J�1v�{O����ntgv!Y��&��g�2�7O��ƺ\f��M��|�	�_�Ȝ���M�2���84s
�̾Nd�w7;��ߕaD�����P�h���/�Ğ⧮ulkm!g�^6t��l7݂�:��;)E|{��GI~W�W�U,L����+��
��A���Ɖ���,r���2�]
qp��nɐ�������R(�1'�j�l�HIx�juY�#���|7�C>s=r\JrBSB78�2��	���7{玟T	��$���x��Ұ*�&�~�qf[�oe��X.>O�����o���V��K�@���Sl��$pҕ���8+Q4�S&H��I�M|W��A�9��9w��*u���{�&�S�4�w���"Rk�r4��h*'砬lA��ĝ?��.����s��ڔ�5bjk�[%���i�b��ʋ��o������w�S%d`B�
���&?#!t�&_r�8�J�`��m�vȊ3����ig����wtY���gԖbN�ޭ%�m�q�Q�q�e�bvI
F��c�s�%�q�0]u���}��V�huGpq.Q���h�?�8~������]SxR�Z������Ok���,�
��?N�K(S��v
��-5�C�'�Q�L��G�w�c?�R�{k���q���9����� u�AW�g&����A�8��6b	����q�'J��2�-I:��>PbN�t��b%h��'Nѓ=u�SO�_�O�~�~�V���:I�IvVtk##讬�uё3�|�Ο=��G¾}��:���>VE��W}\6L��%*��*=���F� v�l�V�Y���D���8y���FV�o`� <Y�*H��U��[��.C�u&�k�fߦ��^�ᙘ;��Z�撚�l����ْ�x �OWsUN�����NLF�|��!P^���,�V�M�NM���?��^	"��q�����Fz��ӵ�9(F�����#��g~�ǩ�X���U�(�J���ʎV*9M���Z[�`s���ʲH_٠�}�݃=G�ty\�h*|�]�n�`mqs��!'�n�0�%'�������r�/�ş���ａ�K��|�;0����_8�#߅���i�w�^���w`��A�hE4��r����\:7�ŅYm#m�N�uN7�w�R�{��?1���S�]٤��i�Z��s�kp��FG��h��m��hx�M�u$3�IF%�y��QlN~kF��?;��g��y^�J��z����$�H��į8��db���q]�3�ͥU ���b�Y��0_��@�%��<�C��;��ʝ�V���?���؊ͥ#Tٞ�MްST��(�����Y軀g;$�õ����:���&$���b��O�����U���&����"��r�q����ڌ�HP����vJު���R������3����JX�䍪���\�}��|O��KrW(j����/��+���v��6)�Kt��tE���96�M4;I���:Bޟd�t�L79E��3a>��+h��s#%Kre�*�U<#�b�q#:V��2#�W����n�LZ(9%��qA\=(�p=1zT�1zo���D䵇�A���9�Ĝ�ܐDY�/ݰ�Y��rڝ���\�5V��S�QnY>�8nꀅF<�Ih�HՊ|�]Q/��UlC���P�J:�����t{67;gq6�Z���j! @���:}��Z����g�dŇv{&%������ƴ��I��a��@�(Hj�����R=���(�8q�$����h��19=�Н�{fp��Yݧ{���=X\ni�1�_�$m�ʁ�(8���	�<��'��1G�Yd�l��/�ՋAL�\�����<��K���D��F�*�b��\t�~��܍�>������$���vD<�_zo�{�վڠB\���I�4�OВ�����,�,�FR��A4���F��-�]f���m��>7��ˬ��.�g��HTV���"n�{�>��B=9��M�bm]�)�֊}\���A��G��r6�f<����?=����Oo߆L�_[�ҙ_ZZAF�qv|W	�f��ʹ���;vߑg�E)� ��UP��}F�X޶����ص��+hd:8;<�D�t�º��^k&�}斅�	xw��G��&
�i���U!�ґiaeV�[[�YH�L7��TM��4�n+O�ix
���dD���JC�G+���D��y�`9W^�ĔwH����e�*c��iů\�CO=���>��51���������>�����Ԡ�ճq�{��s?YYhrFh>���>uw�L�p��RQ*׏�-2�E1��U�/Ձ��/|I�><}��>BQ6r�^D;iaQ�-_ ��޻�U�Ew���#G��e�����/#�Fq�$��J����Ď�;��R���Jd�FK�wm�!C[��h|�I���ykͻ,��{ ���A�B��J�U9�����)(�V4MQmꄹV��捣��V��b�3i��jͯ�������M��IYɧ�?�G�xqi1��vS��~�p��5����
���;�H�섾�kB�ܜ��l) S��JO�7%�%�+�{j<BA��-���d�N@AB�L���X�k�._@���a4s!�z�N�a��Woɡ��ZA����_`��c���
�J�n~��J�4�dd��H�h=�)�����$����d/OE��Kԓ�j+�N�H�15�c'ɚ��+����8�1�i�Q�6pO���(J�
n�Z�d2�)1~+6M�Â��]�ȗm�3���,��6�?�)��VJu��S�K:��[���-1��b$��z�j���P�{F_�d��
���ĵDQ\J>�����YfcI���M^ӵM�Q����Q�sk�PK�b��UY��aD{��a�X���f��G0��f�}A���	fl�D���mV�
8e��d8� �eQ��&N��}7�XZ+|�zj2���(^�QD[�*�CH>����tv�iD��LPwUx�PT�Kqc��T����#�e KIRq��-u�){A=T��p�4�ګ�V�vB�Z�VI�R%qH�����^)��JgjEԙ��u���iZoVޭG� �QB�T�Jay߶�%Y<�s��8�!#�ݨ"fj."Ε옰���Z��p�������p�)��ѳu���wk!W���������G�L �8���.�~D+Z_�ُ�ӛ��yLOO���㚦���af�*f�����GK;����xϐ�
=���2��U	beO�#�DκW�h&��T�K������h��1{�<≸<;�礥heD�Җ��|��K�2~�����#j+��4�o7��F�77 |���,;b.F**94��~����~�:�6<��y� ��W-We����)-l����[c]Ah��L/���r���5��5$RID�S-M��JqQ��H������m�Q���TK-$bR&���a�aܜϛY�u ϔ�3e�By����v����N��j*YS����݇��ay���Zo�xoK�s2�R�\�4�g'L�BV�F���*]'߳9:U�����3Yl�������{"�Y��}��aL�ه���2��ۆW�ë&ƻTV�[�h�U�ťD�_�r˂쏿{��ALL�����s0��0���#���z��?��@o_Ν�����mہ����#T»o����<�̳h�M��3g�`|l�5��'����r�VDg�a��a"q�Z�Y�@.� ǆUW.���L�~)����l �XX��L%Xr0%�ڒ_\0|7^�Y�l����� �����2=X �JY��Z~z_{��K�Z�\nG��Ӄ��89f�:F�F~�N��zU��!|J�{�O�U��!�|�*�����ns�ayvWodWs��$dܪVu0�
�L^��2TB�a�E$���L&�bYY�KŢX���6Yw�d~J��8-6�B)�P,Ik���dK:G�v�5�҈Gz@�a���M�n]�ڶ�{Q��sx�O�T#N��V�/
���;�{;���ӈ�z�(6����x�"*�gU\��2���oM@�P��U����^�ܴ_k����w�7��������\�b�b:׭T,C����\S���䌬�b���G�e5%�(���d):����܋�U���yF�.�k�J�d���0��2il�1����;���G{/����LZ�tL�ݼ��N#�LPɽс`�e�l�D�D|-b���O#�m��Q9���
�04�>ԩuG�Wc��2n�=#̡Nl�"ݦ�T�/���B~������m�j�i5�GUVrz<h��F�PN���Yld� GΒ=Գ�^���2NZ�+r�e�&��6�8�d�8k��#���s3��ؽs�Fe�8H�Ӛ�����'+��9�鹭��5$�9�].���$ԡ}C�-S��/֊U�Ĩv�0�e�\X�zM�s�"���������6UB�g��m
��ʙ8�����ŮB���[[���;�>`���'�����T�}�5��_�3��!��GܥfO�Ɓ�E�`|�vTĆ�Vo��Ե������ӳmq�ZO������Qi+�$��L�Wm`��r<m�t���MvK'\.=�X�UC��ܹg�|]�/�0������T�F�<k�����mң��m��s��Pm�$�bts����U��ƹ�*��űB�t�Ȧ�>���"�2�8���y��-A�����ٻN����q!���	|�e�d!��*����4l���b�o�@_���O�ʩ�xz������a~lS��uS=���&��ߎ`hdX�QSӮ��6v�y��������_�l.�g�=��?���F�㉘k�e��e�u#���Pӫ'�����f#�.�}i��C��F����jm�$� �m��WA@g� �%��C��iD�u���^oo���JR�O;`���>�'�Q95+'�5�����BBt�d�.m-��I�lx�9RIv���u�JT�'L#S��wP����{��/_>�b5u=XMG<F���M4�2���.ǯ �4���\Եr�.�]۴~[�h��� �RS�#'僉;S�ld*(�BnH< %��N1�:�Gr��۸J�����o�W�ڕ�w���[�D�X�$v�@=�nb[� ��C��ݾ���\�L}�9���{	7 �z4�j,�
X�9�m�
� X����`�U��R'���XYA�"��T�ʒp��dѿ,�+����eVBI�~l%��v��D8մ�|� ��>��[EMQ����k�%mRf�b�T�9����D%C(�Rf����M��'%2��k�#ס!h[�	���M��ѧ�W1Z�k͈j{1E�����7b�}�6����)�q�=�
Xp(���V��	 d`��c�������jNn��Ȅ3��a��%�6S�u�tcک��UPz��V���~c=����[��5ҫ�/������O�Դ�9�rKQ��ݨ3�,�%�� v�����E�xM�+#1F5b�����93�y$\�7Qͥ�:�,�9kg�ݚ\�7��s�9�/�M\����0~��*
���oU��}=���5,-�
N7����4#Kh�B�j�nܻDU�hy���`��5��7��B���4Gi�
����=���U���}�����ˏ26�⎼Qq*v�؆���h�R�/U�=ܔ���pܩ�dLp��];q��W1�ۣ�7t��k"ùd
֪�n9GW��@R��9�-�w6��;]XZ�K��Z��%W�v��i��'�
;�isn�[{s�T�������$���s�T�����L�B2�����v�gX�~��V#��/Jl0�Ÿ"��pL��Uː����������d=�}<��&/�d��>���gE ����p��X��7TlU^q�~5uQ�6S1~�\��l�B|���Bf�A��h��6�?<����x�Y��n�%Ƣ	,-����cq���>>���]����/q��e9��.^��H?�l����++���q��e�;uN�ݨ��@��yM$����ٕO�K%��ŋi�V)�\Y/�(�W��h��A�4�i�ZG2�0=�����.�����'���^?�F`b#��]�rY ���pAz&=�n�kA.r��u���A;�dn��$�M.�\;�5�Ak:�,�m�j�����?i3�w|�Ns���+*z�M�:���Xz�S��jQr�'2b�W���ΉQ���&���cc�8�� +rϪ�W�vU�� ��gp4D-�Z��R�T��'a�̙%���(u�`��t���,2a��g*��b�	��bH'�P�Ɖ��z�-��(��(�^�2{��:��+(���5?���bs���I(����Mo���zAʷ�:��h��el��}qM�0��)��9�G%FU��E}��FE#�����8��}�*B+^?S��p����ȴ�p��@~�ў�-�s�a~ji�'��#!��P�j�:��$����n���[�2�`���0e?\�󕴜�E�]qL,�k��	pY���ྜྷ��"Y+j��;Q+9�Z	�Uu-MY�e��&b�#(�b�,Hn8��c�B�f�Xj���Qhon� m�q�=�4Tdm.�ĩ�=��^��s�ʧC�����P}���qOe�)8�[����U���JE�;v�	i�EN\�/�Zj���8��~-ܪ�<��� �
��SReЄ�^tp�QG[
�8Fd�-�pU�i2�R�Wo0 Q���ӫ��/I%s�T]9��(7
��^Ɔ��C*�� ���l�8Ǜ�׮�	��,;B4+�2�ٖ�,���3��X��,�o��U^H[q0�����Z~0��\�Q������_S�V���d�g�)���e&�)�W�Z��"�ZS���Ŭ5�H�)��S[��FT��2�P�Y���0��m�֭2#��;**��>]�&��d�H��e+/J;Q���'Z�**T����ב���IUن��s�\����Z~4�m���Sԕ֕�.-,�\���>��T�Db)� �t��K ��b�w9�k�|�e������JI�Db<ˈ���:4҉�F����ZC�^Cێ�T����|� ���V��זQ�%У��ؽ�{�C˾剮*�t���G�k�^|��i|��oc����z��7d�ػO91%��U]i)I���ݭ�� 5id��Zc.�f�g��;w�y���� l����bgC
�g�gM�vːl��]�,]����'t
H�Y���4���Ԙ�_��gn�hͿ�������ɢ.��é�_�ͣ/V�i���,��d���ʵڝ{�����>�%�=2<�Y� �kˌ���%����V'	�vد��^���K����M�jE�s��*�6@JC��V�a(���Y��²mR�a�����=�c���R�_�#�b���Y�^Hg�L����#�`#���WTcrX�� /�2LV�W�U)f�����j�UĶ�'�0�s+줡��������vFG�v"9~i��k�&��u�uĹ�:�cm�{��F�S@ ��57���c��η��"`4,��b(�K��C� ���N�RQ�\![�Y���%6���Ķ��9�br���1�]a�F 9�h�
_���r���d�$�k�ѽ��'���t=��Z��U�`�'��G�X&���I,�M�Ɖs��@.!6J��R;(fd��Y��I,�EX�Ж�F��r�C)���o���E��U���nMG�hNjDĿjL���ZS#(d�H����Jk_Z�gXr�t�)c���.%!���B�8�ί��hg1��`4��E���RZ��ݷk������"k+k�O'`*u`+"����P@uiY3E��U��8��mVg?a���UĽ2�de/V�'\��G�a��c~�q ����}7C��2�|;vL+O�����X�p����H&��e4�I:��h$��˙�Om���i�.��� ��Zikh�N��!�U�\�ߩ�i:b9���ۂf3����3��˹�Esq�MI��r�L?�x��]�m?j۹�{���3�����q[E��鴡&�s������r,�$�ؗ��!G��P�>VĴP�ZS�bȧ�#��~�m�H����ھ�51�M�D�g+zk��&���,�p�CGo/d*���i��:��/V���V-�g���	�:>/8�M�
i{��+���8���(D�~cpW{=�0炠�̇MBiU>����R�dU=�'���(��޹�22ʡ<;��q$�ys�,�i�K�5m�h��;�]�>��o��	�X��x���x�����~��V�R�7��W�5�A9���2���]5��CM��̓�y���b�C/% /.�X(k�or8T葢���͡C��УGѷw,޺x�a�|�*������]#CA�m;|�Z�K�,AS�32) �/o@�v7���wG�����eCvA�Ŷxس�$�e�B1�͒x�MG��6�{-,���=�R�u6&�E|�]L���tU>��MF���?�vN�r}J+,�|s)��r �A
[��Qà�@ԗj�1P�6�T�AM��]H�"�QSȦʽm�s�ͬU�n6��ŞI�_�~�0>C����$�0��b��p� ��x�����BF7�3�fc��Y�P��b˾=pF��Vl�o�γ����\��SF2��ܡ�G�'!k��*��������K�����sv��^�RMqpz�9q��x�3���G���&�B�T�5�j3��Qtb3��{���p��9�$����ke��H\S0R'�9:J2��Lrf�vl�i��A�UEm����e�����U�v�.ںl*��.���̌���߃h��ܐ:X��u$P�jZ��r�Xx�k�dG&��c�ڿ� ��zɰ8V�-��nЂ�kh���z��z׬^�����i=~�R��y-��.���܎��DX�B9��W�0J%sRDt�VL>��y܎-��c��W巸�M%{H�߂�cG0w�:�W�#W��)QM�ʪ:Za��X��V+��F�0����ڗ�=;:Q3'���u(gɘ�Fj�zO|xF���z�_(+�.@O.�EKԗk�r���/�gbj���G��8�KK�P(��G�j�ZU=�4�*[FC�]�Tb�[+N#�2�>`��aP�_辞,�_8�b��p<�ł�ՒF����U��xkT�{�x_�Q���GtH,M�?������4�,�봫�������SUL������y��b�REt�� q�O��t�&���|*k'�x�z�����X���3��D�N��� ��<��K�g�lm_Rc>�܉z��������j�ib9�ϧ�`��Y�D,�ۉ�:2������\�L<��)
'�g���y����A+����Kh��gU�n��h'�����b٤��K�`[ZX��(P\�B�-�Z��<��߾"�i�h� ă���zH�1~�W��#���7�+f0{�:Ri��D�vEK͋�:FǇ���-ή���q��a9SX^Y���l�eLN�77=��\ܡ���g ���s�����^BK�fH�z]vS��j-�H��Z���}>� ��(�&eɿ	؋��!*ƱE�-�#f;w��N*�3E�B��"f9y{�=�k?�	�gg+�YY�ZV���u#2m�Tc,>=a��~-n���)]e$-��K~�.�KcZ�ei�o��LE8q(�<#����s(B���-O)�Z59=�bУ[�c˗^lQ�����۝ym�(XQiA�vz#;w���I*��Fw�N
��NC�dd�ﶍd
	�4jl���D�ܽ#�&��j��n�d�ic�Ī��ɸ�Gvn�C����M��m'*NW���]^��:��._Z����J-4(&+�W���aޱ/�����}i�ۇW����֖o>-@~�&ku��A\<9�bq��,bU�y<�"F��i׶�,�4FI�fWq~�v���c�=��C)��9@�ڬ�VM8G���BA;�`ЖѦ��Y|����(��n�n�y���ܢV𱠴�Ë�廊��K^����8@1q��L/>'�}?M�21�Ȋ -�K�^it$�t~|���y��	{�:��h��8�e�N�ɞzW�-`i��DiI@�����@�`�^B �D��/�+/��<"����#6��8?w{V�E�51�U���{`]_�Uq�"�`��j"l/�:o�'�e�ũ��!ϰ��bn"���Ķ�vneX�8N�}��u��L�j�2߇�l��DU�|y^��xd�0r�ye�=��ЁO%kh	���BJ�ݩ���o%T��A��/��@�t�ݡ��t�	~Zu��;%-�j#�M��$�L�؊��(�M�9�t�)4Mq���c��75�w�B�ʊd
��>��ߓ�^d[�jTY�@���,��a����ߩ��k
�Q0Y+���e3
��"����t��LvQ)f�<�r΃o�q��03�:�
c�[{���t5���bn�kL]�2�$?]ළq��?'#�v>�aU&nqf�e�b�{�Z���g,c��j;���7��5�+X]�C]&?�׃ۂ$�O7n��u!�C��]��\���Q�T���S���G�\TkT��-�2e*�fih� ����bFes��P)��!@����ֿ�W�#��p��t,�����+r�������C�T�T@aiW�]cÕ+���[o�����P-�*g�J�^r��oe�ه�C�1{��;�;�Z����}-FJ�ؾҿ��Y[�����?��c��T�<|�$���:*����٧�X��u� ����eqb�1��$�����/z�̑��5�L��o ����%�
�LY�K��N���*���Eﯾ����X��y8�&�FM�-[��5 	�:�IF�M/�F2�z,�Ԏ}������dc�X�jt��ڟ����2��۩X�lL	8��2�қ!�._���g��P]欩)$�A��-MiS�=Ψlʜ�) ��ӈ?vXw���3��v���0y����g�z�����ϥ00ܣ^ۍcn��f���~V�☵Q��O�Mⓚ�K${��cO�Б�%`J�����I�{�����<�)AG�鱃{-�q�^��� #S�e���B�eү\�M-���,Ѩ��ÿ�%d�>�j.,Ϡ�� j����\�V��hZ��z�����Z�M9=�i-FFkq��ɧ��#�K�����M��Jwy�_�{6��1�s��Y@��>��C~�(�O?�F	 � �l{+l)�S�~��x�(�����k���q|�z�<��|Wš��xW>_Υ��H�œH+�����p �̋m�:�����/��V�(A��n�iݢiHg����d���L����������P�1'�_E3Fi�+Ӗ�<���nEn�Nl{�Btjb����gRָ��϶/$�szY=15%ϑ��1wM�����rvՍ$O<����ή��۱u�6ٛ���֌�����9h�҉�r��.4
58�!��]m�&q&��iՐ�ݭ0��������(br��=Ks3�DbQ�Ւ#������*5�i�l��5p�~�_W��Y��l �3蘥�T�k5äb���ɘ�tf =ӓ��*�@SK7���q�F�\ë�8B�}q}]b%�1�)�vL�����2R�6�"y����y��W�'%�$�X�)�2���՛��\먇�}���iPB]�����y`Dny~�\� ݲ��b���L��W���PC��Q�V�J�5��4�J����-- �J)�TO��M��*6??x�MS�֨��˥sgq�ÏucS�B�-9d2�)�wK��,"mn�7�R�_~'/�L��վ^D�}�aUVPxh'N���a��C�I�T ,n�ޗ�f�\S�6���Xo��&��:�LU�=��)��A�S��*�QE8j��w� Kb���<v�;����U^P�_^����+���X��a��'������E8�b�V�H�ʆ��"�eCG,#2�B�y�� �s=�>�R_�0�W�*��l�)��y��{��-��j�� &����)�%aK|)y���2br�Uлd� �L��G��,>�s����<� ��V97��wi�y]i��a"��F�[菦|!�:���o�r�ũ�w��-"'�X[0^�*o�4���"���"�eL@��{��?�h:�UjV�y��e�,�z���� +nN�ޯ���q�����܋W0&!?�b��x(������%�Z�S9T�8�.�8�܋��_1�j�օo�l�s9�hO�Pjz��L���/�wd�����ڻ`˧L6���2�w�϶�X@e���
�Z����v��Cx�'�C�s��v�u��6̏V�SB#�P�Q0�PmX��&Pa���V��*>������Qd�=(ח�Wt&�@4��V����=��_~᣻P�1���-�)`�#�;g�`!�`8尡� b:��A��N�x�TD�ئ\N�"�����b��A���q�jͤr��e7$��=6���C�7?/���P�t�[��R	MS��v{�|>�Q�fu�L��cFC1t Fo��=���9��qf>8�謀�Ղ�G}�P^��5=�Az$�U��A����-��חE	�.��ۄ[Y#������yi��=&\���g���╫�p�9�L���RQ�I�c?q �-���(�p��L��^;��W��F#S�0�%7�eǄF�^��Bq��2�l�����<��ɉC.�����d��9=�ޮk�p�����J� 8�k�e[[���u<,k�L���j�Ί��l��%9ê��s���}8�4�<:��Cxr�W&�r�]���K�1�3��hڅ5����H5z�<S!�v�>~�-lO��`��󤪱�j��ђ�!�E2��O�5:���=T���,��-u�?Lg�F{��T�F�A�(�S%=I+��*���2Ǵ�k3�G�"m�XF�Z�MӞm38�~�����M�L��m�'9��kLх_L�k�ä�\�n�ᓉ���Rl�-S��˧Nc_�	�ON�*��ƙ3(R���I&rԒi6jHg��lT�:3��~�{��7�)���
��k��~�β��T-~Ϥ_�G��S�������+�0%`�]���&I҃��K-��``dL~'����ђI�I��:����W�H©_�,��E/+�&�1�dhu�4�����6W��a+�K3.mj����zeɨ��i�:��V*�QB�j��!N��|� e�S��q�ޫn/r�AĈC�K��D�o�掟ҔT,;�h5�)'r [��F�N���-���������NP6�����
�BL��8+�&���@��k���C��3�q����(Ҳ��nUyz�s���$�sHONb��Ǒ�����
�f\�@���#��l��/�j����r5&~��rR���+(-.�a��=WU��V��&��3+�,���b����#_�2�m���Z�ڿ|�����5������⅞V��O����Q8V檎v(��쥺��f_I��ɞAo�{}�C�'�����u$inB�wB�����������A�|��#�:y�}<��^<��~�衸�T�Ջ�>��H4�� ���!�ڵC�=~v�ն��� ���%�Ӑ3���L[!����@6�����|����;;���k@i��VQ-��2B& jxt���0��#(����G��6#Z�x�����ϑ���c�������0�ǡ�����w�!4�};��?	w�������\�:P"�)ҁ�	��k2G��>�Dv���:��=X�[�_�'&z�+����0RO��}��>u�wϊ�C�7�����O1�-�ZXE��u�b����`��
��'��w��k�:m�?�h��=�/oA�?����j�p�I� �TJ��^ϖ�����M���su/��ȩ�E�_�0����n�,�Zs;�%�Z
z�,��I����.kGFs3Թ��Y�v�d#��@g����8>�J��y���l�QəVy�#�5Y����=C��yO'�$�A��w���Ν����Uݺ�<�>�����~�'��J��Z�V3��^�q9�Uo2FK�Fߎ-b���3��{�2p����6���WVM�]���L��rI[�F���n�6��r�5���r��UE`���t�4�^aH��Uu"r�ˊ[�_�b���r���"�A�"�V��璛�3�Gĕe���QܸtW.\��#qf�V���6��*r��
L7ڦ�K��P�\.��~�����Ǐat�Nر��|j�&B���F����X�Ja���^����D��{vڞ�(�
����A�܂	�̦Wõw?�7�,NZX7NZ��P}3����=\��� ��t��y4�1A��`(��wumg3�c�TZ�0��t��]�Q�
+ZJ�(�o��RJ|M	Xٱ� v�ډ��Q���j3�]{�[ō�G�����>{��1����v���A,�ă���C�N�z�!��r�<�د<L�Ю�½j��;�n�ɛU�3����1��N�y�f~�1��=�-��N̈́#��B)Fl�8z����G�:|�,숥z6w�A<�{��[�#��aOd�|Z欰���FQ�06����d�?(���C�
8�����aO���*�w�=��'����ԑ�H�`e�󯾎z���6�O͈��M���	�~�H<zXi�fY��H�֟}'��n�JHˈ��6� �w������d���$Pbʨ�QW[��Oj��X���=(��wxn1A���2��L�:�y_������!��f8�L�*���7�]V"z��4���Bt��)-�`�9e$�� �ح����x�B���zl�ԈӚþA�d��lNÒ�Ձ��U$��͜��mGn|ɉ����e&.�f�,�|��:�r�����;;&�|����f��9�,�WI�g=y�aL#��+ئ?y�5��R�5r�F��q_n����U-h�pF�,�3�������*����7~Bp�p{�v������@%�� c�h�o9���ܭɂ8��l�%g���?��&�s�ŌH;�+Ө��\Ĺw�����}�gB!��wX�%6Iĵ��є��Ǽ���^};�<�ч�#J�������tF�ߙAaU9�� ����^�8E+s�Y�DY\���"�ę](��g#=9%�v��W��2��c��ɶ{�x2��l��n\��5����{�@���Πr�t��Z4K&��!D)�[,��Vi8�{U-ׄi���Y&�ض���յ\�!�(�����G:|$����'X�
�K�x�d�������c���=�0���	�:�5�Ѩu��0o_X^FRj&'�������	RN��aa�X���ˎ���T��m)X]�z/��_�ډ��	�]\;��PD�͐��XN:����01=���<��;������c�^��ת�:k4��-�G������@Ti*��q�
����"J�Rؿo�`�X��]XX��xF�RQU�ۉ����S8|���
8	w�#���_V���h���d�F ��߷��0;���^m����$�ZP�G�6	ݪ������%��p���|}tD�OW�q$Al�b�� ���qv�Ǳr���$�#M� L���~�a&��� [�D�^�\�ݍ�4�'�z��@rK?��S���4�\��/�1w��ʡ�w�˂ZvMz����������\DA/*�mJ�o�
v=y%AbԢ	mC���:o�a��m�6T�����6)��8a�y�&*�ox����N�
�q1>1 _�j���L6!CZ��x��Fd���^��X3��M�R�p7���p���:yF��Rb��쌐H#4�F߶a�%����1��¯V�G���׮Ww�ߗ,������Y`�];�p�uee:�&��KR�vN_zz5���y���|ON*�7�C-ni[����{6]7��k{�n�(e�9��s	�8�`�f1R��+̍�}�)}�<��͆�&�����>%Iy�.|���)���,��́��J����GB��<�_0���e�|��QJ�Ь��OG���nӦx���Ws�h��z�W.aafC����fQXY@�Efb7����r�zn�+E|��ݹM��Jހs����B����j�.)�3?;�����b��e�H���F$X�{��:?߭�=cc�>�����o�t�*?Dĩk�u��9h&A����E�2�v�:��33��E��.V���<3���t�b�b�e2�ѵ�� ��v&�(Y�K遉={1���X�����1٣�ha�z�W�k��JX�C{*◓�Mxl�5MUP���pcv�;w``���p	�ZI?�QH�$i*�T�;��|���oə��W~�_ �ˢ��6��KD=(S�l��.���S�������8��0$ Ϯ�e��Q+�HDu1֙j ��0�s7���� g/�AM �c�d��b]�Qzr�&�2��^C�6sDσ՛�����������64ɶ�bj�Y�RQ���E#�#Z��i� �:!�{M)�B���]�K�Z�3��ٷMPC�'�y�cŏ��N2��6I��"b���3���Q�S�}������y
��Zy�3Z�����"s�d�?���c�1bG�t74��V`����1�N����(��'y6�'A[@%zx��WRSH7��c��K���PJ���m�$t����9��I���S�3���Ebm�3��7�W]��{4�HN`˄����˯�O���|?�R|��ϩ�:���������O��gd�X��H=3�T�B&�v�^���Ɋ[>ת8T��i#��(�C>C&�	"j�|}Y������`��|�ӊsF>56��,F��J2�48��$PwƢ[�{�h�;�Jl-_�	��.�8zF���YJ``;j)��
��=r�s)�R1u�7��ƚ~�F9��7�qT]J�tR~�b��yz�(�

�,��nכy��_�����g�:�J�_3���k�Hk��P��N�e�k��Ph�������eҔ*��5304�~9/��}�)e㒋��	��jE�u��Z����������x��'1�c��/ �t�I�Q��Qk7��'QXXAJ���������ѯ�:R��t=�8�Y]խ�<Y���vF�3�Dn��}~���_akR|v���!݃��W�]F���@"�f���`=y��TX����Y��$����/��`���Q~f<(]�}M�R�9v��l+�"����*����3Ve�lfh�=�to��C<���/��t6����2���r�	�p�F[�J���	����51S�_<�����8a����0�tN=�č�%���C�~qv=�8��}���X����kK�"�4�}��/���+�m�����=��q��|�'<t��Hh���&��;���g��^�!2r�q���r}^<��Խ��?�jZrߣ�v��Ï",H����������)����#�/.�R^��()�c/9�-y�L�r�Sj���w�p��a60#q;�����gZ�j��g���Kq��^�J�xF9�m��(����;]2%5F������յG� ]�Y�zsq?e+kJ�Z��՞�P��+�7��*4�k�o4x�΍c��6*��'ctg����rϵ���=W�� y>G[3.��6�o����k�SK�3,V�����"�Ať����t�����b5e6�:�ؚ�3�(�u?o��ϙ��h�|�q��/8>����_�������7S3~D���
����Fa7�<5�l�a��YM��q�&QB�"��S^AŹ�'䭏R�;]�T���2Miz�\����KEӖ b�1=�����v�4̓颦tQ��?��nI,�wY�u�/=����Y�׺��L�ME)��K`S'}�����j\��?O턬n��1��Z^�Ǉ－G?�9�~�~�ziF9�l�n�������Y��yf9^{�%4�<���ٌ�����k����t
�WLe2 @�3%/�������E����\^)U  ��IDATFA�KjҾd38lWZ)a�]�c}�c���]���N�.X�J؊XiK�G�?�%���1�T�� �����5�n�,ZX�O2�����OE3��Zy�\�[���%O�RA<N���M��醪 ���g�Z-�ԅTL���*Z��;C���^%	�A�#&������q�?lͫ�-s��w�ٶ[���O�2?��¢�䫧a��(5m�!���}�q���������x�s��^Yɞ4	*"k-���}U*\�|�Ξſ���̟��!Aك��ʪ��(KFQm��KS�}��x��� �׋���.�?�H[���N���6�؟��+C��'nٛ�`Xw��>�M���S7�Z��!�{������a���_2*��Pc�'`ߙut/�T}������I����ֽp��߀��ݰ�K���@������
�o֮��>��R�&�>������m\1d��GK:��8�<�C�6](̏�m�U�հX�»���5����������s���Lw͹����U�ɿ�@;/xG��4�C[�u�L	mۈ*�:� o1��7���?�OI{�g�<�����ykr�0QIFa)��i� ��?g����h����Bw|Ћ%��{�ζT�m���v^aw���U�Be�Ep2՟!_j�5�����L�l�(=Qo�5�a���s�9[�R_�h!*�_���V���H�Ʀ]m��г�bC��.к�P��=��}��~ѵ��L곷�V�k�>V�m��F�,��\�`��~n>�#�d�/.`aiY��m�����k�ʔn��}gm�M��P]Z��c��%L�݁�۱�\V\f�f�HE�rNW��979���W���-y]G��""=9-�ho�+Gy(�٘�������ݟÙY���	��gЮ�U����>�ӂ"�:N]��J.�=�{����_� Ν���UD�iD�*6�y �T~$��k���m��jn��������Js����H��#zĦ��W��V,��&C�	��j��YM�ZP�A��yU*SP��4#+1G#9|+U�aˈ(��_,8��m�������On¸�{_8����B�Tٞ9q�Sgpt�!�y�\:ys�- �5L�ZY5%�F���VW�,Fh�� *ν�>��=�8|O~�d����͛b�V[��Ņe�]��W�C���Wĳp��o q���l�C�E���(W�E��\�������\���_�.V�^��&l<oU�+h|ĉ#Ө���h�P�FS	[���F��
�9:)7ͯ��y0��C�@�1e��k�g:2��6�-ѿ�>�2Qè��u3xP�_�0u^еL����ȝ��`�T�u_˃�,#x�,׮/�.V�π�t��X@�F(	 ����t���.ؾ΃0�;��l
�Ԥy��LT�Y���TW$�\���h��)3��䵚��Lp�?5��;���A ��W�Y�o�뾄��z	YF)D������@�=�?A������h�R�D�Q�=��t����dU�fM�}�՛2 O)fg��a$�1mט"������~!@�S۽�,�k_w?�u��]<���8�j�OӰ7|�������\�1�ť=s"����T�2�Y�G[S!lq^�3��2,\��Ǐ����a��O�|���~�v��ˎ�c4T�xue	ͫ.�v�AYn��w8w��؃��`hd��ՁAs�ٴ�r}��|�"�}�5����Ȉ�s`�UV��׃,y�(s˸Z���hcQ�ڱ�~�O?��C|�ʏРd�H���\CS��8��T̓�6{J�i�O[�:za�5�a��Li�U�w[3��y��\����]܆s�1���
�4ԍ���(`j�j4#��	�K�MOT�TS�a{�iJ��~sj��DkO��V�&-"a(ţ����,f�!-�+x��/��;��ᇱ��\�q
��m���C�PB��Q��hT �YA�w�&�p}�.��Ǹ�Λ�΅�G$GU<eV�䕖��p�w �T�f�5��]�n+���k��	�,n�؂��葅�?�#\>���"������ez���H˽���
�)z��FU&��<��,�9��w(�|�8]?���8X�d���:����f����,�!PA��N4�^W��=~��^Wփ�&^�sw��{�Z�4�e�(��������-���}�׃��
:�7�\��r�7�����'�u���6��A�t��չ*-������Ef��W�����Yw�]q�8+���y��=�5S��� t�(��CN�#݌n����'$(P�cD��o4�z���N�T��L�$�3��d���Ǩ�3m�w�A�PD(��C/�4���-?��r�G�	T[�3tZ4�\�?��[i䠋����l�`>�5`cF�Cktu�>������ϣ�&�� �{�MC�t�z:��Ͽk��Y~�&��Ů��Ͼ#����0nY���>� Jl
���}sd�� �m�Ҭ�q5�ςNKU:�Zt�$O��AvƠT�|�j��%�����!?��|�7��Gp��`yV@[?�����ә8ʲ��~�!&w�����'�����O�{`pd�hL;KX,�\��ۯ�'?� �f{�Y�NMgn��y���X�l/*�e�3	,Vqn�:��������K����Q�z��"I�eu��j)ƠN�U���j¦X�%��N$�\�ƋcU�#��B���+H=��`��s�g9jr��}6G��p�6��-=���{�j5��{�A���O����S�4-4�'ѓ�NM���D����-�MC�&v��X,UP���%�^����{r�Q<���(Ξ��?�j�E$�q�j~�BSW!4K5�0K�8u9��X6-�Ak���+�Q�ᓇOR�Ho?zR)^&�ڕK&�:�5nl0-F�����z}�`��;��Ķm��o���K8}�b��p�I��U�S�O1�5�VU���gc�M
�U�nt��91�/Ȼ�a��7���pY�O�/���ֶw�+�ǿ�M�u�W��0ZOu��yFnWz���� nx/��_�������V�����B՞������)�m��Y�N�v���A�����˞ѼZw���(5�����T�Ү�y�����~���)N���5�$���X��>!�ho�/�B�-��?���E�>mCS�~{@F��ij�qS|�j����3����؎��v��s／�+?���NL:�����Q	sK˰d}S�a�9�J�m�*Um�0w���/�B���>����TЮ� ��dec�2z�p�5VgL�%�/l��aqE�!��qD�T�I� @u���k���F�g��}���k�+H�c�墂%ꘛ_D2+8@ދ\<���8o���Nct��3�lM6�P��r� ֮kcb�[f�ݢ6
	ZG�M�l���N�,�w�y	�Y�qB&�Ϫ1���5z�D���&hτ��Y2gEb�pR&b\&�P2�%�$賅��y��G?@�?��|�+x��/�u<��[&}��SܑDθ͊�8��m,n �v�H�U�.)��c����e�Ļ�e��YpHO��K#MΥ<��MoB.��Y�1:�g�+x�cX|�\��о~K�#��5X�6:�}�F���EyXe���2�r��0y]߷���Sc$��v�2�Y3��Y����FR����������� ����U+^����$n7pD��6�-��lqt��n5 �t������^�tmx���V��C����wjA::8;ų�D�����е�&����6��A�ў�䓲*۩
p`�+!�/�������`糏�/	��{��w�5�7��F�X�� �Jˋ7p�ݦJ&�� aG�D��*�q\�H]pL]ef(���B��]�x�ZBX�1噖d'.�Cdr}�3�֝��~��O�A��Uv_��W툑�഍�$^!<�XBD�7%8��V̷�B�ɞOe�i8T#�W(������ʽv���Si�0�jX/h��G��j�4Fˌ&�ZDO	�.����$�è�`�=�Jz���.���U Сid���WCb�CQ����b;�g."��[ػuƞ~(�����TUy�ZQ�L(�XKI���9��摨&�3�H�2h��J~ ۦ���V��N���Z]�\*˵7�[ �_KWvb��K���~叏�o�������u�ˏ�-F8K��m;�SA��w�ʢ�͜Y~���2��G	���Xg�����,�rS�/�?����Z���ݺَ����~�[;�(��j��u���* I���0��m6�K�U�U����x_�5�M# h��/6: }��N�����g����/ǧ��o#7�����C���� D�<��ɺ��|�"��g�n"�CGAB^�P��?��l��`�b��g�ɸ~n��,8���Ҳ�M��fA�/�����tok�E�*sV����~�LK8Ţ؏ضQ����_���	������o�^^E"�jt�!X��{y�'f�6���R/v,b��9Q�i�VZ��s�]����uW52۪4������V#�
-M�i�I�R��ٸS^>��>���&��Ǔ)Ԝ�����X�z2y�:|Gn0�*�M�{p2- k���,Aj�0��7B�u�8~Z� �>���1|y\�茖EO���?�ĕ�`U<L�����TFe5���K�g�X�ޤ&ZJ����4+Q�m[S�;�H�)����>����x�W��һ�������{x�4�h*��\�,��[v�`� �S�|cI��R�k�=��kڰp������i���iǚ��yV@^7|&���MhC��/����GGr�������*Z�����q�ة|��'���(Z��Nن|����7s�֏V��4_��֭�%�1$�\����:ybO��l<�IDo��M�u7��u>W~�����O ��4o� �#Xe���i�9�����~$�i��t
�X��BLF��.O�.�֜�O<f���Ŋ'�d��D(�so�������������K��lc��y��w��$B���T!y����a�J(U˨7(,.�[�aW��V���Jx��E���b�am!�`O]�1'._Fbz�������� �n���x�g?���ED�
,������U4*u�a��n������>��:��9��f;+��`[������W��4XeZ��mĐ�I;S�1&�#v?H�Y���+��]���(���#�?ȝ��b��=��Br���������$�#V{���Ʊ�I`Nn�Z����n�^E�QF�V�O�~Snz_���;��K�w�Ͻ��}�q�];��.�A(���'�C&ugN\����J�p�2�sQ~L�P�-��}[�r��B�M�gω����/�
�>���?y��ɟb������uA�=p{{�y�6Ћ��JǏúz	)>��
�k�a! �\��g�41.òZ�H�"�<�'])Z��$���TU�Ӝ���� ��~dA��ݾ��8�����㝶+��1R���F]9��/��aRJV��k�;?�)��6�����>���f��/Li×�	�d�H���l��O�.��q�������Q@�=^�ѿX~Ϭ%��*^�!Yc�ju4��v��|�G�����;<������~��Kx�՟�Z)#i�g���<w��mz�<��V�R|�`J%��3"aKۿi�gu�K��<�-ƶ�������/~XX����Oq�?�����웤���E�V� U��R��7��h�_�NA�=���1`z:"��Y-����m:�x!�[ӹ
y>���nfG�}��6B���O�б�OKQ�2�"�u�	^dF�D�,	4N%���"@j!�l.��l3�a/�d��!�Պ(-TQ�@ly�2�۬�A�j�(ʵ(��K�vY �;�L�V�n`��	��*ڑR}��l�v����
����il�Gq��˘9}�f��.Vo\AX>�n�Q�UU!Yyjv}�|񋿊�Z���x���K̜=�S��Ԉr�H�}��?�u=+Kh\� �Y՜:W�c��� �p���9� '���� ���A�z���ٳ�i����_��l�w��Ѳ�\?3�u)�_LMཏ �JpBp�(^��6��tf���@
@֝�2��^Pmz���gǡ�:o��42W��N�{�#�?��#���K�1�U���~�w}�V�/ǧi0���J�eTO���ռ���L�����hA���d5��R�  ��l:����,���_�KL?��H���~��yD�ލ�f�"u�RO+�C�����^_� O^f�A����H&Rb3�X*�P�����C����[y�y��".������}��.�Ix'#h�*��
aAI����B�b]�RU���ث7T�%�m�XMUPת�M�j��WZU��YU.�R;S~��ζ� T%!na:���Tb��NaR��"��������ϲ�¢7Z�\v������,01�r� ��C�$h�r��G����-�Q�V�9W����T&��9�F�M�s�1\�|�bO>5����W/���+HEx��_C<3�H"+�q��C���T��^`x�a�^jayE�u���#]΢2� ����ޅ�]{q����6��ro�ݷ��������{Yv�gb�9�ܜo���<����	��"M-Wiͪ��^��r�����.��/{]����*K�[I��H� �` &��n�����y�9�=�$R$��OΠ����ϛ�w�yT�As��1l��kup�TB�\Fd��� SW6sm��MkF,uA{�x�s�|��I��g�׷��A��S�a`u�o��y���/� <[!���ړ%��~���>�O+�z����ô!�"�	�$�i�Gª�;���}�7/��9��V�w�v)[�p�����8���xw�G1�뉨ϻ�E����D<�o	�-�K�_]v� ��ǜ~K�:�.^{���������S����1��g�-F��{�Ut7VP]^�AZ4+���������-	�y(@�+�\k��E��؃9�/O~�y��ߧ�������7X�=��o`��D�����K&7��fL;Q2=��.��������Qʩ��k2�~�v�Ʈ���T4)�!'�������1�W��ܹ�S����- ��X�����SO�@&�ި��@ZP�g�a� �]�ɐ��@>��Cݲx�4��4*�c�<�Ǖ|�e�#��&*+]A��wgN��SY@�:�PAAc�H����g�����>��o)�/��G��������G���M01c����R����޽�T��$�W��t��P�I��ۏ��^�=��>�����+��x�埡֨�,
�q%D^^k�މY<�g/���8w�^QnH��-������p�crJ�0�8sC��q�"��E�����ճ���%��?�ز���_��U��e����O�,T�j�c���[���2�������s;9�8��p����A`HaB�H�_���a��E�;�/�4�gn�o�<>�R*0Y�6�0����7��������_�q)�Ǹ��>p���ޏyp�x�TZ�-)��\T6 �0�э����!������O��"%n�y\��.^��jX}�m<��_�����p������w�t�
n���V��F��U�i�������OK��$�n��
��x	�b	�z�}�i잞CvVp��,�����o����3�S�h�Exf	�ڮ�������W�g!^(����������
VkM8�
�"ٸ�3�f��Ѷ�+f�����0�R����*���F���Y~f��U�t�;�i��&��&��_Ykh^]��k8V�� ��d��wF2�n\�ё4��(��"���~o�`:���18��D�l$
�I����$��O�hkN���ݨ��L��)�/���w��3'4{�U��g���
6>g�c��#����/��SO>�7\���2N����&d1�(�Lf�(%Ҙ)aY���v��?A��a��)4ЁM�-��#��'��3�{1Z� ~�"̕5Ds�B(Aձ������ǐ�ZY1#�6���K$��Y
��?�|5�&�/�'���rȷ���z���X�)"; ݧUŇyd!(��!�_�G���x;�S�� `�-ʶr�B0~>,Z�����DR���n��>�<9*�0�z'㣎��_l3�;���]�L����04���ʍ�j�>�?���A�O/��d�/��œ�Vvy�^|o���>�G�O=��S���pz6�k�XY����:*ˋh�/�{r��5���3E���5���)�Ӎ�U����,�y��~�Z%��pX���7:K�Qk�@ɘ���;��ԫVQk۸���<��_C��n�,3{��hH��.�Y�0�2�;8��G�woW���q��=(�:�̻��`j�%�ЧW�D�-xgO�� ˴L8�_�lGY��3`O�L�P�	��)��\	�y��7p~}M/���C�IFȎ�3��Š�vd�����}A�L���0�4e��q,�DʝE�s/���={�x��q<|<�K��~�ō�ʂ�ӱ8>����b�2����x鴋H��B)�N�&:��;�(�.��S�,���XW΢߸*�$��KhK�ސ�0i���{�	L˻��|���H�"��h����ꀰ��%;�<�.�z�E�����lJ<��mܪd�"|Z����I�1��;$��:V��Y
�,�
��y�ۍE��XvV��n��nЋv'���vfa��Gyy�z���M�`X�z8�=�M/�]�ww|�5 #B�8e{J���a�H���#�Z���r���4��w�������,���{F�Q�c��,�_ǥW�½�����kn#�a�������,@�- �O�Ad�B��%���	>���]\q	�x+W��].+1qq$�T"�z��ҘE�n�E��TF2��v�ic#�@A���_�'�%����ߡ����~��Е���}��6VX�����uL:9 �Í�O�<��c�H��a��BV@�X��P��ǝ���[�� 9�n5�*��&D��2F���8x+�����p���J��|w���Ȳ /[&��d\y�o�*��IgD����xzr�2��)��)�$I'�(��n�c��+��7����Gv��C���	ʗ�����j�x��Ͽ�~r&��;��b�vQ3��k�.V�,� q{�i�Ne!�[���Ѐշ����OL�xa��'qy�:�7��:Z�8����)���blkd
�I��1|D���2��w��1v:�ސ۟�.���2v�����E�7����4@Cړ�<������[��kӋz����0,��*�޾�Z���A��h^�^+�S��H���;�� w���'p��~l���ڙS�b6�J~�R[��%�3V�9z^ad�F��#=	����������Μ����!=:��]Ә��Bq|c{w#;9��<�۬������aխ
X[� ��1?���F}��؆�������y1z�;xĢ�����<��՞�<�c�=���.��_�����0*���b^)����C���x��GQ������7���9hcﱣ0�f�j[ �LR<*�A�3P�]��i���
/nI<���;�u�P��,8#�;t-$�e�fÑ�NZh�w?� ���&Bv��T��1�o�Vb@Ү��� ��bm��L#��2q�E�N�M#��;�IY�t�DR6B>-��av�,���0���������n�כ���(��

�)d_Y��7.ʟN�;�ڐ$�}x�U��;Hgw!���w2j�fG�J���z�l�ْV��F8������y��{Õ2d��	����.�R��-d�����pW�xh�F�QD~�-[|��I���n+�f�=K�x[t:T.jq�>����9<��N�\�OUS��0(A=[aq�N~<���U�p�Rwl�Q�j��"�����>����A��t.�F����C�X�6F�wH�BO��qw����?����>� ��;w�Vo_;���ef�t�j}�B��*rbPu�02&��Hg�6��_:�[DKۚeSt��՞���J�����4V�kx�l�=A�]b��7���ְ߅������=���Rν� �A��,KG�5�U��!�-�4���A�g�K#�M�0]<1�p��H�q na��;h�f��O >"�6�G�i"^_ǍSW���a$'0mcY�%�h*�D.�H����"YǗ_'\��X�Ma)�2-�tbd�F`:��X��6.�S�O�ΠI����Y%�w{q����&�oؓG�ɌGc���wj=��#�Uk͕d3��(
Z��# /��]bu����'@3�܃�G�Eym��Z�5��p�va��u�\�����>~?z�+"p�j&,�ڸ��bPk"�UL����ܖ�R���Z�(N��IcO�y0\��a��i�]���l��Tk�6�򞞡�=�����تN&�#��G*�����|ϖ5$S��㳇�"������������y�����H{!�0̀?:���;~�ǝ�s>�>����ZJ����@-�s)H����>x�<~��8�s�ҩ4�Aŭ���G��ٙOxw����IGQ_�I��U\_~�$c.^;�\e$C�S��7ɱ�An���79���?�1+�ٰ��X�ю[St�V�Z�SƐ��D,_�I�6�h����.n����hF�S��2�!d��hD�J�6�;}Y+#�/�� -S�]ܞDV@g��[o	�k�n�c���$�g�F�ƍ��1"���1\z�-��(c��^�f�����x��F�o�����3_�,��p��y���I���M�����Ȅ�r�1����ώYw���<�M���r���-?��ԧ3hå\ ����;g��D���K��^@�%�����������Epc�̌���b�Xk�oh���@��굆 ¡X���\ũq�n��6c��Z]F����4�9��M����zJД�fpϮQ�����}�E̯�ci���Ү������5:��6p�r
'����z+u��D�
�PY��,���uY̶�W\�(��l^7f*02��)��z�C���A_K��r�EL�`�� ���W��Cu<2>���%ߞ��w�x��@�Ҳ��k(�%ݿ�w�/rl�K�}ʰ=yW�dmxw*Z�QH����
��F7|o�'k�v�A���r�n��=]�׏�;���#n�1�����sR;X�<V�]��;���=��=�,��|���P���]���
'��S/�����dq�(�6=ml��T9��|GriĦ&a	VH���P�ç'ڭ>`�)x�'���=_􄳈A^&&p�r��WK��S�����O0M��Fʌ*��Z>�ۜ�Ai*��E$��._B܅{�����Ckx�����ko�'sp����.��L�������s�����`���W���ד0�#�����[�r|�o zw�;<y��!&���E2�dA>���}޿�����E�zek՞X�	�)}X����^W ��^��1dcI<����G<���g�'K$dR��W4'/�ɠ�\RȃЍj��ml��ĭ�BqR��@IA�׮^���ࡇs�;k!)�d�`2=��Sg�Y}�U9��u�ΧO��ڇlD����8ۛ�Qۈᥓk���|�.-c��� ���G!�B��X:��� ��l,���;�{y��b=�d��y��UF�l���޾��e��o�g���LCL�����N:ZPZ'|�Ⱦ{~��_��c�i_ʰ��v/���z��!#�*�fQ>ȣ�
�Շ�z����Ϟ(�����\�YaGz&w��;<�����gW�%��:!�l������vk�Q@.H��@Yy����3{��n���Eџ�:d�+���7L�p��%��,W0�-�Î��������E|l��qQ�y,�\XkwP-W�uF�u�91����Yd����Fن�a�
&�~�8�;Q�;r������.z84f���9ܻ��k�t��f+7<����Ǟ��?��2���-t��"J�q�J�\���k��]:�L�����?�U�.^Fka}9�n�rBp������~�퇼��b�y�v#�$��W�I|��e����� ��dn���nKA�y�����Dn3��x��#��u��;]�T;�=*�UTj�9����QY����������g2�$��p����L��`}a��,RC&�+/����Qį��P]��ŕ��(�(�f�aq�:&��(e;x��>���7��i�v���bc�6��_�w_��"��V�L��=i$0Zo`��$�����&�ʝ��@@�J���Ou��n]�y=�z#	�\��-(v��hn�&�s���y�y�Xb3�N�� �|�����`zR��v���D�S��Ɛ��pvZ�;)Ovl��)^���J͐���e�):ݎZ�4�aC�?)1 ���z�=��(���������3� N=�߫��s�C�h����F,������s�Ƹ"�Y���~���wO�?�ӓ��j��D����Gu�=���5lmw04"H�����#� �B&�h��d,�{��	8w��ܷA�]�n�j�m`��n|q��g�P6��"���Ɂ{~(_�o��u�m�lVq-�'�fArT�o�6�Q]dJ� ��3�dhԃ����!Đ�3�����ꌀϨ��l1���R��}5e`;���Ct���h
�H�,��8��F�*�3.�z��*��O�J���N�{��p���7���ð���һh�z8���H�i�ڭսg��?��ocfj�<�A�2z�%�jUԵ�nyy�uFlhk��'�V�.��+&��M-1�����}8-��g��+H�)$�	A�2q	ٸ���7G&vj����ų�=�k�
9��6��折 �TL �aaqq�� ��zs���8:�n��� �$�g\lɵ�����h�f�^Y�� ӕ>rY���^����D�A�/	��afrV�����Q����ɸl�aK�6�%������056�b�
�����6	'��˭&�FDi�,5������%�6o=n��z�R���
�=1����p�Je�L���g!����e;8�E��i�Ϸ���U����3��4v��_}� ��i���FHnLϖ�g�B'�n���T�(>,0=� /�E0����w�XԦ���Y
+�������ND�w��q����g$�r��Q��6�{����f�<��ÿ��E�;8C�\����f��a�q� ��a�Q�X&�f�wf���F�0Ew���h�CGP�X��5����<��4�p��Ԟ�l<�gK�b
d�tb�0jU/d0�Kbu}Q�sJc�	T�ťtcc�In�Sv1���"�Mc�0�Z�'����M��װ!�{h	8�&���L$f�پp-y�Υ�-U�q�� �>�	�W<�lY���\ĕ���C!!��g�z�!=$M�R�L;�[�2�o[x��j�8��8:2�Ξ8�����.�/	x��M��5г��Z�.��رc�J�3]�މ)�%�E���	�5,��Z��7��L����R(כXZY���l��qs�f���*]�G���2���HX��È��=�Mڞ���8�u�ڊkii��.�z�0�|�
�v� ��X}��t�NK��+wQi98�'������=����8�X�ۋZ��{��Q��~هY/��D���?ږ��L`D@��
��k58>��u(|;ȹ��}�!������r��q���-�|=�ޯ��7v���N����`����aaI�8��#�c~���J��s�����0m8�s�d��$b����Jm�A���U��y�����=��K����+,��D�i�Xض�#}�#Bu�F{�9����6V�B�~��<��!#�-��\٣Q��V�}s�O�pP��0�v�)��}<��G;[P�����z='go��a�3@��b"��"���[ �#a2�Zu/�xГ��qp�8�K)�;]����7אJ�`��~$�iX7p��!�sp7.]���뻈�rH��
:�����Y[ H�J]_�di/FG��R"��`�7��\���k8"��}%L�͢�λ���э*]c��F��K�-���ne-b��V$* 8���:S�^D�=e��������Յڔ����$P�1/B�W�qv���Ŭ������ �� ��%�h��~���xh�W��ɷ)���c8/�O�2��r��Q��e�o./���2�x^~W��L�+�Y/˭|�ᐡ�LpF��;�>.��K@c\@�ܨ�N+��0�m!�w��y�zsIg7jw�Z�u4���Z�M�Pr�B~
�����:n,�U�qxo	'�/���'����,Εg��6�N�%+�}�9mr]� Z#��@"�,�vLuk+����9��M��PP�`�EW��*0:�_vH�;!)l8\�����¸x�}��_W|N8z��6eڹ�0)���[�N����>.Uʇ���O�oX4�!��-V*e�.���B�tHcD�F������;>x��U����I��]��Ή-��p�^I�^��y7}W������O��ȑlԛH�iс}tW���e�w���3e���F����R��J�],.��7�O�/����IEi3
S�FeCS��[�$�|�{zJ0���yO>� N��*�+K�Dٲԉ�g�#n$1�,�ч���D�t�T�xR���I�j7q��5\�z#��6?���C��w`F�oK��������%S�_��-�3���C0:[�}�2�K�x[��=�8�!. ;*S��)�9�w��Y��!?� ]o��� �/C�6�2�i�f���]���.]���E8l�+@�V]Ø������9dR),�׵�"2���
�^Z���
�]Ʀ\qme=�ƒ��e�k8��`�ک��J
�K�8���d3�^E����xq\z�ln�� �.��(VWb�?sX^�+B8)�1�J��\��;�VOcV��T�h󂆳^�cs�V�Ɇ�'�^�	X���	XK���s(������ܽ���r:�����b��A��X%�u�&�ee8k��"l�fƷ��Pt4��f:x����~�ñ�N&�
�6s|B�?�T=d�	(�Q0Q�W�'���s��_��N���ø��r}W��v�ɀ��
l�X����=��p��h�ֿ?�=x�9��p�#��3�݁�o� |' 8幌'c������h�xD@*��p�9����ʩ�#�|]���ym۴��n�Mѻe��SN>�κ]G�����?��}/�!�ʖ�Ѥ�y�u��,Hp��S"3b��ۈ%�S��c[��)ƅKn׾͑˩6���Eꭃ_�@=/;ô�!�+��z=��Z������I*Go���AN�buv�}Sx���i����b��V�2z�-S�E][ �`�+׷웚���&��0R�b����|7�4��MXY���!6��H�X+W�!����Z����}��n��2o����@pI�c���?�k7���Wq�w�|2��c[�-�4���RCe����8����{�Q~���{�?��js�1�����*ݾ ?�a#�2oϺ��DN�-��w�ü#�᪻߂�])Vj�~�^�wa~�,�%�KQ���?����Ɋ�vm^�V�f��e��^�޵c�%�F�pu]��,��ª,�O�ܒ��M�<xB�=*�136�b6�9wS��(�"��e����*�dBss�q~�ദ���kb1ˌA�����[C>G�����ă��OO��vp��j��x�A�3QLM&�D8�3�Y�T�����c1���єMT��a�I��X������0^�~�:V�W�ęE"mA��|�?�,dP �;��0�u��˕����k��S�%8�;~}�G����s��4W����g�m#��
X&����OBُ[^ؗ6��� @�z?j'
���<'H~���W�>=v�\MF�~W����Cav_�Ie��.�݊����q'����&���3�����4g���P�M�O
�5��o�����gf׋iq#�]y:S�w0���t\����,���bt���Q���NWtsK7�Y��\��4 *�nQ;&x"��&&ħ��r%D&'1��崋K�����%�U����Ы뇒٠A����512�}���3�y�Bu9'ˋ����:��w�zW����4zC8������O��0VLj��^~C#��\
ϟU
4�k�V@�BNt:��N�����g�gz/��9�+Z�j8)�kk�5��2�����7y��z�5pbf�=�v}�<�n�l��dd�b�w;Hpb��
��R?������Ti����:��ʫx�䛸$�%?��U�`=�k�����G�G�����˸|��g�d�c*|;%�y
�f���q��5,����l���t�	r��2��31|8�g7��كt&�b./�,��}M�K^@v*;��9��\���6Co��-Z�6bb!�[]�����T�~���5������fJ��s��ge�<]A49����8�/�Y�ʂ�,;��$�Û��De�D.&�!�b[����^YCk� �=q/r��c�'/�����xɼ<����q3dkX�V��P&���bax;<�������5��0�v��]/ާxa��>V1�W�(�%zۻ=�.T"�3�NL6��n?�|���{�c�?��>�mW����Aa��<��_��<�N�AN���pn<j��/rՉ���Z!8t��X���{������/$Hb���sx���V]�5�V\�<taq�ܐz߰�Vs4�ee��QD,CS�\7�x�:?��Jo��H Z�\ F�ю����Î�H��i�s]Q�}f�
C@R�U� �[���6�c#.:� )��ݱ��E#�&��/�Z,a1f��*N�WQaJ���@�g�ȉNm˔0e*�`��8�And����v7ke�;{W���C�2/t@�����u]&ҹ�Z�O�jXE����)�-7q���O?�a%��'�%׏�7�Ƥ�h��J�+��'��7ɨ�8�9ڛ�z�����j��U����T4������J�*'���݋�S��k_i�hw��u�~	��oD�ȓ��<㚓�s~����"��Ly�K7��{�����v��W��o�{������'O���w���&@j
�~��(�dI�m��ś�x�wqqI����$�l��\l4�W7��~'�-S(�g��Ǒ�����\����4Кp��L+���X�$�$-t����q���I�=�6f��8vo)��\<���-�\�169�+���T��{P,d��M3�f'�S�6�g�F~c�8wiYs���qy��N5}���PL�{<��b'��u,mT0�L�*A9��A5��#3�Њ���������a��c�X�NO]@���<�
ֶ:]�J������{���3�[�p[��'�@��7~����9�=�C�_߽��;<��v�v. }w⵺���~U��m�H1B�o�5�'FDV��A�B<��4j>.�����tE�A	�qg�`<��^���F>�>�"2f����t�,:C�M&a,�Y�'���4����#� �U�4�-�K�ʧ7gȻ�'<��G�o?���O����7��FI��ý���w��}�g�~����fm}x��w�����Y������Q�[��I���]g+�ҧ2a~մ�7/�vհ0�U���,(����������h4�[A�ۄ#��r���T�1�������x/��Kxgj?fG$�I����5��ʶѭ�#����.�1	kc��G�%����l�����\������Ԯ9X3�hdSx����r����V]��OËi��l 8#/�p��]�W��H��=y�"^z�M,,-���� �Ρ��s([J�s��$�MYD)�zZ,���V�,ൢ�K�=�;�J��m�,s�bq��d�P����<8�,�<Д5���gǑ'�1�:�o}�����&G@Y�N�:XH��?���݃��Q��g��W���Lzl�C�a����2&� �a����Kdk�
%��u3\[+�7N��.
�H��3���:|�x�!,\_�O^���N�JyX	mU�f�LUm_���z��˨�MԺt}$�ڜ����?�#���OA�Q
��wU�o�}�]����!�6��˵U>g!��b"�CQ���/>���g��zN��v/��x女x�7�೟�T.�3o_«/y���c����/^�w��������o���/�9����_pyi^ɛM95�0��^{�dW���Ø��o��?���Eܟ/aX��A�"��+�������;���؇����j��2�D���Q�F��&�~��f��GM_�{��^�w�<�,4��yu>����Bw����S���h$�A�����l�y��$n�ʥ�,��#V�~\;j,O��F÷ ݰy;��#�м ~H�*:zN�pW4rkB�VKA�" �Մas�A8Gz=��,�5Ke�pt�|I��P~n�.���"����3�^B}�=�������x��s�*���"�,^;���iQ�6�rk�;�n�M�6��h��ȜFi�qh����[1�P��`���!E�j�F��Y��9:��.���FҾGJ���ј1Yc������.X/�9�~�57[���fP�w��=����1���/�/���\M ښ9t�_#V\��z�{���_*�ζy�3�>k>uԃz���vu?���t=QDT���c��/�X�A�w��Q��ޢ���9���3��'q���-���\����\$ʢ�$�F�Z�[�v%������H˿��DAX^�W����e�[u���`.Z�1R*Se�r�O�į�kE�-ڏ�s�s{�-!*a􅠄G�<��0\	�ZQl�env\эZ�I����v=/ʣ�ߛqF���|��Mά���*�v&�{4ʲmDe���![�e"�S�[�5o��jLXrC�9zX�k�[�H��&�)\�1/�6�T2���QI�C����V��V׮]E_��I.Gy�F�!�+��aT��w�>�FFp��UܼyS�n����K_6FG��\�o�O>A����,
�`� Vd�DSId�%$o��(_���|��~���7	f�N�&���������2]	y�������

m[�u%aə�a��cWl����h2��{a�4��'����$�a����]�v"�K��\Q��6��x���^o���;��4]�y-� #�`�S�'8�/���ۍL~���O���&����Q͖d{�a����h��e�-�����6���d�����@)�b2ް�.Ë��E����n��.�X_�[�Ċ�>�v������� ��d�����E�r��e>�ŬңT66���WN]D��O��&�8�f�:V�jaز4�͓����"�H��Jc=x� ��c�'��	d���W����/b�ހ�Jk��^��G�|��� 7�����Z�{6�5e�SQ�$�>wS��wm�L\��F	ـ��D �8����x�#I3����*X��6���B�Cp�;ۈx�LQ�	\=43��<C]ԛCy�{p���#�r�5���{��Tl��c�o�xiT���x�5�������I����k��^�7���F�)`~�*�cS�O��Vy/������/�6μ�ܼ����2�m�f�B�kk����ށud3Sc�d1c���h�����SbmN��`���G�����_ޛ%�4���(�m�ƒ�T<�;F)��$iChO�����<�-�x��܆g"��eG�[[��AM�-/@�`m��]��7#��y]�Qw*��������ix�Bu�}"t��ψ��@��N�6���1�^p��}ٛ��2W��N	��'�;
xv��l߱�\��>�Ö+$h.rKǉ�\��_$��n~��Ф��jvfP$*K:�8h�+�;����]`H�����Cezbb���������Lu�t/:
����P�x0M�(��R9$�~�\`$����j�d$�Q���*+�}"-T�Q��w�(J�D�&�S��>3=��c���E� ��q�aU�׷ڧ�~�
� Rs��o47Eq݈�{e��P�G(Lvow�z��3�|<Ҡ�p�����9r�r�!� i��6����Y�:�oT�x�)@���`056�h]�mk�l��О B�s�E����!
d ��EmUh)νܣ+`���F����r��te#ّ�$!c���xD=��tm͓6��6���kGL<�B�� =�]L&�Րڳ~��	��!�kr	�P⩘��1�v����R�X�t]�Ϯ�U��!k�vju��0wj�6�P=6;9��W�by�*@��ѳ�o]���{��a�M��~?�2���f�KgDo&R�ʞ�����ML�
��kh��dH�-��9a�9�|m�>��5L簾�������� ���/�\�5��<gl>��;(��8z�2��W���s�s�\j�CRt�%F��2\V��u�^�����̷���\uyƞ��0��g�]��A")�a��栋԰�]i`� �1py����~W������Z��:��y� a��݁`�4�����Ve�eϱ�<�5X��Ֆ<K�Ւ�_t4�{���_cb4���<Ν��7N'�]�J�����t��s_֫/`��^۠ɾ���	���1S�S�)�9�u��L�����I%��9�>�B�亪����ݓ�����O�.N�uq���������x�^{�-̯�`�\G6U������\��������&�ޅJL���6�M1�{�u�2w�����V/���䩖����+�������%yX[�ɦ��3'QE��{�����֌YrpA��0W*e����Zh�K�@E����Y<~�	<��C��}��r���5o4���>�����	�(�|0g!T"�(oz�r�q��s�3O���$h�}���7p�������~��kx��,�nS�ҹ8��pn�.�'���³ϣ_���3gБ�<U��j��o$�x �đn믜��=#����p�{����cn�GQ�x�U���U�3�����@[,���X5b���H��8���`�I	s�� ����Լ*]t<(�!��B@�� �]c��4cz/~��W6+�N�KVC=��'�c��J�(�p��,t�1b]�����Lr�1�C�]Z��7il��1���5UQb��uD�-oW*�F\�b*��œ���%��̇\�)XĒ�F�u^^��xtU�r�zcy<AC)1n�ē�y9�P��>�>ޯ-��14��"����}C���h�C�{��wB��)	��^�+g�T��8������xӛ�ꉥ �i3"*���q�{����)'h)���ƕ�P�u�p��= E_��Rku�ۙΈ��)�\	�O�s�	�w�}��� �'��A�f���`�B�y9�{� i��^=*ϐh8�T�yvr-�a4��-rjuuYޱ,6�����N^�u	IQ����po5}o������#YrxM��3��m`��k�4ۛ�a?���������j͆��4e���� P���]�0\0�4)��<h������n���q��w��3��y�_Y���ޅQ�'��\S�|�( ��z~D�:C<�,�S���}O'�ϕ{ud�Z[By�Wj��,�1�#cb��
&Z�/���'ήV�7>0���K��#Jt��Q^}�;v�R���E�� L����~�Wm,�����.FBTvp0,eX�4Z����3����x��{�����=��&@p�*���*����sCK��U:%@Z BW���C�=,�^���/#"ù6C�F��9-MZ�4�z��VQ`!o!�]�Q�]hp�DL�F/���1B/��
Y����$��~h�>ݯ8���.ä7^ g?%{-�������""9��q��y,-w�ϒ�G�5���N#�F*C���%`ݒ?F\�k̏�����c�k�n\ٰ�m ��W_]�Ь�="<v�3|����e�ʼ����I7'�dph5���Ja�5mr=�YD�����_��o�]�����2nT�M,��MYcG��=��ǟ@it�\÷E�.	�7r �Je�b@��&������3�r�u��4e�ڮ��y�v�`.*s-sKÅƏ7J@�a� ⟣�����;�LC���S�+�`�X�?��|����tqN�����{���=>��._��_>�+7˺'��vO��k<'�T�1.��##h� �+�!Ƈȩ��_O��<�� ��66Q�b���~
���1�g��#�+'7~�ч�g���?�G,\�)�(��,ڠ�GK����
��h�HN��X��<�b&����
�=��,N���E6�g�����J�]Н��c>��^#����+�p�X��l��%\�梲r.v���
��hl|\��X�AGމ�ݻo�s������g��o�w�襗1�w7qk�*dsW�,��z�,�2�G��{x��:zW����ò�(����2��<�uQ�L	�s#4���@=YQ�����2�S��D��Ű�S���TJ���W,j�
pB�����1fM����@U�~���N�B������(�x�B>��W�EA(k�vg�<�����4���mԴ�[C,6���ь6�6�~Z�C���U�c(��?G4E��Hs{�O�OlQu��xI��%U�G���a�O_��4��o�E��W������X(��	�s��+W*��W�	*��Q`T2��{��-�jGΩzE��o ���Oy�f.�@�;+)<b]�9;x/4\��r��~义��<����S���u�+���Oi�RD�8l�ù�sW�]
� ��6�����90���~���#���WP+��g�z�x�9�岴�����7���NG��޲�ڹVax��& r�zt�
���{M�ӌ(�VF@F<:x\��2���<������d�gD�0tK��Ķ�<���P�����Uϝ����~خ���)!UC,\G�ng���s۶�7������!9.��e	���sH��&@S�Ȉ/ǽum�μ#�_v��t� A>+���B�ݱ|V����U����Ւr��<��
�T~2��b��8�116=�\K��h�d0��J�#����ً�'�V��˞�(�"�5,�|뉅F���1�)���r��W�w}�ĳ��H/��n3�.	I7���&n�~�0���˗
bP$�"����FH�ņ�M�gӌv���|UV5�*�ڢ�;F:힜Ƙ�>E9P���G����	���u���L#�%��Z���hݺ>����}�^Q��A�v�բ"�(�	��4l�]5R���YlJ/��|o�EZ�$�&������)�\ x���X\\�����7���T����L(w�*s͎�'�����:��:��-j-�_�WC���Y���Lɵ'˫(��D���"�k� �ҨM�Q�!hyV��, ��Ve�iX�#�<��P���ɺ�"����&��4޻�>�w�����#�"����㵓gP�\�y������a��rw+>�igj�*甑{��<:L�A(ޔ{jOX���犀�����S���o�,hQjs��S�W񟿛��h��YB�����IT���pcm�|�E�N������}��E���bp,�ѓ�sO�b�nK��eљ�Ϧ qt��u$�Z2�4?zg0���Y"�f	_8�&��$�[5����-&/x���x`�>\:w^ݢ��#�~��Q�V������#侑Mk�@(�~L �o>�(�?�	�����uM�����Zt3Q\AضVY���CM�go{�$��ť����K.�L�p���?;.��(�y�,^|��͉�"�����bml��QY��^��G?z��/���{��{Po2G�����[�"%�<�X��I8�?�)��W�����}��XB�v[�35QX/��=�6�\��w��փG@B�o*CW�މ���I��2�=zL)��، ��nnz�yr6��hD��<fiY�w�m�7(� �h9������&m�朰y�iiX����Tv�/_S �-���s�"7R�[o�ĵw�ʳx�����:��6��!�6������C=/���<b�������Ϫ N,.[�Ӹ́��BI�=e�[��ʧ�i����%�,sy��/���Eo$=PT0�fE���p�����{�|��wb�0�q������Dض�yo����ˠ;�**%�e&ȶ�}z8�8"I8J I���
b�1q�}�c�6���.�9Ю5�d�y�J��QX`O��A� }Q)�=S�o+W�):+8��1bRV�4I<�Q��yۨ�ueE��5-��i]sm����ẗD`�s� y�������k_ք0ʱ=��W�5U9�t.Sr:���Z��+����b��.	�F2�����O�T�NK��0��C�����'�z�X��x��y�U��ƆHL�f}�eC@7��\�D��䯍F]כm I�A^$=|Q,�ݓ{��`� ��7u3�gC������|�:^ZyC��*��+�[�CAaT���Z���wd��	t��{,�D�uC�2���$�d�Ⱦ�"~0�m(51�e�{Aw��Ѡ�fݖV;�%5Z(W��i1,�����a=���]���-��g�X���5Փ�6�^W��3jD�lx�5�S�(���M�h��sꊔ�r��p˫U�i`�ۨ`3l*�O��πa�3��ܓw���E�'y��Lzs�>s?0�	�yo+r�a¹�t�,�$M�<�iX*K��A��vi��A�����*%�1�3��凵�}��m5����ػT�׆�^����2�/�H�[,�4\��<�k0���Q9�w�u�*t��~�÷���#$�@���9��k������ 9o�B]@��j�+O����������K�3��F�#9�-�NK�#k��˸* �/{;.�'g�gɿe/e��?��܃��,�|�U,\>��\�fh˳xr���,82(�Y�o|,�T0�����P�ard#�4RrXO��F�Ȣq��^����V�2��9-7��(nH\,�M!5��Z����3�V�g�9T�1�+�Z)jTԱ���~�*޺��#�[8�+�?��������Q�\�tA޽-fP�7l\Z��؏���=.
�!F��YmT��#g����yl��_Z��ͳ��$B�^C�NC^�]3x��	�E�����S��l�Փ���=$�5#�Z�0�<������?�<��d�q��i?�F[��~���0�f�ӭ �N�c�XzA�@Pb�M�ˉE)�������Okx�l������=^�^kk�"�F1U�����`rf{�ǈ��Um��@]�7��DQ�'ʨ ���o|O|��0�胸�����%�C�R-r�S��TK�O��5����r��G����"����D`8z��:j�����no���a:+��ۥ ����!��N�^�'Ze��2�B�+��RtD�1�gw���Q	{���{��Bb��=`H!�J��_���b5�*�7Q�?c2ǻF򘘘�/�*J��`�&�u��ɼ�!�����e$�$��5��Ӥᐛ,%Hi�^4TP��M�ɨ/ӯ���w����8��^�;�[2���4t�/t�s��7�����{l�I������J�9�8�FY3Q�}�V�
=C�:��rؐ�k�y�[{���\?1��V���)���ì�tY2VE)�Eη۩�0*��|��~F_�Q������Q��N��Q��Q��ȏ��r'�=s�t����dn�P��P=U~؉ ���Ź�M����AՂ��ZJ L����W�� �O��q��s���H�a�Ϗ���ٮ~88�z=5��e�%Oȳ���h4�z�sb�!��!�z��}KA���q��fK����XI�JF=�i����m��B�jD|/�G�۞���� "?F����Lz�{��,�����ыP���Ы�Y ���4�ވ�ۛ^=ޫg��c#�7΅C9�����ZI��r�D��@%. ��)������6�93��jk��a���z�yY��9��VEyU;G=)� &��HJރ���<?�u�b8R~���!�G�7d-�Jʱj�}]�B��Yr rX��$�o3}����B�X[�H�t�%
�T�!I�	vY��e�F��E���'8��(����e�<��c�?+����uT�mj�%���y�!��Nو0簯������hdT�Z~�O$�B&����:ܷ�r_��S���i5bp��#% Gs?I��9ޜKm	F�nkB�G�<ϏM��Lg�K��M ,��F��lh1Qʍ���#]*��haȢ#����dѓ}ԒW��3%�9խ-Y��Ȩ�Qo\>�^_�~^?�]�9K�J���0;=�}�E:�.��?Tg�@ޅFg��qy�H���%H�"�ܐ�b�&2��[ �H�(:{cz�ލ}ss�g�>�
�cNc:�3LyAӚ�j��r��io��7�������\_X��FM��k���Z�^���u���v�-X#���l�~bר������A���G����HŪ�.�p�<�$�:U�wz7o�x� ?
waI����T�ռ��,�i9y�M\�|��3�֔C]�5lِ�\�p^^lc��*	�X�ns�"�M��g	��:�{���f�0�(����}7�@4%x�Lc��2����\t�ܯ%�Ԧ:�Vf9�i�������Gpj�X���IdCE6��5d�P�V�R������c%�GS�V-4�%��4�w��Q�O���9D�''Q�w7
�<���
*g/`��(�Ȏ�735��(�䡄�)��e��@,�
�Cn|j6Q6h]��,���P��QybQE��O��f�B�,���볝ïH�eM�r`4G$�m��Mc�T�&Ck^�#�$��I���������>�S�����U�	 ꑅG��1�r4��njNJ���ʆ�M{�O�evL��^D���k*�($�]�-��G��F�G�A`�4
r��f�<��	�d�THw����U�3�˜�F
A&k���K�w���
��T�(
����6y�(�U�I����7R��M�K�v4�����8�Q�F�����&$�6�[��v 2��\Y������R�e�z7���+gd���9)�o�j>"������L��,Q��
�������~z8�Y�����g�ů|]R ���W�<t�RrG)� �^L㐽�+��^*+�ԍ�g	���g�,	Om�(��V��E]����r�ԥRL��О�L�;]�~0z^�б凎����H��H�B�)r\A�i&u}
���=Y�@��?�~�
K=�1�� 8Ov�i[E#�xt�3��	zO2O�#��K9�k��_�C�����Y"�W1�*�Q!B�����t��b9Ͼ�U�IB6�,�0㛚sIc;+�5۲�V�Yu����Y�+2���������	X#A�Lbːɋ�����h*�)9e�l
����j���X�u�4h�Dq@ �� ���ϝ�ԋ��fzV=z��W6Q� ע�w�ߕ��%e̮˹����pCCt���h�q^ːs���M�9��e�?uo�d�y]��3�y�9TN5��P(��H� HI���j�%�D)d��V�~��#���v�����[mGtP�m�-���0�y�����3x��}��@��,�"QU�7�=�����k�i\����&ȟZJ2��Q1;~?�ώ��#wc�͔er$����=2L:�F�Vu��z.
�K&��d�� +7cg�r>jw��Y�6����<gZsY ���`-����[`�¤��N����0�.nf�Wg��bA�裆���p���⒀� g%x������im��UY��;Z�/.��݁wg�w�!'6a��M�EkÔ��>?XXЖ��R������?C�� ԘS>���<眃�Q��H-�<XJ��ӎ�do��*�p��<s�<y�r�kK�F`�����Z�TI���fC���������Ao��Ԧ��w����޼z7�d����ݑ�oo�D���$��싍� �ׁ�^��<֗�X�_��I`4ѹ�w	7w���n��ďg7��+�h�XA��*��������-#�-��8n>����!�x�=�]�bY.�Z�+���?����$���+�X��ښv���ezXG��"aW�k��,~�뿆�<�H�A���0�=�H�s�X�,���Kf���yۇ;Qb
O�Ņ����:V�\�����y��<�C�|wq�����W%b_�?����������Տ��T[�i��O�ʹ��l����
�|u���7p�Np�K����+��l`�u���a0ֶl?$�&�z��� �S�PK��u�M �1�d�b����)��[~")����L�<+��)�����&�?�|@�-���8{AtT����GixǁrKX& �l,��)�/��)�4c�(���KKt7j��u���,)=�L'�$0(K�,�ڽ=��qbu�גg��XY���%2ߔ��L�d	���X1\����q`F�^` ^��їHߛ��3�f��̃Y/rOơ�E!p�Ԍg��
�|M4�Ȝ�yn�v�4ND�<]���P�A"b���#����#��( 1�uLe��H��R�2'�@��]n�t��#�l$�0@^���S*��Ñ9l�Oi�Mhg��c��ƈ�l�XAu���|�Y���0;��ˑX��#�Qdl2�NƜw�����I�C�3:��'��'����qH0�(����k�zY�^W�9_鸦$���D�1���Dd=�L�cZ���11�{F�i�K�+�,���5b2美]��kת)�2{I�F�G��;k���{#�L�X:t�c���f��.ʙ"rr�5�޼�g9���~�p��#�Q`�����gI�Ǘv�$�h7oF;���E��)�Y����3^V�M���m��%v����p_���G��9���ۇK9�=�n� o�qr�y�sz�nyR�WC�xXHe��^Dj:����! cC�aSB��,�1��&`������{����j�ha�9�Q� ��;�O��<y��[~��s2��حɄ�r���ihG�=�F�t~'GR5�:5��� ����+�'��L����T�,NI"�5�mt�\j�i�_��a�|�/��NW3y�B^G�u�s٩�lyh3yJ�!�'�{f����?&1:֬���Z��5L�x�#k��we�}i�����P<U���m쇴W�%G�:� �3V��a��F��:n���{���Q��~:�VS��r����jv��92�)��;ɽ���es����6��ČY�S���?�/>�._ǉ�%;�Y>���5�;+�%��>6V0Ӝ2�|�)�/V�LW��+5<V���s�і��܍��������R�<kOU"F�1��S�֗N��_Z���4	 v����4Jb#$8�x{;�?��[�|E�taC����_�;�����K���Gx��0�DE|��+�_��=\�ic��ׅ�B[�����������2B>Mb|A�`���VA�:y �V�O��x����%ʤ#�ׇɡYQccg?�}X��'��k��1��6�3ݎ��]j��F��K/��[�_����;ܼ�]|�k+���_�sO��a������P"����8�4��p���kj�	N|Y�����j�r�O��Ȅb���������+/\��^GA�h�C�� �8�A��5HK��yC�T"�����=ir�$��rfU�Qu��9��Iס����w1>*/:�&m8P��oHcDCg��;tLǘ�Sʑ�qH��:�6��p�H�#��"zC�Wqm�yO�UA �P�����$�a��e��n(��-}O�GJ(�X��� �{���2Ԉ9�R�v�Z�J�$
5GVN��D@;qK��b5��l��tp$;��	�@��7<Z�F��hѹd��O�ϻ�x�
���N��k�aֹ���b�LqE����D�j��y�0x^�H���0�*aK���` $�k���
��fԞ�xH��f� �ˬ�ܬ��r�"�$/�눼nr|�>����(�ɥS
X�X��uU��<�+ܟ�^dY+ir5h���3=�YQ�9s$0Z[ZE���-��qw�T�4?[�0\'y�V�΀J�PDv<5@4�+h�k�' R�Ē<#������w	����1M`��j!�.�8_
}#۠�]��yY���!AS%����t]���.V��D�I��T� `W2K��lWk��Y��s+G��@����}0�)�I� �_w��X�U
Syf�U�#YCCh1n3`)�2)*C�l��Ut�A�]��EaI��Pi�袰���%k��Loz��Q�S(�5�ꑺ@*�B �@���K��Ͳ�]΅
r��*0���� �p$���e���\6�z�V3`H��\c#�6��f��;��C;��:����F�S���.i��dP��dn	���� ���d�����L0�e�ur�= '}�6������xj* l�b���	��*����PT\fɝ#�J I��Tg	������\;���-��^3��KY��C��!�7Gz ��������{?�1�mna�V¿�s?vt
�(�FV�o�&�|���]�<D�D�r�9�*����6	Y-��f�d,k���痪�'��*������X�6���@����l�5ebs�1�Z�ZF��f��b��Kx���8]�!ޯ��]�
���\eߵ�;��K'���q+�m�$}���d��Et�u��q��^m��X��b[���6Y����>�͍<R�^���g���)��ܓnX���������>�}w�=B^� B�v�P�T��8��$:�P�Hx��N4�D��W7�Ͽ����2V�Y4&����|
 �����a��6��4���|��������_�3O�x�G�÷�\�STC���^��J=��VD�Y�p��	"%�R��-��z4ƽI9q`�6�Wo⃵e���2�h^���i��(O��+�h�C�#3���Uu�1��Bm���h"S^��,|�Ae~v!�E_��"J2%��4�u�I���Ӽ�ؙ�Z!w�����%/�b��j�f�&�n�öD�}��|:�X9d��%�=/���3s�>jdu�4�G�s��щ�s?T�+�̋��H�µ��S;��o���#�C��{A湞�G�'�h�}\�.��O�wDh��ѫc}�* �UXH������j�i��tC2��i��Ӓ=�J�������UYb�Ij�(�)sS̕T�X9iԐ�L��D�P"�옎W�3�7�,Ǧ�D�3<:�!��\˷)�(�qSd5C��U�`�f�X�%�YԎL��YGG���F��#D�T�6�dG�0k�AN"����}�Q��O�O�>k�aF��If���lv���{GN(R�0�1����b�tj&5�>q�kb��ҹ�WƲ�#��^%�H�a22�J����T��12VS6j�:��d({qL�/W�Ϻ�]���s�Sy��5qʆ�ۙ����4���0�N)��}Yxld�
�[z�,*�.���E6��3�gG�I�P�[�aFZ�gsQ$@�������U��g���r�U^_^�ۗ�d����MS�)��[�؁�;��kI�\GU.��~O4�f/��#ՠ`&�d��X2�Q���;��Gٮ�C$k*�
�e���#�$��!�S6^�*I<oc�O�*udć�a�	��m$�aa�fd	�}ϜД� �YJt��zn�d�ܔ~�y�����A�ģ�D�u�&���%��Q�ޣ����!���9�!Θ�����k����K��c���dJ���u`�?�)�\����M2M�˲����g���u<���*�L0�G"�9UE�{3����MJ��|~��)9�O�,��� a�����[Wn��o���7W�l'*�殡�>�^�F_�� @�آ��yw�M�l�eG�x�B�BX�����o}��n��~�2>����g��@ �J�O�ߺ�>��PC��h�_o¤3�~��zF�򰼌����w�h���\�T��>���/⤠�x:������r�~�(�W�Ǆ��$���r���K>����Н�Q,��	.�`�Ûolc���׻�i=���E�ˎ��FQy.ԉ1v�o���H�]-�C�3��g���p�?�J�}��~�BN�ԁ�T	�KMK�0�]��d�đ�P���M*FՏ�D	sp����2$%LY�1���H6rm��"�:3,�.{V���4�Bt2�1,#�֓���k^�Τ\eAN3��$�DQ섚�����M�pB�n�$�E��̍��qޏ�$Үp�/���EE
�lZ%N��0�~�C9j=j���K�I�����r��E�|c��l�z�td#Jw)�Nc�@#��xʓ{�������mfE�J3�$�%�,\7�G����R�J���O����e�F ���T��Zl�!�Ƕ�J�;����t�UL�$3���f��:ά���a:1� S�_����j)��%�r���5�������gږ�c���z�&Xp�Ces�ym��2���q���%~M,��5TnC�����^�T=*+��k<j<s탤�3N����P@�|85�T�u+���7e&��v�����NK�j�4�������ՙ�)��B)Ȯ�dl2�z���F��5������9�&��A�l��
�����\.�<��^�~���Z��<T�ɪ/ C���6�<�#3�ݕ�P餍\ϯ=�K��~�����!Vk��Zb�F��\U�kY�9KU��}��CL%�C{�1�7j[YՈɕ�*0��b��s6�}ԧ�v�{�r,�g�%2̖���X$��x"ᡥY�˹p1��,���*��켊��MNJ��J���Â�u.mH%yI-��Pzƌ�.�=��~xa�(xU�hL0�V���Kv	k�-�325&i��ྉq���B�cx|�}�+���Ǳ#�5� �UDי����i�J&Ő=�����i |���N���W_�W������ʚe�1�L��g��&��d`s����'O��\�3O������"���;��^����7OL�[��҄��m����ze��i��`�k)�x&�W�;�l}7�����(Tj(��`( :��)�o�wM>�!O8���1��q������vRE�����*��g�S'��\��ًO�_���Kĥb�J3�!M�t��3�K��' o�0kv�7z^<Wf�Y!� �PP�ޞ8�.^|	O_�b󠩎��ϩ��J=D#}�if�d��YO������y͓��S!��}������_�:j�{���:(�����@�̎���2#A����K��6[���x2*��`%H��ܙ���ґ�������'*�j8L:�Au�
�4�w��Қ�5 �c5ЌJ�&SB����R�#G��f@�����HJ,�U*��hK6��3Wn��_oˑ��!l�OJ�=��M T8�o�b���_ݎ6�L瀢u��G>+��5e�Y&�>�H-�I�z�i��&ױ�B�)v��H>��Sh�U̕�J�ds9]l`9&��i��/��W�$�^Y'����0C"�c][hhC�b�`�6�x<��d�?SK!�!��R�C���}��=���9�e��N H�� ���h���SFj�%������M�H9T�\FAKb7� �?���Ae#8���v͙�tl9Ț�3�BŔ�V��fp��v{`t��Y���},-�r(A��V�k�yHaP��960q/�%��^V��jE��m���Ot-q �(m"����gp����mqH1�'`�Px%���(�Zb#̔��Լr���ݾu#��>��}r�)K���c��Ժ㑂ʔ�ݢM����[V�1{F������������c8��~nQ�qU�g�)iʛ�1ݟ �gM��˱���V�e)05o��c�))��Z��H��W9x�V)�@�:�������o�ry��7k��#S�wmE%�h�T������J��� �<�T�Bn��)ׇ���K�|Җ/jB�P}�Y��
-b,��v�7󳙝��L���]��m� 6�뛎�J�IQ?�M,��m��W�S���f��Hpy��YE`���#~>o�NΡ 6��Q�ۮǱ�xL�Ƚx����}���y,H@���l%�8��M������Eܓ\�p")A���O>��kkXYZ����C|�wT�iU��h �U��P@ޱ�6���t��|����T�Q�~/�w��^~e_~���vp��m�Ů-��j��L�+�����v���M�r)Tr54e��1	�uܮ����� �h��~��
j����7��ux^l9V���&+r��7���1�4�Lwk��C�}���r��q�H=0�\J��WdYD���|�����.�pr������+�YK�4X�@�� �_�ʃ���)��b� ���2�޿��.l��g^��{"��@�� ��#]4;]�*�/,�����!���hB��@u��8rnY��̪���w&D�ДXj'pR�*�v�Cx��X&;�t���U���?_CN�4h�5�zP��m��m��Y��v���*�i��n�+疉JؿkV�1�F'(�H��x�E��U�ܬ3���(������r�@_�z'65�\�B��9F�B�6�Ph{☱L�!E'#���"�jC&��P�s��}���O$%b��2���:m���#̔�(b�����x%G�0P5n��C�>J!��v���@h�'o�Q���� �L�D��%9R�!�8әF��p�SǗ�ekf�1�_�M�?�9�7�m�oF��Zr��-�N��W�djFl΁�_��&C�/�ZU9�����:5�N<�4#�m`"�����ˊ�̕�T�	H�;W3摖	�b7�����tN��L8� I��06�gf�ƳL��AhǬ%4����΋`��jCdȁ�lb�b��P%G��.�P��%^�s��M�U����\b�\c��,�?��6�ސ�<�uE�Ů=��=��t=��-9���Qo,�sk�V�~Y��+kbW^�+����*�rɃ���Ȱ�Sg2iM"$��ñ^7���1sݩ���*W��(D~$��Z��,�3g�@��[�0`���wuv<��8�<z�H���"N�'@X�3�l^ө���2�ѫF&��=_��	3QA�Җ�a��NQ!i�|Pf9�zN	I�����yHB%��Q��?��[��l���hEǵT�w�����l�
;��Za�h�ze	�*$��n���j6Ir�ӆi��F=����_�����߿����l��H�-�m��'Knv_��^{��N��l����Z��h�{�x������W�(����t�P2&S�T03=�C�ˡ$����1o�f+�y<u�����[���O�*�)K���hd-E	/�RC�Z�j�|�'����������ON*�g����X*�ծl�z%�?��/`m��?����?�����������Ebv(@y�A��Wʨ�߾���x����4�����O������p)��'f�	l�8�J� �a 賊���`��"�,{�@�� �3L���Fr2++�ҋ����s�n x�L�����>�~�ޔcd��i�� 9�;��� p���řnȿp��1l��8f�O��-�%��\+;����cً��#��@��J\���mt���E�+_B�駱����y��J�Aq�ާ��Te[]4<Gu��b���͌�]8��McB��)i͟?��3i�Vr_�]1R�h�QR��M�R��U��PA#�x¬��fUD�FS���X��K@��P��\��-��������r̜A-!��.�~of��30;�T|��?R��7�y���Ck.�B�ψ�(����7���Q���rΕ=V�V�6|B��Oe�+��a;(�{�Qs���rd#���d��䁀f�\S��:��	��������3�:�C�9���b�ฏN�PBq�b}YFϊ#r��t��}(N�N�|�
g$���jig=K�II�d�̄��I)�j�Cd��3���g��f�P1�,k��0
�yqd9ՙ���}��S��<�\>kI�C�9h3E��J�hC�;�U�Md���(3t�E�����n]�B��a��� ���d���YB���V�����;��>��f\V��<3�&�e/��ܾ��~�"�Sm�1�F���tl|`�����L�q��D�c�E�u�3x����eR.4ٲȟ5��H����i��jv�kf���zbG��q;����Q3�SJc��v�o]��hoY;������BA�7c۽��/MD�ܓ n���E,Ԋ�RJ'4�E�4�qS��TΝS¢8�e�'d�Z��bZ��7��7�8�Z�[y�ɘ�63��'򓃮�`O�P�Q���ߴ�+�z�E��hv�Ӣb�]����N}�o��Nl�-��_Z�ɦ1ȓ�7��`*>ڑ�#%�:�MqKr?��p2b��
0�n�&%�r���p��,2��>��1�EF�E�j��A,��-Yc;�!R]ξ���7�r������{�;�À1�jA�V�*G���p���t��Ў9��ek�U����Cd��|���������P&?��?n�Q<���#�U���A���{���\���4�M��j��5��0�� E��/<{�\;g���e�-���;x�>&�ktf	�KG�ĩݻ�{�!�?�������8h���������������<y���kg��bT{L��:Z�LɇUГ�^̩��d�N���ٓx��'����ñ/ɂ0<-WX���u<���s�y�gA���>x崹F#M��rr���������>��Y��G&����(Nw�Ny���j����6�#��r���"S/�B���U�Y;��}����6�T1N�61�x���ۃ>���d{�'�1���d�-ڃ�T4&�5��#%�y6룎�f)�qTN��J�ah8P��c)v��&����d���Ȯ��M�+�'��r_������6{:�਴8;�G�y*w8�<�0Ejw�s��O�}�Y�"��t�\W���N��o4�/�g<fDi��Wby12�T�Xo&����M�K��I�X�8�e&ǖ5#TR�b�b(���J��X�R�(8�F?�G�R:@~>�la	8�W�2�c�@bA�~_��("($64��*���׊'�a�Ӽ
����zG�����}y�}6�]��G�R�t���f�6q�
 pT&�X��c���lFK��~5̪(��ם*�� ��(��/Q��V�<z��	�LQ�,:%3*/��L��nJeQBg��$X&�q��ZZ)���蜌��	z
����k��i���	w*q��s43��FV��̺5��|J��K�eF��t�IW��}��<&���͒R�r<�,���J���o����f��	H�pؑ="'�3G�
6��/�'q���DK�aG._���
AH��쏱8�QqM�\��B�:*��hJ0�88�ir|�>1+���l<��%���Գ�*$$�7!�3�����?�/�`|Z�_춃��ߖ �I�� �y�SEJ�ɟ� �����?؉�U�Ѩ���M�3VR���Wyj���Gͮ9��ѱ�R��mA�Y�G������,] �2���>˧��ѱ�GR��`D+F�ӱ�e֐�L3Ґ�z�ѡ��Grc��TU�6j���*�gl(xLTy�3A�ru�L k�&��$�  ElO�C��I$`� Ñm�,��"v:}\����^Gm5;n3�ze�X=~Jna���m��6+�R-uJ)}��g%�S-��ʥ��ǿ�k���^T�	%��h�c7eg�Z�[ҋ]����6��~y�7���;�/e�u:����l%���$0���'� E1������} >Q�ѡ��L�Q���ņ���C�F�p*>��b�{��'<s�1�s!�������D*�f��Z��g�YEJ��ljw��po�����;�C���bлA�� �RIn`Io^�Tą����ʆ�4t����=�������%����l��$L�qE�u��p^~e��.��Uu�P������)�\:Z�U��C߳=��� 5�9j�(�1+�쵷�����G�<���.vw�Qb��(.�K���s�� �1����?�kˋ��a�t��xX����A���2�J��8��D�ƱN5�I�l)�2h&���ݯ�Md�R.L��{7!g�$�!�
�G�_�����ٲ���~n�	]����	�O�f"#��Yk7��I멺&�R��� ��P�vE
�z�v�˻:�/�vuH�Z�J�T*@��j�3E���,��sf����^e1t���L���izr��0�ɬU�ӓM?��V֨?��+����o���X �펃���n��?�)�#q����6�l��)����1G�A�T��p��l%�'˝rz�[My�wuL�8��vq�>I:	�f�����Ϡ�=�PF�U��
;E�Ճ]����?�$����t�2��)� ��^`l;{gA��iJ>!���8�L'p)���@��1g�`9>K�9����^�����h�1T�,�K����[�}2k��>I��L�o`�6S�N�@�3#Y-���w����.6���E�̈�k&��=��df���t�λ��L�^l�<�
g�i�Z��|�z k�6zp.0�c)���˧Mג
��*&MA	�t�ˁ~����[����L~q$��ؘ����~��d�{7%��|ց��)���������ʟf��������T�*���f����$�JQF�{0��N�t���C�v�M:�9�z��PN��Ց�2��L�ƥ����Q�|&�O���6cL�E�8����8������iR"`V��S͸�� ��ޡ�O��v��)��C�?�t����Xp��MB��0�,�ٹ��F�tŵ@a�	��<;@���6��K;a�H�.}��T�:�8AW�]�'�'8!��r��]���Bg<�����&�~��Y�-40����}�h�5�*��,U�1b���~��W�'��]|��K�MT~G���Ʈc���d�P?��qf�_���4��&%��&��*Ւ�Em}�ZT��٘}ddO�x���E�i�]��/#/k�3��>�r8�\)xu���rͭM��ƖDL.���'g�KF���6���P 7��;��R��g��tNul��ޭ!��������Š��<�.���r�R��5w�4��>�����l��E�H���Z~.��,"��/���h�����{X�`9d"�&��1�5Xn���
��8CQ�7���e�UXʕ}| ������Y©�'p��m����bY����iA�yy���8��o�~2�Ѕ=��#�G���|�d��fyvG�kHͅ�����}�%F^���-0�\v�1�4e)%���#�{�h�c���G:���;�WF�)˙�L��[2�!�Y�d�@�Q����X��TL�%�����7�ɹd��R�r�++'���F��:�)�Dq�bz��ru�k�Vki��/�t<�pK���h��SZ�2F�)��� )e^86J\�\���5_;�i7�}��}��)�$-?�.��z�}1�v��U���4[
�i�`gk��]q�}Y�1Ni�{>6}��]��ىg�8��c�v�y��|^�C.tQ��D��]7�Q
<G����a���� �������^� G@)����Jdp�dQ���h�)q:(���,G$C.��l1�X�)�?	�Ӊ<q�8�Q��d(��ӑ}ڱ��x�k��)���R+䖱b8>� �Q�t���ӷ���?+�(S�;��H5��5��-�E�n�-gU�� �ϟ�I͒1���ϵ�uK����-T�e���H3�̭��k����!�b��笳L#��3�e�N�]��l���IPy��+�r���)QQ3{l���Ɍ ��0���*9�3p9Mݎ�y6~���O�*��7���Vp}А���Gt ���s6j��eUʯ����Y<�;}��T�酲�߸u!��`U�{��2Ui��k9y~������eO�t�Ĕ���%0e�ͤ�(p�4p���Ԭ���`���xI N��qTn�Ԧ�<���<'/ׯ�{�M;�4Sν��h�*|�CNŠ	8���Cw5���U<תG��w��$��rYM���,A���iD�i�����I[QdĹ��ɪ��K�/{����o�b_�25��hu����&��9�P�&I�o�s�uh��
B�C3�	%�ț�e �����w�d���-�����IX-V��q��]��6v��%T�u	T�j#^�̓bS�xp�>�i
�<V�b[]���0s�l� @��~����_��x����E��9t��l�p�����k4�k�2˞��_��t�Y�l�78g4
t��.�g�u�;����yo�\��z�̹���ED���n[�B�+`������Ar��)��yS%䳜����7S��w�/8�+�C��6�l������[�G�q�&q���1*��D1�-ި�٧N��(�+M��K�ڃ4n���F�b�4V�6���G�ְ�Í��F)�y������W�v����y��|�+�� ~��r)�{��h�1f�\ʠ3�"w�q�m�`e��q��àh�G��`��y�O���/_ǝ�(�R�r��tQ�r�F=$1�wM4gkT;���H�q�TYN�6�M�כ�ޕ?���&)b��1�3Z�p@�ol�,f�M��r�3	�V���M%S����*�9)���l��@ J"�8�|�r�0BhF� ^'������9/@M F9ˮ^q�Y�8���(eI�wP��T�PCM���c����g�:�!p�f��%���1+i�����]���r��b9��TS��0��)����f-aO9��4E�ݒf[\?Ќ`�MI_Pi6W@UΫP*ai�*c��*V�l���	����Cܾ����wqx0PB�^���n�;�]��U�p.9㑆����A��S8H0g�N+���SfA���|�_~Cq���{�D��H�v���p4��N8�+]��ŨMC���l��LK�+R_3�7�ZY�r6�����e�����L₫�����" cƏg;zi��KJ|̪��;m}M0��0�C�Kɗ㨠	9�i��N�P��xƙ��$3��\�N��F:�v��崚L'�;���ơY6
�I(��Ќ����@���|��	�=uBbġ66t�r�m����5BKޥ+v$�c�<[�t�Q%�t�=r�]��q���J�
&r����Գ<�8^��o`���0�G�76d��A��N�P��$@6��x8�	��
��:A�͟���W��P@�R5���B��hR~H����D��BF���|f�\C�a��T��g���ԧ)�y����=3��4��Z����խ�ƾI�1l%mh&9҄�r��ASC�x�3l�V�����1�m�K�?#u�G���S{�Z����IE%�����>~����8P{���
_\[�g0KY*fb53��yh))��M�q��Gd��1�j��:L9�S�=�D��賒��Y��l�öN��V���;��붴��f9m�[t��i5Ut�l�}5�SڇF�/ΪV����Ư�O�������G3ݚxx���xV���9��dB�y�Q[��O
f\���I�3�m�����+/=����,���ܠ�W����H҂��L�7s�s5��]|pW0F��q	�6Κ V������/���p�kg�dJ%��,xv�䴳�����xr�㹃EܸQ@����|V�wL�瓈P�ᢿ���']ș��2V�X=qz�O���{�����:����c8&����8���j	���}8;5l���� ν����)��#F���q��/by���kx{{K�8.�  <PB�H���FC~�:?	�*r�G3Ό���]��I��$4�\���c�hh˙V�A���~�1
�Pc,��8H�_�r�.�M�'��������WZgzb����,j's�l�Jq,�I�HC�Q�2�V��j�����3AVr1T3����,�)y�ZN+W�S�����,?yQ.)��;�ϪzzW ����s,���N{�V��Q#M��%j͹�Y���H�h�12C�#S���w-�f!�bwš�B.����8m�~��������P�bi����,���p��Nl�`�B[��q��=�lu���B
7&I{�ɽ�\��5..-�!#�,��"I��ޢѦ2Ƌ�CF�99�ݻ����_h�����N�T��~s��v��|�l�"}G�;3<�1���ຉ6�L	�+Y��b��7N0���*
��t�0�(�Y�Ĥ����2"_"�G b��W~p.[V0W�,@M�+�W�R`�����Ĕ��5rM�	��i�����Qbx�Z�����u���{��i�q�bأ�m��q��X��x�)���^3St֮i�PG�4&�����O��a����A���fCy��*r�9]Ay��cY��6_���S�&�	t�{�<�3�c��Ϙ�w9�,$��(�-�l�0|��<gx�3�s<����lKy��8-~��Ǹ=ŤȮ��.z�+5yv��b�Ƚ�hv��A���5��N�z4��(I��f�J`�9��T�Ll���ihj�L*��#{C��~�ƾ��)V*������N��>�f�d�������rOi6&��+*bc�1,�^��z��tf�"� iu�;- ��݉�5��0���é�w��ڝ��!��FN�4����6�L#r(��5@�MCj��7�a�$ɍ�&0B��_HeN�
���^]��o\��ƨ�%{��\����6n����Ԍތo���`�B��o�;]�B#`�@�8y~c>y��~_z����Gx���p�=�|�wq̰�y�@�{;`�̄�v�Ͻ���H2���4C��>���������L�h��K�j��
Ŏps�l��aR�T���᠋7?�����g�~k+3�>I�]C����y1�y�3�0��� F �i��D6�pSd�ӫ�ᖐ�7t���f�6IV�߆����'��w0�ʃ������н������}����~�w��N���ϝƱ�%<�rMG����q����o���ɮߔ�#V�R�M1Z]qT�|}kK��b������]F#�&�&S.ht�F��?���$��#��O�D��\�E�N#��։k�naU�d���_eʣ�*r��t���1S�a򹮙��4�k�L$�#Pm(3�Q	��N��'�[�3�;��m�=2�A��og�J���!EE��T�Ȩ�bY@Q>�F�aa����XZ�hv�X�O�jv�A�C��wp����fI(as�00P���kY�{��~����d@1]:f�Ɗl>������8�B��U�w��f�-m�}cm�3���h�2�		�ʓM�TB��kb��!�\@�+1���;�&��������q��Y�c�������N�u0h�#�N�d_�!	�L|�	��n8яL>��:��D�+�J�o"/F{ ky��V�ͱ���Mk�ɛ��at��g���( |,�-3+˒ޕ��'r�p�u�<}Zg��sF��@��Rf�j�(rK���9��#%�������[9%���BuQ�������=��B#��.Jv��F����N�%��QX�D�/�
r��v��F�ڱ�����uql����mܽq�F_�~J�,��Rr�Yvdc32�M˩.Z�M�Kρi����@@σ�[�ܺ�Hr��Z���	?���%��]�M���I�	�e�z65?��J�k	f������@�%����6ZZΏ�]��ܽ����]P�����e#��?����1�����V2Aؽ�]8W�E�ZD��a�TÕ~S��,w�䷎	x_���ӅJK!�匍Y]N�X�b��Y�����̜�	����:%j��
�
V9��?�"+�L�]Y�i6��ij��Y��/>j���NŁ���Qز�.u=�v�^�2-a�"!�X�g�YF��l�LY�O2��&'"�G�y�\��x\�r��0vxc6٥ȉ-;�)��*?OG�y���_蓣�l�-I�w�?��L��It�⩙�-kk:� ��~8~R�-	�����K�$8`ƺ(kg]CZ�˷n���X1�r���ə `Vj({�Z��7��|�����Y���$�Zӏ�����X.�?щ<5�E��ǁ�Ǳ���1e\W�̂o�K��^�g:���[ǆ��M�t���l6/����T��Yk���^�]����`ii����T�d�U̥����P߫���`Z���$oH~e�Ź�ϼ*2���SQ��x���J�<��}R��=�I����7b<z��3VG��9s�<�~��8������X"�*�}�*|��/	�����<����>���nb,h���ˎ8���0M0�\H��~��x�s����u<~z��-1xbz��tLZZ6��]hA_g3"+��u$Qr��r�	e�J;���nhF�m�j�:��V��L2l�IhJ�0@�C�9��Y�);%2`'��pj7Ӌtt^NdG\i�6V�
�2��q�z(�B9�����9V���j˕��+�N��Q��.��P)����iq����v�#�W��0�x-�y�} �{��8?%·RW뮦��Uȗ�٧��w�w8����9.�_Φ4�E"19EqU��r�	�}+�ˬ
˒�Й�#�N�'�e:��ۭ��P��C�Ӿ6\� ם��i�?y�.��P^ƙg�r�~����%���t1�0��ۚF����)�U��C��S���L9�+�OM�S7eWU��Ү���P���ޚ��!z�f�h|2�(w(�P۬/������|~��vK�E�U1��j
�:��ΜX�g��}��5T���N�C����c=�H@N��:?�#�*�cXZ=�0�-��+�ԮY�)pC���Y=�Ŝ8"f�i ��0f
UzD GA�r�\T>�^���F���G��0�Q���$��Z�u�7T}���e�J��9�̯ka�a#����2�:�@)+_'�O�p)L�4Mi6��3c匴��	G�-P��x�L��Oj���i�P�_��g�n�N]vhf'{7�G� ec�����=ܻy�v�ݖ��S�a�e��g_y��U��m8w(`�\WY�̀�ٺX+����2N���&�"��D�CQ �Yu��tt�����
�X�~�f��i-�U�A=�hy�S.܌,�,j��Ʋ?���|�\�#�l��3��9�b�C��eՑ���S�=ʸ|�>�:ع18�s�V$�+�} {��1�OI���6q������33���V��$�J�P��R�F�o#ս'��#3h@�y��?�d៸7�n��� ]�u�7�'��,��L��XZ�!�;=*s�\��ۜ��u>v`�䂵%�	�m��UW
ɝ{�����Bf���j����!��ZU�a�'*�)�{6���׿�|��KF���I�*�LN��Z�����ǏH1i*�#k�7
�/�:��c��w��5�V��2Ո�~�@��r���,�>���.�w�!(�ZY�X���˚�g.v+M�G�%�~f�/>���������H�>ȧ�Ά��5�RVd�ā�A����=�ˇ���e!{K��P��o9 ����?�'_$�~�H��i�H73��"��g?��M(;�~�>���5|�O������|��Ȗ�ь���XEm{r�*�>�]�4�S�lRo��>�X���%�&gU�n,QC0p��A-yKr���]}�J��G0I�(�A>����	}�	Q�cd����p�'�H<C���br�ڥ
�lϑ64.��ٞ���#g�dm��kl~���~]F�#y����g��O7�z 	W�8��YJ&��\�'F8�Z�r��bX[�`]"Ǎ�
N���T)����ܿ��{4v�h��^�d��J>2uy~�JAm>�+'/��u��PJ��^:�K6�iF[��y����4�`�1�Mw���|FfRh,uf$�@S�t�����~sT�D�WvmKd7D:"����`؏q��%׵���[?� ?��P����3pZ����N�#{{�6��u��@���q��2�ԡ�,���g�4�PϘ�G��u]������T�+�xZLĀ�0�.�{��9����C�x�q��+�(h�ѵ���}dN.�3�}����7�%b�|����Ψ��X [�uG�Z�?gh��:fU�MI��a,�=���R#�S��Iؔߟ���TK��&	�ƣب�Ob��Zn��2`	�î�N?��ǟ��������?|S�v��9%G�n.�)����
���9OL&wvD*�t�3��d��|b�TX�P����t��9隄O���Q�-y��`�gĦ�|�bM3�|!ς]�Y/5W���=f����>��������GO)t�|X��]X��_� ��wpZ�'�L�]L��E����P�����զ���-���(?X�h�0��\ ]!Z��lf��3yf$�G�}�˗����,2��)�l�*r��E��e��̜φ��!��wt�M��H�ڣţ�Rj�����J�	F}ȊEy���ro��bR���\���{*7	b��	���9�Ve~���(�aO�Rn���D<�= �$�5�Ŭ�6w�1;���})��@���T�Jqѯpv}h:?i�f�e?�5�G],�M��q�'�h�+��v�/[A����Ԧx�Q�I �)S��sr3��^='�������검W��|�Ў��;�ڝk;V[��ת��L���I����<�����|gV�X�LS�S���
�~���F�T���jm�L �����������?�p��]ܺ}O�=m�u�
�$o�:4C��%��0o1��\YKj�:�~h�|(a�º��8��߳���l1�C9����RM����zo|�;��O��W_��^ Q� /}�E?�����{�G}��"r�`'�D�b�,;YY�͟M�:X;ߍі�q��m\�W�|Y��&6�)�}G%Z���R'ħ�A��δ�ĝ��Ȥ��5Z\*CaS'��Q`G�SGQ��ȝ�Bxl���ٴ$�sp<��NJ�cN@+�C�8��*B�\�9_t8�Sr�K���5��9�Ô��a�{��W�#�l��r��H��T^�|�b�|�S,/t�����J]��k��]�����+�qㆎ��,�b��J-�2F!?F�&����Oey�x)#��e$B���%',Te�L�SNU�O��Rz�$��!���*�P{�33l�@�"��QGf�JcH� ��cɑ6�'�`P��'F���SR�e1�c�Lv���{�!7���)ag{;,~�w�z�.���WU�a�VV	�<S��z�)�Qc�@�z-:1klρ�fcC�yJ�.r\�4<A��|���U�?�*��<�z�{��geT�*���#٣_VDU֍/��psK��6N������-�l��ɏ5;�N�����XX^B�^U��n�:���EK�O�Q^�q��8m�����T��v_Kϝv=���Z�tq�m�-N���t({�o:O�PK5qXQ���k�6�rm+�N���~�P�	�Xr�m��E��)�E��~o��/��ӹ) �� ��g$P8k��Vm6{�42	�ZFU6e�R.�Σ���Mb���R��\�/E��/g��@׎� e3�,��:���\�Ž�����!�z�U<�,�U��D��_�o�t����g7�zk��d��f�k� ��a�k����l�df���;hhu������c�5c�CFGZ%�xܹ �׫c'�@;���}J�0m�	�m�{�ʐ�G�r��&-L�ׁ����tSS�I���P�uo��o�u*@��
,�;%y�'�oȒGژ�5~����/"�,k��:�b��癬�`fj���Z<# �
w����=�}�
ǐ�����ꚵ�D�m���Z��N��J�0RW1��<��4��$�fQY�����7K�1���o�/h��+��i`4�G�&�yMhg�Z]�gY�I�����O�d��se�:Vg�a%���k�E��o�^~�" @��2��>5��b?��ZԞ=ʿy��ʩ�Y���kh���s�R2�6�a���jS`9ߗ�Q�)�{�<y���ｯ�6���o��0�Y;6�����p`���q����ǭ�p��i������v!#$N���K#����v�DqF�8��L���..����P�/^�znRW�	\\z��9��x7�ށ؄�H�|�\�$��'�TF6�䘖ZR~)�5��{�gI
H�p�� �I���[��=��D
���˟,��8pMV$T��g�TA�ح�˧f��ysQ�a��H-�f}���G���O�����{J&5���\�+��F����@w^�e2#q�9�v��G�!*rM'I���Y��T�Dٮj�)؃)��� q�p�5��zh9(���+�����X[>!ѵ����l��l��<����8���:��j����^�Q(�*7��?f&�l���r-|T:Q�M�S����C�R 3�ʵ��PM8L�W���̈Ί����L���S1����D�Q�7ݗl@���v�ȟ!�{���_R ȑ8W�q	YG�n��L�N>qBK��;mܸ���w���?]�lY�����+y��c}q����*�q��ǘ�y�\�L]\��sk��qpZ�2A��-�ִ?�5���6�J���nFB�e�XѱJ�|J�n_tC\�&�3��ǱۉQ�TQ)�U���/j�Ѹ�gC�����+7�e�g�·֎�"'��9�JJAA��D�֘�|_Fwؗ���5�4%  �.B��b�?N�V��Hf�rv�;�y�>��*Z��r4Y�]��Q��}�c�!Ps1���7-�R�Ζ+fbX�"�O�GH�m��jW2;��S�UN}-�Ŋ��<�h����X�43��z$�P;�Yf�A����C$i����2:�4�����Ӌ�;�51��`�HX�Z�k���{�q������:��]�,;}iI��m
s�Sl$ο?��`͛�F�>����9�����j0�\K1^Z8;5�X�pW��X�����>'c�ꉽ��N�s$�A������w��W"nm ��gq��6%������%fC��ݺ�Q�%k����5p)�Y����8��1'�Ŭ����D�Y�;�����*��	�_Dܕ�mu�ڜ0V;�ly�)g��Z�g���Y��][��L�#�j'a�%�3�B�d�^���œP��j��|�1mAz$��Gc[l���(bem�׾�,���P�����T�	.��}j�~�u�;�{�'bƲe�O��5|�W���rmO�CӘgN����9��_��VG\�d��2J��m4������?!�m�����*\j}��ZYZ�gN����wؕϨb�k�`���U`!(v�_LI�(�m��({�~���W�NXQ&���Х�(3�GL.�b0�iV߈�_���*�\����3�YUf�*l�����i�%���K��<12�Z>�����8��3N���Q���[���w�hv%��;���Vp�D�����o.��0��2H*�q1nK�����T��{�<h(/j�X�H���n_u��#R�X픆�8�/�?<t���2}"�݊��(؀��Qn��Kvu:E��Ӊ�8c}��'����ӹ�M�iVɜ��4��k�1¥�F�wa��8��7�E�����}Rr0��sp�Ј$jL�P�����bD��q�s�C|�fn�u�D��¹�u,.��P+)��\_B�XB��G� ��1CS�� ��>��	��*����i����"�|(@Uz*W�{�%��0Ġ;T͈��r01�K5�jS�ćZ��6k��E�#nf3(G3��̌�W���+,/�/�)�L�s^��qy�)�=�7'pw�(��Q_)�zu[���}���cJ�__�"-��y���KX�.>Yݜ��\c�%0��`��)��	*��2�h���#�f�l"`����A� �
sy��"\K�"v��p(��2DW�tG@Cq��}y���3yx���8�bZγ���t9��v�:��$�74C@P�3��y��l�����F�rS��9�������m�m��̐�'v�%%�B.�t���N�޼��b�	��TKb+r��.��F�$M�*������dMb?��dsb"6�q[lAE���:b	U��SdO1#�#�d�Y��H�����������H3�=	�!�S	l2���0f���B(���	&2�il#Ne�;���o��_c�#t������u����Ԗ�����hJp�{���ݎ�s����jk��^y&=	"��	Zj����c�xA}I{,]��۳�O˭^R�2��T,!��(g��kGnV>o�Xޑ{�Z��t�,�S���� ��Ha������_���+�BZ��#���،)�ೞ<�Uw�'L��]��OI���eT�;ȥ�7o�;��¤!���v���ttOS���|D*�ǁ(�M�lz9�v�������$�)�1�.`�u�<𧻓�L�m��3�l�f��7�×����9��'�:SBĬ6	���D-�hҕ���-��3"u$��MIqzC�P�xQl�˙��H�Vo��YK�<uI�{P�榏�7���i������agG�GjY��6����P)g`��ugf�Ƶ�~�MA��p¼�mr���gs�p����8�HN�R_��-�����?�^G�c���2�2f�%����<���<yf�O`����h��%��L"1���^A%t�Şi���9R�x�P���u��ϠT:�SC|*�j����{5Y�^Wb�s�͛7�/_��A� 8$Di�	�&b�#>_�0!E�E�0
�B!ƌ�C�р �pmѾ��WVeV��9F{���[��&����HdW���|���^ۭ�$4TY6\zq�5���3s1���cx�#��,�$�cT��צ�$/�.a8۪H4�V�wW)dr9�Ɏd�ʁ�Ø�
k�ת����Z:$��T)�-�F��k&+Q��3��o8籐�g�Kc�i !`i��.\c�b��V<�'�G�*D8���Ό��_&�5.�:�0�Z�
Nʶ:�e���)B2פ~y����ςR���~��غev\�z�(������j�1&ǚ�߸8���0-@�Ƈw��]C����,Ξ�ǪD�K+��JI�\��� �������{���5W�_{m�Μ�d�z�vG3��C�R?T��`D�A_A�`�5f�|ٳF�����U�\�`Sw�L�Ȏ}C��� e��P� �=��}a�]A^!��8��r�sS��,Mǐ�M"6�!���B���)��+eq�������-��>b���8=_�x�v���\r&���C�i��,VV���I�l8��N��MG�N��<�k��\y� #�$�i���6Z���M�dk�	���4��x,��z8��J�$�������ߛ� �#�aV�Iy
��
���:�ba��+(ͮ*{ �6%G /�;ڽ}��a	��`�#���$��wG����@��5iZR�*b�̕tg�Aՠ��f���8��*=�P mO�N��1��>�a���15���[~Q�oQ�
f���a�:#��䳇��{eHys�iĺC{���׀��2��zW�=d�y�G��SL�I�=��3�]���%��?�Y�b�����fT��sGx����ʍk��k���-ϢI�eY�cg�<HLƏ~p2�oO�?Kw�=j�Øt�v8I*�p
���i��ސ�M����_����4G�]�Z(�J��8�è�����V�w���I�Y�Q1(�*��`N6���*�Ͷ�v���qX�a��ǂتiY��Úf�2���WE=�ҋ?Jgb�Vȗ�R,�Ft��q�_Ø�NF���X��'�KQ%VIѭc�`r�+��H�G{J�=��(!G��(��@+*�F�,�o��$Y����I���T�\�j�ƪiֻ�)�x!���Y�;s���՛5\�5���}\��D1w�>��\H+L�E�c���>�Ǐk:Wp|�p��u.ڵ�T�3D�Сq�N���2���'k�v�?t�	?+��RI	Lή-a}yUR2�Zeſ�^K�ؚ�>^�q�b(v�C`���̼� {��X^Z3�T�H����4h�1��	o�@$Uj��jE��r�c��-���h[�|C'+���$��G�hT-d�f)�������8�����,��+cu!���o���
�Rr�%?��p�#l!/�r<4�1�zK�p��[�S*���+���Ҥhw�qL�O�eE`�l�㾓�&^��Mn��,V��g�a��¦e�Z	�87�O���O��1�|ai�@A?�{�����LG�acHd����ha���v��ģ�q��1޼U�ݭ��nk)ll�S��P.���|8�y�Ħ�%
��
�;@�Z�PU)��D�:{�F�(ߨ�U��B����b��$�@�̜��Fk�\�cRئ��i�֒sĥ$͞2�����`8��乁�����XA�!�*P��Jd�0�,��L��5�l�`j� �*�X.�Di�%����%�2
�����*��x��D��Ԇ�iH�B�%�6|푢#b�x��\��fFW�����$�&��0����L���B�Z��oli�'#��P. ���Ý
2{;�=>�$��j�U*��GB:7(�!K��BF�IN^W�XF6_�!7��w�*�͌#����1���=��
�HH�>S�Z����W��hԴ��#g�Wt�։��f��L�"I�V�)�3���.j����OZ/m����F�I���r�	B�d݁����i,��~�����?��8	��洶���0XL�Y�Gk�2�bK�1vo_CO���-	v�d����~�>���)��˿�˗����W!fj�㳟�*޸���Wo!%�켛Q=�1/	r�s��Li�fR�e�~�iVG�W�U5��JI,��b��e�z��Z�f��e{N��N�����l���C�r���X��fL���>�xjZ�_
cj��6Q�]�}���!S�C^@�߮J ���!&��.�`W�\�px��)�&4�G��ںc��W�"zT��I�l����6�>~œU4ek��R�WmXB޷��谊#�t${��9/5@4��l���GM[W8�#H]�̔j|[�X1U�ω܌ �RyY�� �T��)��k��w��,�-�y"#��[��杔؂�x�5SV���+,٪-N�>���?�҉�2�����Pa@��c�3����$O�f����Hcmeg��q�֦ ��R�91#9���@�uL@��H�}��s0��M�#sG���-p�>FZ�}S>�p�4��Hk;�w���÷�P9J�$���<[�G�FD֏o<���51N.��@4��Tc7W�ǝ-/�|�ݯ>�_���4��sO���Q�G��p�c1����)t��N�τy����J��Q�ă�a${}��HD+Q	V�~7� w�TG �Q9�?%F��OC�k�)���a��AJ�D2N�F���'�Y���ч�=2����8b��x�����9DJ]1n���x��x�.��� �]�=��3��_,i��c�K0MG/@"�A����b�ޡf��7L`�m�����(Wy�iZ�յ/�I���@� ���%�M"� P4�qq�l�p���S�Ǎ��E9�lxgϝ�Y���2�o�N��=���@����`����i`_�c���8�A����9��
���[���b�gf1[�;G�����9LIL7+H�we��z���P���w]1���C^D��V�a�K�]2��Ĉ�z��o>�o�Ӻ�����# m^�����LV�Rܩ����,�oA�)^v�j��z��A�&��}t1�rϋci`�������x���|����/b��%��.�k�Q^\��',���	�i9`���s;<<ĮX��o�������N��@�4]��j5�7o�D�.�b�Ph6j�,�������?%_&-K����MV�G�H]���蜇Ό�d� Aн��O^ħ?�y��po�@�}���8�.>yS3�b���ʾ��ҳ�~���wQ��PE
�L�BgΞ����&�rf�)�Q[�	3i�%��Ņ2�������C������h܃�r-������Y�!|&e���'�f��.������/)46��1+���r *�L8���{��,'��fK�体��Tq��)f�Qd����Ğ�7��>Je�Ĥ$�lK���JB������X�'6��'�F�4*R�+n1pM���?�=�dV�m�Z��`ש�;+�K��������7��t���'1hb�d00�`��9�"����-46I����kW���a�!��������L%�J�WI���LW�,�������1W���y�۳�=)��*Þr�,�#?�"�9�����p��i�[~ԟ�8���|o��䈥-l�!_*_�6�O�g���@���SVg��!�V�?Rz2�v����of2��&��J��s�׬4z�U���Μitr�-&9��������1^e���� Ϲ��g���K�FٗY��f�n�IG�\Ǵ�p�eXV�f��@���	�֏��O���?94���|����X��ut����/��
�W����ӟA:�����TY)'���B�wG�Q�w,`����{�{h�|�q�~_K�:m3r/;�(ʐF���9O��3��F��;�N2��E���0��F����R�XڛC�L����&ʬQ�%�
��Tc�B�F�����<�4Q��3^cvE���s��/���p���`k�xy�Fy&��rVS:YPʙq�E��WٱV×`�aJ�}9`b��0�k<���r���}Uň��+N����e�e�i������8p��8��>V`�=`�XčTX*[T��^;���i�$�M9)zO�Gs��Bc@PA2Z_�,����B�IB��=�wyؿ��Ý}dr�Z�+л��*�y[@�4��G���¼�H%��Ƚ%p���t���z��-�%�������R���Y�Ӂ^|�T^�̵_Fۃh]?lY04��1ɔ���z��C9K.��y>�������}�i����s>:Z���E�P��~�l�H�����b/� �����3��8ǽ�f�y��RrF��-�aum��9�f�h�����𠦚�{�5ē9ܺy���O�q^��3=�-m�f"�}x&4��,l73�Qפc�t�՘���9Jp0F��a�S��̯�7�s�{ؽzk��<��� }fE�R�rr���A��E,��_����?ǭ�Ѿ�Ď��7vqyf�򫿄򣟖C8��w����zr��r��f_�[ܵY��q<��O����x��>޹}�psԂ/`���y�+�|R,������ F��NI4R�t-�XB�ZH&�l��~@�.��f�	��c�A�=e�D!�YV������c. �EN��8\ǿ�%5��	}�A]5%������X�]w�AR��ΰ�ٚ��=��~�H��s�.�J�	*s���a�QS�N0�� 38���%��	�#	s\�c�hI�]�*b%\�؞��*m9�$z>���Cy@%�A)��f��M�4�|�����E����/�;%6lJߗRI���֨P�MF�,+>R�k&gzc����鄀_�WhJ���xF �P�F�AV��3����9��a����{���̠���������u?O�Z���Z���X��9��'�2	�/ڧ��u��8�nzB?Ǔ}��l�PF��y�ik���!���z��xZ{�)G�AF��+w�a)���\U+1�(d}Ԕ�ʡ�CA�1%�4��j/}�.�-K�q|�K��������k��On �8G�E����N��@�b�	Z��N|�C���Z���V����}?���167�?��=�N��Ĳ���&X����N�:)Ӊ���O����r�=X��u�����S�=��@1,�ZFn����02d�R"��4�����&S�7:�NrwM|?�\�M����|���e�.�/��e%�~����Zx��sx�5,�e��Ő�L+uJ[��-qF���%�ݧ,ِ������(��9��L�d��_�z���h[��I�L
N���,է����`&l���Ŵ�F1yKu6a�Q��¾'���X�N��7��k�ZO�d[�+��G-�~��*��Z��R�v�����j۷+�߽�+W����U\�����d�8�4M��tO>��N�4{?-U�` b�I�wdG��I�2��xu�� 4�����'pF)�������D���xVV5;ԑm�*aٛwXE1�����>j�
c[��9�ĩN�q���"S�!%����6%�x��� H�$À#P1�Ȱ�D��i���IjMB�AO�yM1���=�5X��:���}���ˤ�$qgg{�ZS3;�DJǡƩ�* ��ό��[��u�%�p@����AN�ӫjfL'��x��������x�C�g���?Ìؕ��|��"Z��3�s�p��$Ϭ)��Q6�W���P�Eo����A�z��:���GJ���D�7�Q��7�����R�BN �m	�~�{G6K�X�:�$����|����M_n��}V��᝴���cT"b!Ӏ�!�ii8(�9Ik5 #q�^��=cou?�x��A�:�gNξ� ����*S&��l�Fa� ����t��Y����7g;�V(��\���_��o��Ⱦ�o�L^,�B�PF@��3
~�\p
�E���@ �Xem��s�P#���԰�)��#2>��jĚʝg�9I;�s����c�_�4���C9T��U����'r����K���[��d���}�]y�C�������r<�+��I\�%&��A�<6�|��$����.g�ίV-�83����G�����V��y:&5~��ǢA���b��=�J������]�$ [�t_��*�u��/�	��))�h �OI BnDWl�۔((�
�pL֏��	�˞8j���68Fg2��x�9}0�I�\�[ox����h��5|����b��;�e<�t�<,�U�^�����I ��Kx��Z)G˽/і�-���w}ܺw�t����.��Y �b �t��e)K �r@l4�l���0-N2�L�a�w'ێO������:?j&�����{;~m�4���̇�0셆�t󏻸]X���Xh�����]�8��|�L񏨼 ?;\xh�x7�������3ϟù�2S9��cԪC�mUq���oVШ�L9�C2l\�� [2��,%J�	��Mg�sҗ�8�	ܤD�������D:��,Q%Sy͂��Y��ʴq@Dy��0���<��faj޶�DF�6���<~VmH�ZTPI�c~��x����여�@������6h4�+�����l#�@�Z	и\�����N=W�Pcb�����)m���%ĳ�	L&�� 8��by����� Ҽ5eQ��\��)���tqB��/6ݳ�Љ���-d��\NA���;�����5' v��޼�t1���UOK�_�cgaI�k��`q��D�=d�i����� ,��lB�h?��J
Cղef��S�GG��bA=Z6���:P)��h�\�������Gm߹���3��q�����B��/^��@t^��m�mmV4��=����1�K����Ѿڞ�8�d���D������m��EN��c�����2�>�SE�7�*h�%�k4;���>�~�l�x6��Ⱛ�4�޿�~�]E	@�)	:�&kBm_�T�0U�<���#�3i�gp�v��nMqPl��C�Ϭ���]�۾<��o ��~cՔ%�d�u�u��:I���yf���<��v���f��A8K�I�,Ͽ3�s��mT �'���P8JD7�N{jm�T9�?����Mq�l�%8Y���Α<�1�3���N����䌺G��e���P(����)1�}�G?�r5��]��_Q����
���za���k�ҔJ�ҮܫJMz����P��g���(���$��+�a}�q���/���W��.�=��M����W���$@��� ��ؤ_��a*ncV�R��t9��z�x�A�9n&eꋸO�9m���P:)��.�! �OZ����l*�1�4({��tAv8)A���ˇZ��������1hH�t_G��D7'�IԔs���X\�_9J<�l5�;�	v��.%i)[(A[G�U����<J��H�:�W�����UK"�<�d/|fEX����E�Lo��^�uQ�=yL��Ⅵ�O�2��N����.������8>��g�jVp��c���wvqW@^�ˋ��,�-ۻ�A�n��l;��1Q\6�F2D��p��څ���9%��Oi��ŘF.�F3�2�W2���B0u�E������w{�'4�U)S|?4�a�:���La�z��k����D�K���m���]���������)��r�U�����s?�"�f�j����:�y}W��D堇vm�t�Є��d�cM���|.����	�R�I����t8ITm��Ӱ�Š'Bc���NI���D�0
�8
�#�5~p�%��p�4K��8:����ì�8[7�t��RQ���aFmO��������1�b��9̻6:��v�h�:
T)߶?��M�+M�<�m������b���Y>�`�7h�]5Q%�z�fo�����9�� G� <fF���}����f�;n�B
6��G}����8�^��S��X��g�-
�8v����Z�LA�U�icY�����ܫ�<5��;;�}��r~���ѯ�t���h��eL//�	fY�2$l��*�`����Ҕ�f��e��ӭ�;�7�������8��Z��)�3�dM�n���W�쫦���؏B-���C�����R-�c���5B���\R���z�.������{(P{�#�t��*ͰZ�_�a")��g�����_�*�*]|���rg ��� �Q�������e|jc޽mq�Mt�y�]�פ�p.�Š�����_�'�����6���6Z	G�V%y��J�!��Kg�u�X58�;���T(8�������l��sU�n���ݶ,�<�u��ٔ�u�tٳ�!+�a�M
����[;��2N"d����d���G��r��ѫ0�����Z. ]�@b�	Y�m�`�ykUy/�4�4�'��-��Z�7��ߵ�a;CԲ���=�&;7�� 8����Ț�ᦗ0�t��⚾�/�:n-2�&�w� �]Ni���pa����7_��~>���-ܸ���G-�
�H��4�nL�{��y���յ~�v���E�8�&L�G{�9 'v���ϰv�m��e�C���x��V��Hė����Ӻ6+W�f��j���]ʆ�.)��e[�Gg�~̰K�����f�~2Z՞?m?���!V*�~%*�$�L@վVjU��x��x��)9�.�ܭ���TNo���W���9��/j_���Ͳ�L%N���gd��#�[�!.^�k�6��ޛF�C<�W��:�����i���sRB��=r�cѓM��/����&����',�X�I��,��n���������O?��WF�����/�}��_n���y�
k��U�=9X2��< K�$3N���
�V�xZٰ��D��z�
�mm.fs/����/�5C]e#y�)Y��DҝqG���E��t4�=��`�:㶦�G��ÁD
�H9i�������X&�Mu���f���$���fn8�i�v�2۠�wRA�>O+���cB~"f��W�u�%k�  �����Z5\��.�s�_���ńNP�=�����u|x��8����3�m,-�1UrQ*�15�2 ɓ����B�I�d&2����`]c�e!M:��S�p-R�aE�x�b�n����4sh�y �����z*���t�O�|ji�S�@�|�~� J6�$(J�	��+����s�{�F#�Uě�H�Y('pQ���}���84�����<��9�=����HV�&�7d,��~��H�mY�]..��jV5�{hF.���"�>؃�����ZUQ���78��c<�`C�_��8����U5�֕W
����+������{�jt��JP[Z��	O"���DM��'e�ey�W�~]ֿ��Ϋ�Wsp]����}��JE�{���Ԉ��ʀ�=��4#-������]%�f��4�*��h�͞� �r�W= ��k	��NF�q#���l� L�,��,�DF�����S��t\�GZ�#���IY�H� Y^�GS\��`X��|Bl�iO�{��=X��/?������8��������lߒ@�-�`h�p��n������H��+�qH��%�8������4�3�=l�W6�G[��ZU�^ڭ6�)��ͯ�DY�V�l�&9&�Z�$���\p̑���PF���>���m$��.�A![ĐmG�^�`�r�J/$�9>I^�qf�<%�֢.iOd{�� =�����<�� Eyϱ���

�>j�ޅ_�+�#�@�=6�y�҆�9����i8!�s�8sbr�V��Q.�1��I
��>g^�b;O{���x�F=	��%��=�~�H֞��)�mɽ��|CU��}U(
�ڔR
(��@�'AH"=' O֩)�<����_��~y{���ի�h� ��A��e�'�خ�8��X,����8�Y'���[��Q���KPU���BV��>RS)$�y�<-����h�¢�7�vK�9K�1��s��eȗ���q���$�T#wC|���	�BUVl��%i=��_-�A�wܿn���&��m<���D�f�5K�������C9���W�{��8�^}j���giS�u�HJ���N����$ͯ�*��6�^`HM��>���}n���^����}|�v�-��x�pf��¶��I�?��_U	��MӲy��'������o+�����/�iK)����.����O�4ÃlYq�-�U�b�gi�f�_�������{�GJ��+��ѯ~S��!�tڋȮD��'%�:Eƈc F���R��?�}�a�h���	6)KûG#�=w���)+��L�$͊NU�up"l�`�2�f#��0���"j+T����a�#đ�_��ʼ�k|���{}�g��rY2�eCW��w���;;h	@IJT4;[����g��Dq:@��C�,�.ϴ^�:��̿4�F^��<����lJ[đ��xcu�ڸ���}�z䰑C��8#K�����f���x�����I?-S[�:	p�Q8e(F�l6��|���[CNX��gIZL"6UFpp�@@�Րﵛ���*f{�! nG9No��+ g�?vK��h�����*�t�v<��qƦ!@Qh�⎣�����8�o��<���,UT��8�n��t����6�(���BF�0�o4�H�X�'��~^��ͽ�6-�e?;*H�K�)w�]�u��z�����[�[�97]yƉ�8�)�B�"y��<�!�a�H1��
�7�Mͨ7�)r(DUb�;��|`�hM%�B�FF�%	e+�:���$�6��3E"����&�������*U�	3��,	AQ8Ko&.-}?���� �Π���E�g�M,O/�ΠR���3�>���omoc�O����֎�xT��3��jMw��P��G]�=���!�'�� \��2#��'I�bg���n��j���/�P�u��.����(:t)H�>�V;&P�ҿf��cy�k���Q��pt�����"P�H ��'P�RK�l�}�<xY�,7�y�O�c|�g�Y�`��N�����:�g��L
��	4����U�E�&S�4��r���Bn�Q�C&G���� 5���p���`≽���$�|��9J
���{5�~K֐��i�25`�>9��Vk����?$��XH�E	��������r���������<����ii(�Gl��jJ���s�Q�p��M�kuzy��|�'c�N�!�қ$�bsܑ��j	V��gs���Usگ���>xꤊ4��$۶h�Â>f��G���ʚ@~����@�z�b
����������G��?r�|�S���e_�4)D����H\\��Ͱ7�~�xl���5`})���"n��q�5�߳p�qO>�oaq��S�!�'�^�)^�7̃�x��T�N��(e%��+K�Q���	���9��������������;/b,���d!&2gV��L>%�����20�2
�B}��bf����\r]��jbt�g�@ef^��ʵ]���Ʋ!v���w���yW����Xxዠ����rí��Z��f�lm��M���q��4���;����L~Ǜ6\ODe���3-��4�k�Q�n�- �/�$@y�P½;�����\z�Q�H��9�K߹�W޺���kk�X�/ʇDAs�MC# (�4gZ �8:A�̈Q:�>�Ss$��5�&(�������={�������T�������F�dEW�Dq���"�?�s�Y~������a���pk$�?&�<�A�t2��=�fuı�,�c�,�3[D�����1���L���ɿc����r�Kq�W��	�n�{�s�{="k�D��&��Mܺ>6CYt���!	Cԛ�d$X����pZ�W�� ��{����>7���n��lO�י<z��5;�,�Q@��_N�U&������3n,jjA$u��%g��/��4�� ����΂%���1Xa���FQ���<|K��L:��[O3��!{����q��TQ5��lM"�T;������l�U_�ε��7�̔�L�Ʉr���ϑ��*F�lx�9n��D�O�>�A=u�z�K��<��~�Y���+_�Jsӈ?r;r�^�-L�H�����*�?��.
rS/���ͮ8��E�+�km���T'<W��jA.ű���x$1����Y��[�+�<>[��W
�(
 �:}3)�S� ��OO߫=� �&y<=j�7�?��Jf�J��s0�{4��([~zm	�c��eٹe$J��m�$. �bf��
�-?��e$�u��� )�P��=%��8�Q�!�x¡�+��2j��ZT�O{�f���S��^�^��rL��Y���\w���[��f��dLm�f�̞H����7��̪$�7ځݻ�'�j�K/q��9��S�=���Y<��������ɳ���n��n���WS�ę�8s�����q0�[���5"7���5�hٜ�w��뭡 �ˍ!�*K`_�k���u���O�1;&?��"��w�>�I;s���n����ޜS/=��s3u�y	K�x
�Y�a�v���� "�M���b���xړ؀uk�g�t� ?Ж�hc��A��u%�/���F�6���o�- ����%,�B'��!�}���N��Yj�����+�9��������?���2�m^��AŅKZ��D��F�}�T�D�t\>�j[�lvS���9�l����RjP5�(,̣��#��y���F�&�M��n��;r �Ͼ #��8�ƛ�p���O<�Y�=F�#��|<�ѫ��#c<5;�e[a�P�Dw]T��(Z�q�wC�;�޽�A� ����HT-̏j�)��D�T�l��	P������e��.kEL�js��W_��W^�!J�i�9���^W3=��� ���<F�l��j�icCI���8G�� ɽ�]��Y^�h�ШT�o55����ѧ�ِe�@"�!z�Ի�3�R!�3/��H�;�*���
 Y"doW�%�+�����G�!��l�O	���H�}0�U���)�uu}YN��ffr�LM	��#7�!�7Y��M��0�n"a#����f��q���]�VC�3�{
+�+x���۲��%�6�Z�
33|��F愥ʌ�'��p��z�fb0������;�;C̀�y� �~s$���ٜ�3W�F�uK���P�nGT'��Y��H�S�uZ����P�«UM(US��!�%R��'pJ�,�Mk���ur2�K���[����zY�%ג�x�[w65�8P�	�����TL� #iG�����p��`��k��  ��IDAT4��]�)fK��r3:��y @����[)$���u��?�0>��/c��Gw����̋���l^3u� �/>�<�y�}c��vG��X��&]�Ғ���C�'�]�M?�RrV����ё{H�יm�x��q���l!֨`]��W�����T��7�����^2�G&J����G����}+�@�˴�$X~gٝ�UB���Յ��>~V#�>5���r�k���ׯ�fi!��#f���-
H��n �o
����Y*!#�(ϡ��Q��CU۽�}�(.��6��a�xP�{����&D1�a�������9+�4b���;���P���|�=qGp�K�}�L��*ΰ�=�$ϵzu��}<�X�VG����j��j7�XzosuO9�H2���E��ʟ�)��<����M�0
��I<��^}kO���H�t�i[Sz�ú*����mm١����i|륛��oܓ��a<���r.=O���/��i����F$I���"F\��F�X�`,v~ZlҬ�v���#�6�Ё���-�t����5i:�yfG���c(FF"�B~�g/bn����.��|���㨚D�{ ?���U��Nʿ����"r���{���L���bl��D�\��6��)�䟟E�YFyfo_k�Ǝ|O��-��e=�,�����H3�0EO/8��cM�XV�(p5�ʍ_���|��x�#�T��W��� ʫ��}3�^Ba9���^������[��̗d��qO�+�����$d�{�2S$�f}%u�޺轄@�M�J���s��g�oL��}L�a.JsqP�Y[{�p�]5r*^>b/ML��X�V��~�'ϧ�ŕ)�����J�-|�[�7^�ą�Kx�����Õ,Z�O'�`���A_6;��ӱ���IF޺�/6���V�b���Rр��؃U������t:ء���e��3�n�w���y"��R,�j�Y�c|%vu��MN�L?[�\F��x8E���T�
�w�X��9�~>�`*/�% bvnA�������s+�٘M���2��C�AZ��&��+�x(���������wU��3?��D�/�h?��w�q��)`��*�F�,Ş�i�d5�5�gu�1�}A&����]aϙo�0�`�nE�L����"��B�8x���X���e�<���X�_­+W����3CP�N�Ҭ��D�j
��0ό%TFŜX���cO�Oɿ3֖�rs�<��l{kGKy9��O��:<��,#Au���RnO��^���9��ӌ4[0� hfʑ���AN�y��
��x��	�������@╂N��8In���` �bL��@��w�/���3O���T�%9J��˯IP�`\���`��yL��"���єg��K�EA΂-g )����%�Sq|ogW�J�,r�HP�K�<k�s/�&���a9r�6w��̡�h����a��k�[	�y�w�FoT3$|��8�A�=�lʗFB��X�������X�̲��mD�	R�ĸv�ܾ쳴�{�k;���`V(���.#����p�x�}d����<��5dWF.�|v��U4�} �yGI�A��8����]����ˊ��W��w���+�qPL̢>fV8iڥNj(b
]�#�N�R:��;B��/�b�*�� ��
� �"�@�R�kƲN���ؼ/��P{�)i�>���8V�%h���1ܩ!v���\Km�H��\�qKLI_��-�	�d����r�$�|x���m
��^��s%��:�A�<s������������|������V�/~zS�9�S|V\��s�I�$˴��<��O�_��O������&P�1n!!g�9s��(&{J��ʿ]{���A�Da+�)��G���	�N9n���3�W�XY]���gVHh)��?�(G-���?�W���~�sJ�҃�$�e(L�@sr[�@�>f�b��U��������/~;�-�_��'8����/cX�Ӟj�RZ�\g䤢1bi�)Yr���|_�RN�&(:-����Y���o���X��4��h��"���t<1����܅-�j�4�}"1ގ_��p"2���Rv(���@4�d�v���r�G�b�e퉒��r�5Bp�)x�lf؎���8�Yi�f;e�7����̼���5F������ù��x��s�x���N|\R��P�	$se� ѯ��m�qpw;�w�:0P�v���Q[���1�ƨwZ�_���gOdN]B��t��d� X�1`n�ƺ�R�s3#陹
ϐ�:fW����o4��� �2G�)�'(�DG(KHNŌ�|�|rIx���c�t3,����'�`��e��佗W����A�@�V�r�g8�y�*�|p]�h�_��/�~�>��ݝ
X�,��Zc�&��L��������S3w������VQ�<0�f7T_�8Q��<ѥ�U�-jM8�<zl_���p /?=]��_Bi~��^{�ܼ�����LJ3w��ᚖ�y$Τ�zG�nOl]�%l��7�i��J]�`	�:������<�S
�ID�j�<����g��yZ�z?QV���D%{�F����+��1��4�JֳCC�A,�\��d��_��آ�[70P�����ذ�=S�۷�އW�癢N��W1/��`/��JӸ$�s�2��m|p��J��r�N"�g���
୾�:�-L�ō˸X�ƒ ��{�7O���1��/lC���(��dz�2m�&���}�٦�e~�6ƖP�$�.+?H��	Hbf-j�D�f��6#_�4G��U���	�^��"�P�irF�+�/�9)+6���Ϋ@s�L��Iz=tvo�Ք�n�����A�[5��m��I�!�9���-Ӵb��|#�e�r���Y#ٶc�m����t�R^Sl}A����A���Է�k�ߠ��M' �u�6f��8�YA�4���Q�u1��"���x�F��P־]�{>_~��}<@1GNJ�sH$e5���H&S�5�J2sKȹ�+����������N��>�ه��?�JSq��J~I���Xo��Ǜ��4�t��V��O�rT���$�'&-9����yt�rw�|\۬adeOl�cS����9)����9�+� >J+!j<�⅋<�>����<4���^1l����?���&a����:�����iIc�����z�$�W�����o��5�Sx��%ܼ����o �y^��"����GM�1NΒe�3�S�c�����]23��̖dh�-#��c�Qm��é�����xo� q1�g/>O�+���Hs�����{W��q��gQoUq#1FQ"���b<��-��503盜xx�&c�S�u��M�Om���$GDol[fzP0,�G=yJF�%��Ij7ᘲ�?��r�i1)�ॷ����a�L���e,��-�,��p5�+ �+Ghvq��}��&n��No���vo(kK�%��E�G��r8F�Ͱ6� ������c5�������t[��"9q���0-���ݫ,t*��:(� ��tn2|��f�Y��`x����R�Q�aLr�!2���������Q�{76����J�Y|�?�ܲ�EyA�Z8�����S�[M�S�R��TT�募��g�]���\�(-2��u���X�'�3�%���Č�1!�X
Vá���$��x2�T��#C�l{8%I�	倕uiv��Eitz��[���UU�ɑ�Z��X�wqV��z*�Z��k�&6���	�s��6�'�'���o�s�XL�<K�=7�d��,�4�j��}���M o@�!�v���=Wq���89C�%OKL�1�0��@��nv����}��Զq&�	�wRl�gl�B�"����Lb�#bb����쯖��E�����WL�wZ5��;�{eY��
Xk�<��K�n��h����3�m<��[��`  J�_�ev��I,�.��}���ؾ�������oK�*�E�JF$Pf0�R`�����'�C��YOk�YJ����W=P�!%�u|�uc?,���I+�յ��h�"
B@v�*�w�{1����0*KUv�mb�w�$g�ԁ�S$V�� jU'彝-���)ؖ�]�u)ȟJ�$LϬ����B*���DŃ O'�ý��� ��w�+{5�7�#A����]Wl�%�I����eŐ�H5m�l(M�QИK��M�2E��d-X_�`H�?7l�dpc�J�� ]��CY���Yi	����z���٘�ߡg#�z�d�<!�I���b��)x���z�+�_�����J��b���Z��1��L������4=L¡2bПг��ΰZ�$��u�xrN��§���~qU�Z���P{��2cm�,+)Je���PH7a��l5�x0H���k';B!YDr1%�1�6� *�y
x`N��u���t\F։x���F�+���[7�/g���!��f_\�t�loW��<��gg��ʠzT1r;���l;U%%�u4����M6��+��"=[��t�O��ڗT�r��yd~�k���xVս�[X��Ul{T,��~�?��ڑ>��蟽��q�Q.i|-:
+�O��n�<~!z���G,�1��OX� ����9���jLrJ�b�T��1��Q_'�JSi�;��+�~���O���R_���ca�AnJ�W�Rf-ұ2��c=������_G�h�F}�j�����ā�� �Y���z��-Au@�9�<IJ�"�#u'�����z������L��f��&r{bB�3�^gN�c��?F��<�C%J5D�Jdj������Z�����4aR 1{7�=d�\�vO�iK�������_���������=xu��2/����.�}�J�fM{��[���3v�ۏ:�$��u��d1��̽��3�~z�t��{��a��,R7QG`E��r=\-�C�|O@y2�גw{0֌\o O��E6�G������A��m��$p�[H��u%�"���IY4b�+0�|}��l	��{+O�����b�/.���Q�D'�m�f�SW@(3[���=u�!G#u���R�'�ľ�����#*�s�yf��@����	H�\#���eI��n�n+q�t��白��Sl`ՠӭJ)��=���7�/����������M�޼����|���_�Y4k���{�����1��X[��Ͻ( ����O_Ǧ��'�����C!�wP��^iSx�w1~��ű퐶*8Q���-$�;��rlȳ����t/��NH�m�ߢ�ғY:�~W���M9n5�=�4f�7�sճ���@@0y��I��������sHedm��@���d���3��
��X�3�왣}`�Y���yUHª��ʇ���H�l����b�_�G�'�jh��h��64=n��P)�Q�X��;D!� ��9���+e�\[z�K����>>J��ze/%�1b�<b�:���m1�E�e�&�-eV���7�"2���2gf[�����!~����[���Y<�\?�s�am�������ޯ)YF��G/>�+:k������ ��p쪤�R1�#I�,�_:�'�P��|� Ӆ�+f�����2��}iU!����Jz���=E�C|��yR1b�Q�c;b8�=9�+�SP����O��5�� ���g�<,^j��<�v|�O�6�nf�8DC��;�	�*�,��?���U$��w��N�)<��<�}j_�f���{�~����%I�CI�l�IܗHM@JSP@�`7p'�s��O������ѡ�+ؓ���%B:x�-��\,�0ة�T�A�S�J>Ym�0d���1�/�&N�h�U�,n�x<���a�!�lf`��3f$�&0�$�D��N�o�!�v���%$>.MYf<�Sh����D��^��^���(�a,�~'�z������%������y,��C�D�b��R}`�$�p3�|�6^���m��=Del�@�u��Ӡ��� V��<���B'����@�q٦3�C%�ㄾ5n�n�0S������k@4f��y�p/�'8�"�s���!��%��d@ݰ��?A�ꏵRC�Ggh�_n苣ꢹu���#|��2rO��]�s4�G�QεL9�g�YA�n���~6����Xݸ���2t>��Ӳ�������6;S&��M���<�<�r4S�T�	b������ �e8��$�-���PDi��
*):���<1�9P�i`�;k���7.%ͬp}#�Ǿc����Q/!�"��U)A���(�t��`���x)˦l���X$W�i����5}� B�@�Ӽ�����`6 ��__?ف���V_�=�\�6v��-y
S:I�Pg�f1�}TNZ[�Z��=(U����2�XV�#�>�`�����H�K�&�����Y���?�-�.f��_�Ͳ6Ů�rE3)�����&���8���?�ޠ�p~L?�p|P��M�)[5<��"b��.)a�b*���L_�ccw��S�V�_�b �Ӳ�b#S�� �Z�~g���Lu�;��i��
��[���,�EJ�6Ɲ�Y�SK���Y�'�C�{�n�*?�Rβ�$�2	ͨ��O:�p��=�ݖ�a�o��&,�AdՁ�$C��Ŵ��uM�V¸�t"���O�3n�zHfdf�ŋ�g0���ƺ�uR�7 WmG"f(|�����X{w$�/{B<�Ø�e.^ZA���yRL����}Y��-	^���yd���\���@��=lj�W�l����+�g%C���i?b��-����*G�\��t�I��ı8#F���I�*'�뒍C�!#]wb���]�X���c�4���?�`��ӈ�$x�*�7�B*1��8��!�$��G����W�Ci�����b�$��$"��8����L��M9e�y�r�$bi��b��)C�lD���G�)g+7�h�R��T*+��}C}pzl?a�7���?.�>(�Ћz������j�i`������o�7����H�8��#fޚ^}���r�dS��)O��1>%��Tb��s���^.�
N|::)��@,�6�`�}b1y&��=T�ql]�P��%�V�Ab�|#�氁��E���*�x��d�34�u�gjb�)0�ޥ\<�����I�	{�?:e�_�Y�(Åc^(�(�e�V�dako�@�K�%ljw��a.\@>?��|��>��cX��L��)���ҥ��Mw?Pb�w�qTo��pH�5����sY�Lt��41&1y���q��k�p�O|ߔ�<u���ò�?�cBmLa�or�,�`ʖ&cc�da��$Ses�u�h�~��vFiT#�&��}�@E"�8j:��\:#�o���߿������c��W_Dr�����v[���t�å�`�'���^k�8ع��1�0I
f��l�|Q�L]R��1�x�f��ۉ>-OHê�L�1�A8I�r�����\#g��%l7O�Į4ٝ�?OlF`���8Mb����-
є�?�@?]�d[���'��`"3�L��$���:X�WӶ�f��^��i+�N�fP�	ꋛi���\YQY�h��D�8f�yH�h{d2�$V-X|G�������_�*.]:#��
/�4噛	�
~���W7w�s�
̺�X�i���u~�W�v�7�X'�=�r��t(����]'��6�8'lڢ=9>J��H<+�e�m0��tǧ���lf����"���]�����g���/i%�4�ВfL��'��L:}ɭ8RBwG�ݹ�C�s<��dϗ�8�M�
��y�$���U��s��a�D�)�lQޏ���1JF�)�3��R$�r�3�d��#/%`q( 3P*�b���^��k���{�(��[Etj�2��r���q=3Ĭ����E6���=¾ن��p ��Ґ~uЌ��|/Iʢ��	���կ|���7���\��6�z[l��W�-���<yQ|P�C9��l�����O㊞���,ٳ`��+�g�r�;F�ёu;;����U<�6'�>��76�'f��1�u�������P��ͪ?���Y�$�F�㴙Yb���;6�V��iw�uq �pve��t���#�@|b�F�~q�}���!�M����F�< ,ܽ��;�����]�hL��u��?�����z�Uu>���l�.�d%Kr`S�N#i�D1^�F��a�*̨�r�'���Ѡr2��
-��s*�5�H��(������e9 Lf��W�@Z+f��8q��`6E�=y߮ ��|�IYUU��Y�~Q�c��?�P�8��H�&d�l�QK�N����52�Ѥ\:C*�$O	�'tBT@�����5��]��N���ǓO���3�H�Gʕ�2�2b��z�~�����q��CU�b��o��H[��fIlJ#���t�$�i�O�H�ňX�0�ó@�Bk��HϏNF�_�c�F$�͝�c�v�2���3��Fw20��8#���h���)��df�
�?+�%AÉ�=q,qJ @������\�u_�)�Ý
��5��*U�x�k�B���w�`�2�/��K��Ň׶�2)��+eKm����6�BgR�����vZ]L��&2z���l�]tN@��}?2����8��;iT'�+'3��#��@�����Wt��1m*;8Yn1\�VP,u�Z��B��WT��km��A^�	�ctG S��'��	I��3�`ϛ
��B~ðWV��f�öL��B~�qjqJxD�dW{��9��}����a��ʍŹ88a)	*k�!^{�}����!%�?[ȫf��4c~�l�-�q���l
��B=d�#Z�8���s�죣ITG�ޘ���KV%�b{�r���oE|�A8�k���Edr������_���I�4�{���Z��j��G��ٽ���xb�A��4�� ��#�#�$�h H�aF�x<��'W̊����Q;�#z��,-R��{�EVU�ͬ>�ȱ���ʌ���ܟ�?~I��7���."�[6�]*d����c���%��5�1�	 ��{Fg��B��G�7U&KMZ���J�J	�=���y�R>�!��}�O����xi{���Ex�'�k�ve5cz���t�=����mL#7N ɬ����]�J�7�'���Ns���Kyk&�Up��u����9=|���q���Q�c%�S	��>Nx���)<vi[���k�\k	RK@�k�fm� ��u�1�~f��p���b'���[���k!��5ܹ��sO���B����m��O9������8@���T	��	ʒQ�"�s��=?�W�(���^;�b1�b����N��M7�}���{���/o�
����R)�\��ze����oZQS�ip�a���$m׵%Ǣq8�]nN��P�b�?o��T3�Jn�/?T���	�$�z&�+�1��1�H�h�~x��6�����@��+ύ7���3�蘆1__�wF��}sU4����7��k�,@�Vd�N���F�%S���@2"��[���G��2�"< �*ӻ��ibF�I��AZ`��7��x<Tm��$��F���}P5�^� ��5�l0[�����90���i�ܺ��&�Y�>c�8����|ˤ�#�,K��0"�!�F��^z���⅟y���Ő���]�H���_�g��?����z���ܫc����"�l�Q�(��]~Y��w
ὑ�H�)b�0�x�4ED^w�N$�\N��@��F`���L#N?�4�,�/P�2�������ω�fJZ��oW*p��Y��(@�N��{C0�n�tl���d$�,�?4�
�#�Wrj� Ŧ*�C����E��������N�#�|Ĉ��⥓�+� ��`k��e:����{Q�%-�Z��G���xs�.�w�9�������Q�?���%�ß=xv�#��,�G��'��;zm�kH�N7�:����X ��G3��]N�����,f���i#K�4t��'�*�ƪ	�d����"$�lZ&)��{�
�e��]x�"��Y���m����(�q��/k�D�h�3���~�^�-. izx?�!�Dԟ����GT�L��:@�����?���im�L���Y�Q��M���)�I4�{H���`"��+�~G�J=k��W1)�4V��m��(�#��x��FB�b�Ȑ�;Ɣ��M���E���=�%�$�L��8����A�v?����S]ծa$���nEd	B�p���s:�Xi=���ʳ������/w�qI%_�Ō%+õ�%u��#��8��`!G�_�2hp����`/q˥)�W1^�cT�weo�O���/�0J��;=���8fh+ܽ�f�&6��g�\��[��(f�����'^���p��,^{����h6�����g�AU��������Zpv�q�����ټ(>�ӛ�}�������i��r�K
����7_E�_�/��y\���[�����h�y�+�T���H�;�tdϝ;��k��+�Q��6�1,(��1	l	�*aP+�l�����1z�&o O"������'yF�qZ��}�A���~�k�ڷ�ce1�M���cߕE:<|���� t���5�P���tl��	���cG<��p��_$��4l���do�ಧ��7�dNbl���|������
R���Ξ������I��G�2\zz���
cJ�y�s�0�č�Ӳ�e�f9������(�"�J�3��L���%�^:��1܆��S�<��m�/����v��/�����	��K��n�_|�'����q��W���}��N^_��.�E�"�e/ӫ�<�D>�[	�K[-2�Ʊ+�eFY)FXC1��8�x]F.��U~I��H�S�w���:p��@�:x�H��37,]Je�L�F���A��ۤ����F��INQ�(�H��s���C�,�v!�n)  �j����e��?���o	ٳ��C������g���V��m�˛R�0��r/���Tݟ�Eܹ~m�L�}uٓ�#
m�8�!�I�D�A�z�f�JM3q��f�~��a��cV�|�hϚ�f��Q�W(��g��j<JR>�����8����\�S4�2΀�,�8De���d�J5�7g�,RJv|�4%����ƶ)۔��96�W��u傔��̀"��?;#�+P)q�6�OPr��s�����q��i��<���`]Y�Y�?��w?��[�����Ǡ$_h`g��m�2%����M�@u��������e�bU4�'c�E�>�@<C
����؉!�f�:�+P���:��g��X�#�f����r�,��/�o�����>�u��n���O!���y���ɝ���y�@%rm
�]�)W�P;���J݈�� �"���Hww��ݼF[��L��2E֦���+ǵ���7�}�8�^X�3(�1͔d��M�" _ȕm�|�/����?T���Hso;Dܻ��~����7��M�_<��w�h��	lm���h�/|�~�����Byպ���{X\���������?��œx�ګX��lb��1����Գ��5`�V��L�Ђ�����0.���������yO������1l��3�*U	k&I+x?j��Sy��̶�0e����ㇱ?�"�L���J�(���l`��$���/��X��d����ܾ��t�2��߸�!��cKx���X\�ps��z��EM�u�*��c��ju�jy����;���T뜥�
����'���1���B�8�4��$x�����O�?�iOܿ[��<���+f��F������/��0�lg��\ O��T���A�F�U477����ʯ4�*��r�@��iC3����L�@���y����b's8�K�S�W֍=�q�41��%n�wJ�s)�_������L�R�!u��9��XB�E� tR�iV"9���md}�FR��<�6�-�]��N�#�zؓ��)��ltg`����>V�Ν��^��|A��������7��.:�Dt3������ua�����E�Y�Z���K�7���;�L�e���`s���bd��ڵ9�� -3ىǃI�J���H�^ M�ƺhӌ�H�8��:E��2Z#nr��l�Jػ��e!J�9"/�B��5Ǯ�^5�U
�j�G4�����9¿�7��1~���,�O���D+����<�����m�`����\AR����E��U�2������3�3�����T�u���r�>.����\��2������Gȣ���3����2�q��s��?9|�4�8���l��n�C���3�) =c�+!Jyy�6�t�i[&��k^���"G���#�h%�R��ϸ4�u����4i�Kt��������I�Jn��j�\�`Rk��{��F��ik���6���/���q����O5�"�t
�h�hO�C�*���
7�$�T�6�G�GMX\�{q,;h#�"�:R\=t�AA�o���f3�k�{����k3~���SJ%T�n���n����rs+�ј#����x"o�<�	R�.2`>F�9GG�ʵu��4]��`\n��$��7��륙o�ċg*y��@�ߐv��yXD���&�5�25�1�������Zc
[_�2B֍�-��r
�o�·.{x�~�'��޵��J����5�}��}���]�;w���)���sϜpw�6���j�/�{zs(4J����^�~;B��Ʊe�j��z�w)�q�Q���H_�������窸xaww�;�h����CϺ���}��l��r2ӗ�I.?������ɟq|T�ej�T>l�l��G;���ƭ�{����%�ʕ��U��ߴ��hԢ�X�W�e�r	K���Pʝ'�8m�Q��卙8����"I)�]��V���8���_��+o�c�B�O}��Y������(�e���?�l�:,r��W_�;�n2+"`d�\�PR긍mv�i�UJU�6���Ť��J�����:	�i�4�U�;U�,�y�7�'���7�c�X4��8y�q�Ly�G8���?��c�a��1�
5 �q#�f刬���4�3����&g'b���C	��.��N���v*���ps<7o3�L�.�EG3�,k�v�xVJ���Y�Z3T��De��HȡsНNφ�_8��z�u��pp��w޿����{���x��όyM##���ı�2�涤��A;�d�2�Û�%�D骙nլ���r'WSw�"����)���efԵ��MȘ7`$95�-�~�M@_��O���%�F����ԺQ�m����������o6i/�R�e���� ˼ݓ�����G�Z4#��>��������͖�rd�#��df�w'bm���3�xCy�37;1f�~<������>���{?��Y6`�)��ل�#;�;�$m&H��X�:������O�e!מ�z&��׭F���M��b����x:��?)�	~��jB����\��J�6�Ɲ���J�S��j�=�3����&6w}4w7�k� {C�ʹ�5?���N�������6�Q�l��b�v~�Z�9�/��>?���.m�vFv+�
\	�(.hJ����)��u�f������΍i�ld���X:����F!��b:Pt���0ݿ��N�q{ ��P�#�:��?o�=4���ݱ*@��*�#�?���j��#�ƻ
���8���S�/`�Wy�n̥	���n�@ �GN�e�<��3�T�:k�2�UcǞF��H�\7�O��g+Tfm_eS*���ަ��+�	��U�/�D=��,͍��D�.�����÷��2NWC<���T��v��/}��~�;tF��+Q�Z�6���QoDL�EN�0�gL�����6��<�bD@<�O���M0��5�h{�.�M�vE� �Q���򼝋�,����O�K�������u��#g3�ٟ�i����c2N61��y��v6Ls0�����N���>�Y�g�by!�� ��nגp�N�Xq��r�Q̝�4��hp�v�ȇofM�v2�ȭ"A�I��nގ�տ��?��nmCgZA���+�_ũC����������,�oo��o�����ߺr��w�o�Z�l�U�y��к�Ƒ#��ɉ����x8��?A�F��_�Lf@���17��b����
��!�e�܁8pñi��pN�=�~9M.f �f�h�i���!uY�Pq�O3X�Л��bK�ds�Z�:���hܖ+U�R���E���wna��`�u\&N�'栎'��qR������8���<������n���{�o���7�'�u�����t9����9�x��N�.J3cG'r��;��xq|H�t��iƋL��]ql������t]Ӓ��Sw.Bq>�1�KV&������!/%�k���8�4b)����U�&�Ne`��8��R�)LQd�l���Ue����d@Þŕ;���ª������|��	���>�n����67k% �5�)�Į�x�U,Lj(I��S�l����Z2]���g�Q2F��ɨ%iǮ�J�n��>:�u!9 �q��~�E�f»"9��r���6z`��a�"'�]��g��۷�_���Mc7ZK�75Xd�&	3��쎂���5���aZ�\�R>p�L!;�NX�Dف��B�C��!�l�=����������;�[i�1q�Ⱥ�}�4[%�EIc�8�O�ʯb��~��ް�եEk��M�F�G��}���.^<�g�y5��=�4���L�L�Sk��qp_���Z�����p�f��͆���\�A�K�k$�H���x`k���ch��Rz1���]EVɥMq`��jv�.�����kl��p�=
MJ�p�Q��#�8�pn�.��&���ɝ�;)�P<v	^���RI�:,r�N�x��"���8?Oߐ����n�;�P�$j���{���<�|�~�{��`\8O�H؂k�p�����7#=��U*䫒!J�Ϣ��^g��Ɨ�k����?}�\:���+�YC�9<��Ӹ��U�l��5=��gţ�:ڹ�x����7x_��{�Q�6��j�O	:-M	P�� ��U���oL��h=�h����ۘ��\��]���� vF�qt��́-�����DN��(���ʵ?��hcg�8{�Q��_��	29����1EXg������Ѩ0l�_��"޺|�������?�~�W���K���c��z��c�un+��g �h�4��-�q����Ř�Q�C�揝�����f	��=Ɵ}�&^}k�a��C�|5��6�W_�*���ĉ��7�����>��񣣮��=L�!n�Z��y�����d����|��~�:�q{}�������X����f"=+5��kss/,̙���&׳;�b����
�"�O<޸���t�6�-L�!��J&^���*�5Lw��Г��C%W�ٮ���S.հSf��,N�C�����,Ҝ������*�hR��T���urI:�Ï��(Z�.���[���؉4�%X���$ur���(#��x��T��ˠ;�[g�u(�yFC�8���\17}���N;���}|�;����"g(����ƻ�����
��YJ����5��x�u���J2�D�S�8�QIK�)&5E�z�
�^+��,�V-X����U�y6U�M�'j����JhT��f�䐜dK���&��!�j�й�5��P簷?Dkw�H�����(H�͛��&��ƮM⬁(���2>���q��X�n4��+`zmK�]Ó��@�kڸ&?�Ջ	�>Do��[�]���W�-��gP��G�?��qJ�G&Y�\eid�<G"�
��tn'��.�^�V�)s;Q_�1�=u"���K�D�MR��/~���ײ�����Q9��?���I� �I�d�;����'N�u8t���L�ֈ��Ǿ%Ӌ����7�BG�7qݦjj[�L�n2���\f��IF�)# ��j+��C>_��Q��\��cp�2�2�5:�n�v��&�-Yv�k�����~TŉK���a���i��n���^���m:���:>����z�x��u���O�C1��@P���-˴�"tN��\�B�n�z�Y��[�z�{�� �"�VS����ĝ]iQNW�IB�������>U��.���&���M���k����c���i�|p����e� ��`�[y�bWc�u�+�Us7I"� @������1���;�9k�����	4���-X5w�j+ܻ-���uo��)��Cl�� �G?�`��}�O�Cp�{�q�ω綷u`;>���fw�.?Ki�1��uiK�l������'����V�2�nH�㒏l�p�{V�#�̿9�I���/����-��6^��e�W���o��%��]��(q���3��W_�{]���~��m��K�_�Z�&
~���l����1�c�����kzX\��X��C�D.ӯ`�O:���<m� aA�bi���{����;���[6�����I���A-�oV��F	��8���}�^7�ПنOB壿�R����5¦����HĈg�$����| ���U�ɠj��iɛڰ�q_�\�wo���yw�>���GjzM~���׫����e%�Y�/�P����w��/�V?�#�ǽ��;�o���=��16�+�M��As�����>�|_}�U,��/�X)��x��'>�<�V|�����z����G�c�H��� z)�KQ���_������E���o�G:q��t�L�bh<F͎��h7[��|e㺻X�6�Izǟ�q�kV��q�����	ժ�^���u��:� ������2�e��0�7N�J����T���s�qg|���7��ǬX�5ld�`ԁ��Kly����e�f�1ﰴ�&Qfl��fB>�@�f����'��4��lӆEp��v#���:�n,�q?Jkb������M�[�5k�`zj.��cˬY�4��$�d\֭A��Ae����-4Wʛ�B���Y��,y6r�eh�rY�P�#���O	��s�ȁ<��~Ɵ�S�����C]�4R*�M�o�ߞ��G����(Ka�?A�{k�7�cL���'"�{�mP�pQw��b#�B�c:���}o�q�}�$j�Ҟ�'N��#����m5b�K��%�+�j�������y����ќG��F2�٭L��
X,������]7�L�����(�m[�l,qeG�wZt�tf���td�Ne}m�	o�eٲ�9~��J���`h��	���[X���&��7x� NA�(TC��$�TJ��LN��abSQ$�k�n�}et��% ��*��h�W��q��a>��A�;GF$K�����E�ʬ�	T<���Ex��@�c�&��$��|���*��иX����kZ��a&�F��^:�A�n`Sv��_����ַ�[h��-%V�X7��_k�i ��Z����ĸO��:._ż@o䲗������Y�|��g�{]3Gd��kp��p�<ː�v�� v��x&�%�Y�L��8�;��Ա_=�����M�p�)WҳD��{0WZB�4m��G\������B;���-�P�,#���a�>jL�$U,���x�~���@� Q��"A��n��X���C΀ڨC�X�t.`0�t����x��nq:QHt��;��/���h�f�R�%�"
>׫�t�s��Z�:~�+��ל��G+��&Phז>�{�w��n���.��_]ƭ�'.<��F��:Z͛���/�g��L�܍���%��P�uH;/�ĩql��UJ@{]�l�Z��àͳ�B��j?w�����J��q>]�� J�R�৐�����"*�w�B��DYf�h����� ��vi����}�����g)Q���Vg��߼���7nmXҢ�&��9�ȳ9Ζ�W���P�v��)߻KD���׮���1�x'��D�%:�B5x���;����:<�_~gΟ�/<�j����g��4�{ d̜�	�f��k�'xL�.����7~vPf(D��*�x����/�_��?FOB�
��9l�JR�;0*�.�7L3l��-���pJʚu1�J��N��ƕEh��Ӟ���Fy-�a�V�;�7�&�y�Q6c��B�,W��8mnRI㮒?S<���	�\Y�Y�Hс��"b.��b7�c^�Ojw���nj��N�C����\m��K:(�Q�V��$�F�<8�X|��ޔP/�GGT�f�;>�k7����;����R뷎[^�#���X�R%cz�LB��q%SM	XW&���Z��;-#�<=G� ?�E�XF%d�ZʠJQȋ4��Z�S)�+��]IQ]}��뇎 �N�N����l�Lǟw|ES|p��%��o%��t���iz�9%��84�0�2R����]�1:S}�9�!�0� ��� �3����>A_�D����h��(1�o�x�r�%څ/�����3˨���i�S��Ͻ��Y��w��Y�&nd��|&㜨�^��� ������J�8+7��K�{��9<����]�t�y~�*F��:1c���t�.�N��i61�!�SΆX,�P�X�7С��t>����3�0�q*�P)W��N�]������0X�@�ֳ�˳;Ip��3!�	����� ����g����+�k�-*$�'c'�|����5��1�-
e;Q3�We�� Z�F��l6��@�QGW嶮�g߲E�:�tm�C�q}�8���ߣ�]��;��k~�$ZRjM�IqC^�������:�}�Pt�%�a�H��j�ے#!xW�]�R���:ړ��!�k��m�_ƚ"f�m�5�	�gR�@�w5`��y/�pN��e ��y��;���-���	C�r��e+�x�4�����)=�&���?�&��\YT���5�����x6��m��B{�B<4���8�Yk�*I@Z�[2c;GS7mN��K���jV���:f���H����S7A%:Ж�L�#1�n��@F+v��4MJ$�	��NYAA�i*�~�y�ƴ]��Y̦�/�<�y�g]|/x�������k��m��r�v���3�f�˸�~_zu�8`�r��4�p�i�X��z�~�|ي�k�������Ҝ��F����#z���f���d�����!����y�5>���]\u	O���(���y|ķ}��Ѭ�7 �"�x���x��:�K�^�J�	2��C@�{�Ƶ�|oQkUt#Lǫ��"�w�*�3�����f�gv�ӧq��I'-�q���j���D�=���.�x��w�m��ewXbľ���q�k&�vjh���u-�q��M|�7qie��
�mm�	��������iQj��� o�=�qV?���^�M��+o�����mm�V�[J�2�@s�1)g*rQ�T��Bo�e]Z�T�b���1� ֕���en�I���?@_rt�9�)#��{�xo��cG.X��!����`r�H&O#�\�wX2���왢�5<h҉����xD��C'�Ó�(3
�nmX�A���x4"�FN���f3�q���:�{�F>�����Cag�]��{F���j�,��j�q�tt�0�;{����d^$������AJA�#}�ƈa��?�4�B>a�R`�*�FCH'_'��<FC*Es���7��'`S�G;e`�y����)�[tVHS�* (귖0�^b��蹁�#E�ڍ�e$>ߌ��K� P�-�5�hd@����2����4�{9��-��`�#�([< h�����ή������V�kbsOeQ.�H �h2=�So~����Tp�X͜z9�1_5�{w۸�����}�3��&�����Z�Q
y�!h��s���o�����[���EF���*�汿�os������"ϔ�T �pE�j�� k�&��t��cx��Mˈ��t���r%9n.���2F<c�n�J7#0J��{�!ww���E̕�H$Sf 67O��C�=���*�qg�aeނ�rوұ2,�[���'���%�0��9� [VQϑvX�g:v�Z]�ɭab�Sexd��Ә��
����(�������j��V	^�ʂHwjL �-Jr���<k��1}�� 5~N�l�� ��T`01�\mJ��� 4X�j

D�=��=��k�b=7E]����*cP:�ԙ�vg6��OǷ��N�>f0�i?�yC2?�<J̴�f��뚞G�ິ��*ǽ���»�C��u\
��iTb�*:��~�M��X62g�4�t���ؽz삮"�T��pz�'bF[_Z�2ϩ��i�	|F��u�ۏ��q�0?1�<剕}����5�n^|��#s�L$�4�̥7�g7�Pv/=G!*����+��s��Ou��S�q�$t�u�DeЀ�����NUU|Z��*�z� B@���]��A��x�Zi��|��R ���S�N;����Z��Υ�ghW&�n�^g��L���Tt�Mq0C8w|j�:�B�7��)���$�X����^H(X��~�H4;���m�n�����$��CR�~���	��,�GR�EC�����oަ���_��:�&rDO��՘X��РM^`P�f�=�b��GϞ����Pzi&oB�,>�W�����oр2r#zgzƁ���w�V��*\��m.��?e�C���[o���+�h����X9c�gEt�� 9��(>�Oд���%:�M.��h<�ڷ����ރ1�(<���,}��W�?���o}p�F��Ȍ]f&��{�4>H�F�AgB`��G�F�.�0�Y���&@$�@�����PdinNu���Y����%���Wgͭ� �q `��5Ö�J���A�B=�Of�c���>���Ʌ��%ǿ�n��B��}���g]�su�;i9 ��8̀�R���>�2ct@�u��O�۩i�=<-����.��xOI 9���/Y�D��cTߢ��ڧ�����oO��He_#q�&<-���\���0W������WkY���	=T��%�Ra%�B�br�l�J�ee�Dl&���"�B��(�2c���$Ӡٙ��'�3$���Lp���Q*К����k���{g�N����P�>7��'p����]G�G�	����O !��2� �`g���#�E\X�p{��7{XoG袇���x=�;c|pm�|r��������pju�`���`_�-T2��2/��+�g���X:��}'q�h�1�� P��O}�S&�ܾC[�' ؞~���P�[@�����ig�D��l�����M,,,�P��_�T��9qrU�nm�رe\�Z=L�]ԫ��94��f]�vm��e��E��]����=��:1���ԺLo�0�[�rS�y�l���3b���'(>6��d�a��>mRQs�5�vȳ�?��6f���P���m�:��5־Pf-r6V"�?��c��rύ��ޣ�E�,������
8�eK;L]�"�p�e�7�xS�l���$gM��sx�xd�te���&Ď��{�|�8r�K�EC��uFQ�l�$�{]�r�|��}P�"m��t/��C��٤>_�5Zؘ0k*�kɹT[VRB�Z���>��]m�Z=4װ2g��K�1�k�f,��xܳ
�::⁕���{�0�d�����&�����C
��5mJ���j�vm���2��uL ���O����������#<r�n~
򼴪�&u�	� �d=Fηi�d����-�w�y�c�$	���"����Y7(@MQ���k�j�>q�r6�xB����QV�~r�-���q��kx�y������"v��������S���\�m\8s��i���|�2v:M�gp(�A���;m�?��)д���4��p��S��=��!�:��2P 8ow���s�W.�s&5��r��A:�O�(������5��u�jv077�u)���O�}�t�������Z�m��{{��^z��7�"�)+��*�X�#t'�'��.퇤��xߏ/��>�lꑴX����<�gpf�X�����:�F��`�:7 7�f�uz��yd�Ay��<׉�il�ܼ�?��W�P_��|�qT�FYZ���l<�O����i�$�gY���ћu���~�w�?�����=��s��3�kb��9�����"@��x�eR �W�F$q��"=�T��v{Mt��|�g܂���X�qY���?�\&�ÜC�7B`A��f˜�����ڣ�Z��>�������i'�?u]�|�Id<�C��k [�_�`H�3���
>�rɕ���|]-�qڄ���-I�f�4#�!]3q�&���Jx�ݵ�59>�j�:��`�	��j8sr���%��k���>����V J"�X��c�C"���A-��-<�X���L#�Z	zTʓb�{飾DPH��hIx�5� �2o"y{ә��7g����Ӈ�w�f������y�qE��+����랓7U�|�{ݳ���j��s���t�B��-�NI��!ʍ	����K3�����EJ�e�hHzm�G�r���(��F��nn����'6�W����w�l5F-)���F�W�ps~�L�x�������P��4eB�o8Q��T�Jr��Ig:r������~�_��W��@}�k�U^�>Q�G�,`ps�g���}�H���dr�W�z�Uh����~��#��JX�<rO�{n���8���{$�:��掽��A�R{�#��>��Ƙ���<�$�Qn`�?��y�M@���G��A*v-���<?{NYi�w]S�k4G`\�9n��lz���^pU�S�e�l?H�����)�d�l��Q��
�Ǎ��D��)�V�m����6�c�2�@�8^"�k���bl��
@b�Y@K�{�$MpXU�I����ԉ�E]�����%j�ʹ����	�f�̑��JMv���JO*3�8R�4�`�=3�Za�7:��z^�:���C������Vi_��<��ak �o�x.|��h��e��'^���9�	�	����)���e��J�&���=��������+�'͟��g�����������ܰ�jH#g���
�d˧�,A�?0�}/�����Y���T.Z� v��W��8W)�=3;�3ĠO砢�	�e�Mw2ae��2��c�4�������T�ڹЌ�u	琜=��A_׺Ǡ�C4�ާغ�t�,���E\�ٰs�R��n`��qL��@�=��bh�Q�Yq�����*\�3��9�S�NJx���x�~�ÅS��)������Lh����+�U���V�U���9��m<��c6��:�M���ʷ��o��x4������Y��ԸO�k�g��2�>G��R����U���k|��P�9��K	�F���������-��"G������D�K��{{x��������m��8�%��ȫ\4�UFܿ�_�������DQ��}���GU�~����Q�>K�#mAO	�>2Fm ���ou���+����|��׬�S-�R�c�1$��,X�Ѱ̔�y����]�6w �	߷��(�(Uk�Qй&�����-.��*��{��4Vz]<�qaa	Ν�#�^"�(Yj{cc��K]������֎5*� �K�Z�ь�+�>�z��b�xP��7�᠃7i���&��>#����Q�@��7w�b��t�|_,��oI%��ެ�?0�����,���m�������8˨џ��gck\��`��w&��ch�$�x���\��h�ug��J����3|�
�e�������,2���Ěf��t`sC?.�O:�mx�l�˄$��i�։9guYjb�6~L ��/��N�k�E�~�mH��5��fC��@H9�F���}MPR�� �;i@�1�yEobA���E�s��-Wk��Lio�
ױ��`���\�{��}y���#i��7�Mq��}̝g���9ó�v�c��P" ��%�����%�in�8�q?�o��Y��7���������}�4�D�#A�Vsw�֍ =%���j]o&���G8u�� j���m�0�]�s�5�u������ 4[���,P31�� ���� M+�a�4Vv2`��)Щv��ؼ�^��v�f�5���+t��s{��"��g�yt��\s<�e�ƕR�JQ 7�`�n�N-�]�V�LBA�����i2�<0,Gh�Av���}��\{�� �ؾ����r��F_� ��!�X�Hvɛ5�+�9u��T�2��߄⯩�6m��x��SY-RN����c�+���#P&�6A�@3��i���Ƞ�hl��qb6%����g �&^�s.I�F����� �%П���������2����.^Z���v�`��b�����q��>LY�i��q�m,Y�Ny�er'i�����c.���&���dd�S����d���u��J��_���1������aέ�,;#��4-����/p_kzA��v��W��C��,k����C��¤h{��)%<k�=�0�������k�,�Be�յ?�1���>��oJ�ꌏ��:S�S� ��q��� ����Asg�'[-��#�ps����3\@#�`�&���Gk�C����A�� ox�D�U�TYڄ㹮�8$����M|��{{�����/,���e�䉟�oP����	2j���>���hN����s��A�,?����h}�\���y_z�M�7ֹ��/���8k_@U�F��S�[{?z��ޫ���~�N-/�#�6@�$����Z�P--��䥳��;e��'Opnu����<����K1����q��qfI%gr��Z��S%��1��_�7�K/\B5�s͏|tm0�TE��7]�A�3��G�?��p�Ɍ5DD�$Jd$�â{|�O�=-�H�~�&���Op��];q�?j�f�t���V	INE�C:�阀j�wm�Ҝ�"����NW"��MO�}F��Il���'�b�`�s�ʭ)WPh�c���Et��E�J����C�s�p"2����<z��e)
!�x�M�����l����}I*(1EP��]ZF��zgd\_�&��;�B��E]D�F/+��f���	�}�6��aҎ������?�
t�n�a�q\uKV+!�\�ݵ-*�Y5��n�/;n��	���!�u��{fx��N-�qz)o%��:�s��9T򦁪<�e��F��sj�f���)��s�;!:�UAѼfb2��xy�9�5��8��uq`A5 ��._t��̑��F��`k*�l��ȕ~�ne	=�.��w���N,�v���$�$�H����7WÂ�*a���ݱY�p�'Xh�c��6��븵a�8�~g�f'��b�Fz�ۡ�z=���n��py�6�lvg��}ϞĮK�Nx:���*�!�Ac�_"@S�I�؍$�d����ɲD�ӄ�$D�ߴ��� ��������[��qGqz���$��������P����s��,]��2�SebVUfդ��~�N k��#h,�,��a�ϟ灮�gE����b>/�5��>�^�2r��T�X�)ݹ��.��C��o�F2��#��X��ʶ��\Mq�
X<~
�l�n%/ce�	mN{���M�Z�qjcg�Mi���Á����S#p�s��r&��*�hD��nf������|�@&Nd���l���hr8���i�D���B�4�F�K%����,�wj>!���^�FOYul��(?6d����X�z���a�=�2��^Y!P�;�������)�}��Ľ�.6icK��.�`��OO�w]�ZJ[��y�Av�`����g>#M���y��@�+���$�ҷ� ��ٹ3�� W>Q�UA����'emn"_S=���8��f��o�\��mt{m�ӓV�<�O��pauqO�6Q9��)}ψ o�2Đ���B�eE�SՅ��lb��P�nb�!LԀ�����y��p�<����i��䌼&7��Z��>����95.e����*{��ǹw�Xk�������W���WG!����ʷ��c��,A^�Uwz��`��3��%=Q�����F���>�2�G����#�䥇�z4͛�	���/�ڍkV:�v��sfK�kƱ���yw��
����'Ѩ�e �0T�ì��C�wb��y�$�u4U���/m!V�'���GkX����jx��.����=?\�6-�>��L xm{���_���M��/�,Η}S���i4��s��~�i7S}��Ip ]g�i	i��@5I�Z'l(I�<�~�o�Ew3E�:ތ26\�-:�?��K�?����޽5�y+�H��W�A�h�B)ϟ5L_I������&Z��)t ��B�꺌i�[��A>?3#�QPDWD�adJFsa�h�����{�7�X�4�j%��(B���@㱻}׌@A|/b����?�1����IzW|�=5)������[u��57xI�m5����x��*��{�(�%:㝉8?%�x�
.���./aN\�A�^��S��|K;�=���XY�5��7��uGY߫�]�ܸ�csY<~�5St+����#��PC��UH4��w��쉳y<si�N.��=7?�V/�X�ӱ�,K	<��F4B�_�)a�]I�fĈ^���f����(!`��q%/Lz�^�9sesM/A�Au�6��I\o���i<Q�C�4���ƶ�U�S�JY.�:1�A���纹fT>V�E멎w��xyO���f�i0��k��"ِf����]ɣRn��XC�IPXj�A�ϰ�rq	��ֵ>���݋}\8����=��V�WDX��~O$y���plx�\ŀ����ة�Z(4��LN�X��X�J�����������Lo��2vC�&Q��p�u+�\�s�=U��(Nܘ��Zq�ƽR����%��st�C�M\]�(ʘ�{��O|Y�V�1�C:�>o��N}p'����^�<�UC�]H5��Z�މj�:amLY9�ci|Lgc5���O�I�P�L$���r%k�*5�NC0r�_Y:e��kCt���S�mn��%�X]d���~U�.��Q�qJր���6� ���ٲ�O.��YfC�@����u� �n$�c�:SW1Ps�2�H3|��ӈF�'�iY�Z]�N�M����[|�e����vy�'��&jpo�e���I��~iЌ��Z�S9.��3�T�m�b���55)�9��=��~<@@gZ��C0�L����yA|�>j�߾�l�����'h��Ni�ij���:79���^.ƕ����a�ת}>�UȄ��3倃���o�:����ތ2��|�vg�i7&<C���K(_�[�1�ˠ���wv�&�T�8�����)�#��w[֠Q�u��]C�*I`��\���/�͜K�?�x��9��F��M�=����o��ո);���s��,���˸qo��q�-qm�;����k�Ĺ�u����\A��e�Kx�_���_��o3Ή�[�IM��Z�7_�k<v��H��\[�K(��>H/k�2C�4�x�v��5���7���Q=�Q�z[y�U�\[�˖+�W�&���݌����f"Oy�Ifb�rq����U�n�Q�y��c���|�3��'�5�k�vw��4h��].Tp����\����W4�����"���ŅKS|�gqn�Qe�.��[�ۋmV���a"@%i��]���;���U����t�+X��a���hl��/B��a+s�,0KC��C���j׊��kȥ���#�>��9Ȭ�Rg�!Qw����������/�/���u�{߳!�ڄ>#�	7���4�&�j��O�=���|�=<�lݠ@��4|%?t㤬|��ٴ�B�y@�<�&�Kv�<�z�U�H�ڛ;��z"�s/2�xv���-�����T���j*��Pⲁ�H�O�h&����&�F�	^����2l�����}0$(��sn��uP�:7ZM݁���3Tor���_�.�����M��8iN�*����t�O*�0�7�0Ҕ\��.<e�*Mn�ƀI�:��VGع��W��Tg�W�ʢ��<������G�- ��3pD��/(��HL�Jr���ZFk�&t��#8�d�bF�C>7����$6ɛ���E�y�&>����o+�7�?U���`y'��m�H��z&��;S�\,.$�;5�b����>_1�\��s��@���}�81�V)f���U9��&��)/��Z���u����^���ׇ�zy�{��M��A��|�����U��ÚϹ��k�n({>v�A0�l�<�#�_�?�Q��e?���FѺng oj⡾������L�)��P���[���:�3h� ��Gr'Uy��*��L}�$U��(������L�0��LƼ_���d��Q�	�ե������a�׷�5��Ƞ�4�ҭTPG��I�/��4�t�����tԛ�P�O3Y&�ʳ�b�)�k�p�a�Qi� o�0O�V��4�m��d\�L�>��q����9r�2�#���8탴�ud�c��i������+��>K§�ky���g�:��F��qK���30�vtwo�Z������pWxn�8��g��[�]Ik�5>҂J2EڋU�ݓ��3jK��6�&���Kܺ�*C��5	)K(Z���y-��!3�F���#`����^�G8�N��>�|������:n��w$��yڣ.B��8N'�<�
�}�u~I�&�*v !v��wDS5�$�7���̥皮�S���K�+����q���%9O��(����۵�I�`�;�^�L�0��˳-m>/�-q�y�z� 㤡��N9i)�v��4g�N_:b��J�	V�W EO�
��s��wsm��{%�\]Bm.��0C{�5*�;o��+����ˠ7��P��x����1<e����+��Wqj��FY1?c\�tN���a&p�	U<|�-i9]R�o���OϤo�\/gps#�����񕗿�&�xno�(�(�[��]����6������u��'H���VB�t=��<��X,,]� ;B�Ɛ����.���^��ï�����q����,A������
jܜ:<�B�����������M|�O��>�.�Y��Q�70/	]����m��J]v��a���������E��!���r*wE�|iQI�����^�r���o~�K�K[KV:��a)����D��
�:\1v՜���7��߳L���YD@U�YEى8U)a!�>��M�f���R��P��X]An0Ag��Gä�{w�����4�X~"vsLu�f��l������b�d7fjҷD���!�
�A�����-��&0\����r��1�ӡahz���:u�d����sx����cf�f���C�!�K�l�\�V�l��k� ��%6�y0vIe���i�s���P�'m���:j�
��:�L~1ґ=���ci�$>��-�AO���J�!��+�B���7� �)}������ްG����{�غ���w�縘��q:@<6c8�Ė�T����Y�������K�&�P���
�Pk������2C��g�B!�qH�J����Ɯ�V���AJ5:��$}�Ab� �LF�k�PmF�?��~�w���	��\�q۬F���J5�K<K	`�K���޲,�8��|�(��ڸ���[�1?O)t��O�U��+ ����@���&��K���y:� ��;�����#G��������}9p�혗���3!Ul�$��!�g+�h-�˴5��g�<�ݶ��Iu�el�@<�^+�T	���ؽ�c=����UN�K�$pW�l�#��Ͳ=&�!7�X. �M�6�D�m��r7��`��G8B�D�K:��K�0�g`���\���\���$��\'��lT�<�I��������D���d߼{����j�aAr��D�}���!�D��k��5�5{-�<�N�������E\���t�����͗@��_��qfMb��?y	bV�9�CK"�V1ʩ��d��#M�Q U�:��wۻ�v{Rt  UsB���%��T��3q8wʼ��jc�������Id�dҠ'�j�o�|���Q!�)Y�K�K��g ��3�������Z�JH+��ھ�L��G��t'��UHf�7d�E�*�9kl�"��U3e+�oGn̥�C��5̞-..b���[woX��X,�Z��������kK����s���jz�����Z�|���{ElN�Ȇ#�����I@�&ͰQ�͝5���[�x�Q�[��nb&��&���ǣ<�ٶ2���.�<>�8�?]N��Nr��u��Mq����}�x��w��?�$M�0ۢFG�<$�q��y�@~owY~���Kx��\:y
��9��2 ��֫\�a9xO<1ŵ{�ߺ�{;YlwT:j�R����>��.~�7V���"~�_���Naq�rh��D�-$�� ?�{ϴ��w�<��%���Ӹxb	�ӼU�f�(k�ߛ�����B��8�������J�0����� �9�@ �7�����Y7��_��w������T�X��%Ti0��dl�5�j�4�CܹwW?�;kw]��YN�I�H��g2â��Ĉ�ͽ}4G�fyh�9,së�~�&ƃ]�T�#TI�p��{��ȧ��*���OWۏڸ�ķ��"y-�0�%#�;�ŋ E W���M%Ȫ�J�]	ʸHG�;�*a���(�Wy2Jl�t*f9Od�ĕw��M9nV>�tb=Nԩ��6JN_�V
�)�h�HY�$s0s�Nsa��g/T���<.��a�FEݯyIc+4�^0t�[|3�NƄ{�'E�!F��&GEQ�.@�v�1lvi�	T�#��w�L�����0�u��M��K�����N�@GéF��j�7.2�}F	�zn�|ߙnG]HRɏ	�?�t��S+���:$�]�Κ�Q!�H�ԜT�\@��,���9=�K��EAcor��b���U��cu�ep����z���\��eF��7��U�cǪ8��G�Ll�h�$�������E�fб(;b�]�/gK"����� 3!�0#���jJq"��CP�ĕY��ip�3���$|�5�P�H:(�;@��_��%5�X��3�mU�����R��(�U͚l��>: dq(���r��wm`�͐M�Ϝ�̭C�`v�l�_r�<�S��	7�ᦔHwoF���~��x�tr�5�?��0ɤç}�+"�Xwo=W����e��)�C�?��%����!�{�[���k����2���!z�����k��6�ϸ��j�׶̑2���Ql�������5�C4�w0iH�g��^��I��*�jzi�Ls��Թ����ߧ�ۀ*f�q���S�\�����-��i▲Kah�����˧qBM�{5�˴�,�����h�T%�<.p�{ζ+8OR�J��*�2��� ����tP�V�v����6<�o��I�ǵ�v=�R�QœNh���"Zq���K��aK� R	���&%է_,�D���&��&[�H<�ڥ����m�L�m\��U�cܼ��<�ub�ݮ��Op�����k��h�ܐ1��o�j�&'�	�%�����ӯ��~���f�����|��)�_*��D������A�����{>Y���a���v��ԓv6G�@"aJa[e�X%9|s����d���(Y�`R�H��@d`��ؼ�wb�tN7�����w�gv�(�d7j0;3������<�?ƭ��0�<_��/~���ʤ�x�����&�0rtEa��Av�^�~��3�m��<�礦=a��W����a�|���Hϟ=����P����� ��V
�=��m�OG���}�pRN҇���� #��"�/R�j��[��5ؽ��ׯ������=��8��g0?,*8RLe�����`�R�^��,�g�)�����n�K,�6EW�1����������۸y������T��.������X4��>�h<���9�«��p��-T�%^�$�)���R�DWJ	���H�C	�r��b��(S�Jb2?��?�����[�w�!�9R�>߯)]]��3ҏb��Ɠ��<�j�_w�srJ���`C�&2m�A/`d��A��+e�3YA��*{v��?T梍`��&~12�'U(��5�zn�G�DS��V��);��_���5��1SC�p,G>:k99M,�xЛm�	�Ö��������r�b�w:K|zgr� ��$�X�p�t��q�D7���S6e�1�V�f�ET�h��7��?�3�<�ԭ�Y�~�HPZ%M�j�@}˰��P��3�`w�ș5��lm}ZS��{}��F �Mʎ�7\�C'y8m�4+��9�M�H�]2�ƿ��^�tRQ�x�R�G,�*�	x��u?��j���.\���\�A�THd�j~�1��fB�	�v	\�5�~�˦}fd�!V�YoH�ޥSՠ @�N�K]���`A�V%I5g�G���7��y��G�`�JCqs�㲟��w���9ue�&�U�4e�uML���s��QU�^]�^P��Ͷ�ze��'G�JC��芷�74R�$�!G00���@��bX�e�vI�G|QH��TY{<uy�w�X�vZ�A;�.��8;5�W���F���ŵg쯣����c�JMq�L���!�C�p#*�X6�AF���ZP6�9Ӥ��|���j�ˮ�q����a��)`16CkNK�JS�������a��S��Md��)<w�$���B���	�����wKU���Ӂ�IW	p��XY�����K�R*�G�B����t���#<��`������W������V}eKyq���A1�5��4�]'dJ6M��t<�/���{\�^:e���Eڝ�䦐mwm�D��V$�cƁeU`V��<��A�1���(s>W��hχ>����%L�t�}G�#�m�{�@R�<j��a��i%�-��F�F`��|U%���	X'@zrw��jK"ۣ�,U����2Y����QZ[CW)�,à������GKm+�'jsZ��\�ZA�����%S��|x�����B8� +�G�'��{4�<w	�UIY�t�f��c�NL`c���O�����>��@u�V�����~��"�q�p$鳭���>�Ԫ#�y����×��8��;n��������~��b�h{z�����X� v�Ϊ�ȷj8ML
J�>8@���S���t��P�?*~C��I�F��l>� ��G�QD�u��)�`������[���."/�|�$��!~��
��w�emz��o��n�1�G$M����5����ҥ���g������9>X��*B��89�h�k:�&c�CoY.�`��W&*nNF=fw$��;wP����~��Wqse޹����
ԣ�� sf2g�P��S�
�y��e�Ztf�?��R��8�tu�;�51��FcEWm�P�|�v0`%�ǉ�hS"�3ҀG�?'�c��Eさw�^�:/W�F*1�Kk}Cؐ��Ri���-3
��h�]5��ȱ�^^F�g��*��F�E7�D�&��
��2�iV+�:�ejeB�����������j�7_����L���@�x�/�����[��ie�����w&��&~
���x���H
�lӂ:*NΆp~1���9�hZC	�9��s4�t���	Ty:�j�&Z�-F��u뛫���ml�V���[�J�C4�}j~�X�7�J��VX	�o��Bh:�0���)k�(Oӷ�q8��7D#>1}V�pz
1V������1��8+5��Xi�{᳇�=U�Q,�@��Z9�]8�8����XZ�!GG+J<h�|�l�|���<:͑����6���H��D��ʗ
�.�	��P)8��1t��҂7���4�A�	J#jS��iڕ�;��}O���^00% 7r�k�N����M�TΫ�l���7p MA��e�C�ݠ?�4��#[�/���M��x�ҽ]ǚ1�c*j�?����9e� �����n�̀���wW<دï�2�o�E6�9e�%��@��s��A�b|LQ�7;)&�t`�w44u؂�@��)8��.ꄏ�+,��/P��N�C��Ц& �yܪ��������?�S_�
�Z�0�=���?G��W�Y����e�tN'mX�g-']���'��r���\���I�,��$:�8ޮ�[��W���"\e����ީ��$�Bf���mT�PCm*}�F�����v�t����I|���jc��������Sq����B�*:����rG�25C[[J�0���$���c'�#J@:�dTn��-x��L�g�"�O
X|�iN7���N����vW�Q�|�s��Ǘ�{�>��}�Q�c�0��/���P��K�*��0}� ���&�(�<�/�2���d��Nf�IeQ�Ա��/2e�\��v��k�$FF���1ob���M����4�]�6��S�h+0�g�*��_����\����uK%����h����KI&��Ǿ����,��� ��5���j��,�ݟ��?���F������K������ya'ov,|:e#|���sXL����0��#|X�[A�oL�k(�5=IZ�e��g��o��^{E��}ll{�K�4rn��o��辉�|o��%:�%�b]t�i�+E'������`}��ֳ5�v�J����v)�L�L;�X*`��	���M�4F��/��k�1k��h$_Eg\�����ǝ�u\���߼��^��W}��L�t��7I���~C:�#���yFE)᾵z��\�q�hD�;H�Ŧ����ǆn�\\n�U��KVU&�����3"�T� ����<t���b9yJ$�`�QSa^��O����pk�����pݰʴ~dN�������^At��,�ǞF�0�����|�-�'��NeQ��!&n֬�Ac����?N T�/���g�vǍ�*��L�<�5�۔��q٦�k*�!�q�����t�wB��yo��Fn�V�K� }��!�u���"�>���GO�q�|� |�F1�Ǎ���-A/d���f�FɌ���:�Z�`��u�����H�O���ʅo�+n��*k�k{LGa��q���z>*��Uf~��	�u���	R�������1�L��^fQ�\d�=���� ���k��NvJ+�U�덉�E�rM���&	�6=�tp�4��a$�
�ڮ@*4tS�(���wg7�m��9:�B��[��Zvߞ-6�#�M��g�F<t���1�?����D'��0�T��U�K���WQf�^�A$�a>K�1��>��T0M��U�V�b���t��s"�NJ.���~��Q�s@�� Ǖ �@�]v6L�����zEa���7l�3������j?��P��!U���rw#*�-�񍻩4@f�&K�Y&;�PCp$X)XT#~XF~��Xb�l�(�������C��ˊ]P�(Gz�r=C��:�{�ٰ�gA�6��4��d<��$~Z=��������Ơ�I��q��@��w0��X&`����`P�UZk5�{�ӣC�{� <؝x�Q�C��]o7���`���Ý{�m{6�ƹ�4li�|N�����^wPGx沼�uOY/�}�¾�ؑ������eЂ7�tƱ�\�f3*����ܷA-Q8�ugD�u�_����1}�{q�}�o�V0ΔZߙ��U��;E�#T�g��Y�Q�9Q�V�6�ͳ]�G��>�=�8���;�]�gp?B+1��?���^��ˈq��S�؞�h�S�̨���6vJ\��y$��<"�]����F!�Q��9�&_(p?ɻ]��`c� S�H%&19�Es$��:�:b�M,���M�ԱJ�2޺��@4˽�E���Ź=Ԛ<	>��õ��?�!�����O�T6��h���?ܛ*�$���e�|����8�PQ����0�hv��Ymٛ4���;�7?���.��C�����=�lj`$�y�~��*�c8w��Clol�p�K��C�36E�Qn�P�R� �֐�>�gϞG����rQm@ع{�����Y�2	lm���s���}F^�׻h�����v�E��C<�ثH�����D�=.'�f��(�<\�V�O~��~:�T
���rB8=��#K�dX�����v7Y	�.�>(cck�b�	Yk�^(><4g�K��ɩI�Ifչ�A3sǐ�䰻���W�akcǸ�⡘�sK�"T�Usk� aH@5�(A�G�u��<����G� �Q�Y�-�	/��B�OL�GGV�X'����N��0�t�Wi��������� Qk����O`�Y��p���JӞ�����B��I���ۈ��,�Cc>���}~���xY�h`%=�����~����Q�[��Qyg4��,��S1�}�!yGn8��=<[v�F��#X*~h@�w�KPyT��5�;F=�T��VT)��qvy�Ĕ��=��&�Y*��	��{ulll`����{E"�%��x��h�;�q�kH"�cB�"��5tQ���<�1Rvm8����g,"��h�I9yo�;�������a&���OCzb�h܏6ֺ5�L�Mq��#���w�G=���aG�ǻ�F��4F��!��V\�2ʕ.��m<��	d�|�����$�<3�yL;�{{��gâ����v���H��	��?��q��G h��3�O�+-Fڳ(��38���#Y��F�]E!�0�[���ࠈ��<�}��6��|�eZ�$c�NU~�.��/�v�ש �>&����g8`���*Z��{xHwm�҇��30Vn����H���4�=^T�e�&�䮕xG`���s�"��i�F���\��ߵoY�nN���hw���Ƶ��X�L����M�?m�?Բ>LQ�����6�}w�}t��t��a���̒Ⱥ�~	��4JFm���ET����9������l��ms�_\��u�����غy������%��y7n�Ю#L'������S�^i1K_��ȁ-+���k4�������*�m���V q����xg��f�Nb*�è�9�����4$TB#E����~c/`�O
PzRs��Y~vU�@�2pcy|i���jE�P8q�J�z����8��3[i���SK�o9����6;*O�!B�fP�3�c.�hCt���]������?�}}+�;e��}8�5������\~�}��;8h5���7��?��X�xx�5�~p	�M�ΗI��K�F���ƥ���4�g��F�Ӎʁȼ�m|!#��z������_��7����hV����I���US�a$��G"�����|m�v~��-���;����~��_�_��i�Y��HrP��}Ϥq�������k������dC�[4[����4k1~N��r#��]�GF�� =߸��P'��E��!�уk���=՗ �~�������+X����"}��/�{(�teZ��)HV_����M���,NO�l>��r�%x���~:>���9���؁�R�z��C��/��j_��R�u�v�_ÄtN�a�ֺX���G�xd����3|�U����E0�8��9~��A�Bu,��&��8��é%��v��m�;���#�;�w�"Ϡ�@2����\<�����{��!*�+(d46t��^���km��΢.��Q�� hC���X$aeZM%F��\! �v��4��sg�y�x��x㭷	R��he��2���_5p򖪏(���^�۴�qM�ť�APZ' ��10�+���lr�h�7x8����	I�(Z�2܀!��_��
t����(���F~a5��O٦6�w�c��1U,ѩ隴�H4��2P��]DyP���&ff��r��&���~�z�f<�����*"�oAs�*?�p�-c��2���Fw04r��Y]c'#�(׼�3JBh��q1�����l�7h.d�%a=X���HY���ᠼki��'��t�]�r�n}��&?E�ˀB��݃\���+��pw����DlpC%�j�o �gm�F�q8��s�@���~�Hp�:-���3&JG�C�Xm*���]�M�������;;���M�c�e���#�T_G2u�L�>�m��.��gJ[Wi��2�ִ#B�Q���6��ģ��3'pb1ja�7���H���2�u��+�r8�����8�&����ry���y�����2��@SO^�V���U���h����o!�H�?��������/��������>x� �U�q���&��?H%��ݮ��q�5���:C���%�*��=詌������,�y��De�����
�p���`�q.�6�"�AI;�I}W�t�,���:a�#pM��5H%��~�d�rD}�Yp�hT�=T�ӲIi���=�ƙIɈ}�Ub\Xqqx��Dt5a�OH�6NE�$ú�T_%��ݝ�钷FNWZ�[�%Q��Zݖ���qt���n]̬��1��5I�g����B����wq���z8����(q�����f��Dt0�w���	n����zۜ��{�������K҆���2���l�Ϥq�@�j�J C{��XP�bi�A3�Z`����x(5�-��V�Lۖ6 ��N74L��RR����te�m�~<����r��{�4n���2R����|���pè�e��B���ʝ���B�o�=�s]	�����&af�~��י��'�ϻ���AϦ�5���)�}��%�U<��c6I0�h��ɹ�Z{��]���&���R�<2���%������S�����{w�s�3�l/�5���p�ǱO#�q/�TKZ��~��i0�v�.�h��MC�����6�%������tz����c>�ŭ��������AL/�����8�w��C�{e���l���crӅ	tx����_]Y��>��ӿ�%���h�B6rjB��,�tܚ����BU#M��{�
d��C3�C�Z��6
6�ox�i��%��(�K�RW��&?���U�����ҫ�ѯv1�=���y��}k�P�F� ������]��l�ѡm�=�盟���=�Gyn�7�a�:B?5��&�?@�z����hI�(�s���?��cg���h��@$^"2��W���7�D�ߊa�X
���26��x�F��\�ӗ\�ȴ[�#5�ב	�p�d
�p{���$�"���o}>��j/^�O#B�@S�i Z���}L���a86����ڣu^�{Xk��N,�Q��AF8s��kKil�;e��Y�|�gf1�J�ڵ�p�.6v]ɔQ��UvJ뼸i�qC.�s�C@�Ҡ8�F�YD�{�Vm�u(1r�]��?����Өo��ڦh��-R�L�e�3��k��v:��0O�>��H;7�a�X�P�m�Q��_m ��4�Ӂ���j��;�)*�z�����e��B��JG�&8G�UE5�*���7������D"N�l�J�N���F��CP��8��E'!��E�]4�Xg��������Z�9D<�W�k�O+'B����jJ�)g��1Ex9;hV��G�ߴLM���#�7?Xa�	l4Mɹta�S:�b�bB�Ak�]��3�1y�ol�=�AǕ�����9ȇ������0�y�;��򙶭뱃I��*�Bl�v�i�O*�y��M=k^vT������cp�gx�ʦ��#�P�ň�|�}K�.�E��C�Ս�oԸ���7������GA��Έ� �|׃��J� 0�қ4^��a���@��"���i��Gњ�������Cx4�aޅ�?��DE������|�y(��T[t�*�
xi�R�5�z9���xN�Ϧ��n���G����s@�SG�w.���x�d�j�
��<���Q9���?sjZ�v�ў�[��p&��3��� U9��̡��s�I˚˹�l�ɤ8��V�~TM�26
d�c����ˠ7�~�M�#�7�hi�z�\>lY��Q=yFCQe��u���q?F"~�Y4kmԔa�N�$�N�k�m�{Ь��)�_I:�vh��R�C� ;
cD���1�u{�6��d����L
[�*|Lq�
(�3�?:����;��Y�,�"�h���sy��r���y���TY�]�RU��P�ԩ�k�wҒ�2��.K<K{�
����<�*ۓ�Zu�mt��G�I� ~�*��AT.g2��k�h2������O`&��s�X�p=��D��z�kO%�S�7p�+u]�u�@��g���T�<"A����q�*;ח�a��	_�c:hu�6� E��k�m�㑩Y�NO�� ,L���ţ��'׭�v�ϷS�`���F��,s���g��$������3FU�S+��[C�ϓMO�)�N��<�YYO

G���]�T�]8}Ҩ����0*�0��`JA����^z��ݍ��q漇���ӧ�<7]�������(���%���я�w�?
��i����������R\��?���'u�{}G=f��C�6�<.?s�7t����!�]����~�M��:rL���|c�4S��͎����[�x��+��;�q�֊��l��P�S�gX~�&�T�����F�(�C0/��H,����X$�h_�����x��-I�����c=yF3�s|^!��V�!=�l(��D�<���l������m\��A�G�XG{��o�q�\��l	e�����*vNoO�U_��d��a|2�(�4��h$ⷾ��C���:/S/�F,��hL�7�(��	�<<�h˧#����c����Z��sި-D)�LN�F�ȸ�j��%)>ɓ�3g�?���P,�P��YSy�z�F����*z6�`5�+�t��M����D�<t`I��JK�Ƶ�/,��h���ul�[d����vD�4�~��A�g��hr4N㞽� ImP���u�ͨJ��CNi�wxP�����e(Oq��b��9`��F��<f+�����i�eHOR8N��|�{�� Ͷ���,|b���J���{�\Ild�F�{"�P���Gz�Uʘ4R����Q�!���N��!�=qg9�������&��$�*u����}|p���oV�Б������Б�Q��=�GWB}p�?�ù9�c��kK��<�#`��{I���S��ᴹ_-e�M��ᦋ���~�__W���?#FWa��&E�KM���:�4>�>~�g���*a�9g
3�9l���?D�<M�%�m:�@=_˸}����{�/�\< �<��Ѱ �2�uF�Y�C1Txv6VVp��9�����8~q�r	�j�����7�P��%C)#������d��V�J|y�Q�N���k:2Z��i�o��}����|�_�*�&s(|�dO.c*�7=�6�
��l!�J�Ѵ�EN]mUj;�	l��df��Ƕ��$
���Ǚ7R�n����gq}���e���	�g���/2h+8�`Z��4 -��j�&`]B��_��h�@@Z���=s��A�@.E��oPUF*�|&�ʄ�6D�_+�#X�sMg&�$�h�E�[�`�vM(�d�@��a���\#: �]sWiL���ы�by��^�nf��/�T*c=���*UD�ˠ�N�` �k6�-m��M$��9���ڠo���
�Ari��}ӌ�L��yz6D&�䂒�S����u�����Tg =�s�������x���xX�ڡ�j3Z�,c���6 �~=��!���cπ;g�&$�< �H*3����T�
���`�l�2���b&�ll4��G���g��������~�C�����6��~��Μ:�ϟ>�M���y�Q�S��?�W����H�|�������'N������)\�ro��㾩����O�q�`3ŵ�E�����6c��1$�̭V �k��=yE����U�c�x0�.�fu��ڙ{��_���n�H�2~�	���ci��'z���m$��x��$��+���1�,�PRtk���~�S�u�
>��5|��E�v�5p܂f�W��$P0�u�/"c���f���;jh��g���y'M?ٺ�b%x��Cb������wW���&C�1�:���u����,|�]C�[%���窤�_����cxa~Ӵ���wpPe���kHt��_�ܓ7���r�*jq�7q��&:+�hfF���ml!��w�Q�"*/��O�b�|��g�H%���D&�Z�m%#�l,�g�ƹ�g�� ��g����߸��u|�i�r�'�qc7�ap��(��<�޺���;�G�>��	��7�wn�P�E���(��9�gI��D����s����?��r�[�����QT	E:��J͌�x��4\qجzCx�<e�z6#	יF|ǟ��pu[ֳ`L}�^�a��e����++w�k[QV� �U�YԲ8�p��:t`�(: 7�kJL�ϵ��^D{�4��� �E]x�k��j.�"�S��2���UwQ�U���M�z�����*�m V�"͟��5H�IƌY?��g��C�����<�S��k�^�Ƽv�>��"�̓����`1e�R����jX�7R�Y������=s."L#Wܩڔ�M =�cm�������"n�ee�����Mg�+�:�F�17�i���2�>�>z�FGO����R���L.�\E ��������0m�M�>A� =�1>��{�O�BC�w��x)�i�cY/������g���Y(1���s�LD���yO��ڪZ�h4���l5=��Y����8ǟ��_�p�����6��&e ��a�d�光��/���Ү8?������o��Q�uro��Qѡ�TY���p:�=���Z~×��=�ZY��S�!:��;����ƾI���W���1�	5k�+بבP��� � !97�[/����׬��[k`*�1�C$l\s���J :G���<����/|
�O\��{k�ں$wjF�4B<7�a����>�[o�0i���H�.��3Ϡ���[����ӱ4�-뭋�5�*^5����:�s�T
�u�6j*˖kHҦ>����]�hC�&g�պ�t@�A٨�Y����k��N��}���k�[�8�Db���Sf2E��X�]V)�F`����7��o|�Q�������wiOo��;�?�6�+? E�&����ZM�D���Y���:��_�����M�*[6��Mτ��"����k�`еË#�'H}�������˗�����{Ys��#UD4a�1bߺ�e j���,x��d�zg�x�\�����L��o��6�&eU����~^Ӗ}ss�������2�)>'�vhж���y��w�s���}\���k����/���6VjE<=�!4�5��{q��q��_�:��Wo�B[�|�?Â�x�o�˘��<�90�ѤY�W�o�W���h��!�����z��]�s�)�qb�����%S��1l����͟��:�jc��c*���|���|��A�g_�v��I��3�н��ͽ}|�������̓x��2�f�Ȥ��{�Z�d!�!+�i|���\{#ױp̯�C�p(Ӱ�h�{~��#\�^�n������7q�A��CՖb�F�T�ZtUV9R�����x���a����<ǟ'fYT�v�>:��P%�i�����������U��cJ�q���)�:�w���������L��6|1.�9>�Bdol�v?��^�`��&�������1�T0���/����T���	Fz)�֭|�o>d�u�s�Lb����o�	�����4L��i0*�@ןA4�{�����l.��[��Kkؿ��)��a,#�0=u���ir6Yw����@�uWZYI$Κv��N�����:L�!�h\�tC��rPa���Ӡw�4\=�^/_�o:�D�t73����cmm���(;����oM��P�s��p"�͍.�i�t���&��!z��hT�I`u��yzv�L��#®���f��p��y����t�b�+�WR�s4���u��F���xOh
*=߽��k0�P]���~�8��׮�����L�x��8���ex$Ť��h(j��`@����^��"×��%,�A6��0t�4��(�w�x��>������t	����=4Z?2�0݋�h��;��=�+q���!�st0x��8�4]	��oG:��_��ݟǓ�HȦ��8��f�y�>����f�����B=�o��{<����er��2=ԁ�i��N+���f� ns�1�8�@:��N�G�36y\*����� ���ߔD��2�`�<l@�(H\���\�{�%�DЩ,T����n�or��q���q�������ف��;],�/d2�k��N>�t@�@4GQ�߇�1r��a��D4e=g��A��Gx�F~L��ɟBz�֕���_�	wP��|���݉����F<�B�QC]�U���X,��2�x�g/�Y����:�=��5 �PIY41�ɥY�q��m����6�x	�z	Kg�0�g������nD�*�!)_O��o]��[����kw���˘;>�J�O��E2�0�)�txG�FaC/R����@�.�
���x>�զ�C��gҀj̿J0�)`�1=ϐ ��D
_y�	,.G�>�ƻ���_�^��!��úUT��m�z�dBr=�X��Q��h���s�8~��g�����ۯ6����MG�%���$`mSP6f������O��+/�� YYS]���Rv�:PDR�|�gTUy	'l�^=ӿ���(�w;��cS�R�h�g��*�;��|ԏdwR�%c>Q��L��/w~��m�@����Dg6\f�f8����N���P����;�$��1E��7uK6�	���Y-����_z�%�	ԟ����R����*�d:o��2�>�8����g��{[�P�(��ԇX���Q�����'����K�	N���S&�6�s�x&�Y�{}�8��T~
#��ɈJ��E�R{�ۃ ^��^�a��'��f1�����7�L�^m�Ɗ����oS�%K���\�J/��2>�zg�paq���ƅ��*�?�A;jj���g����.��sRrC�+��#�=h����n��W�	�n��C�)�_e��~�g���t��)ޯ��{#� �P�� ~af���I���i�b�0�ggf��ġ���,"�E,����:��w���[A���av��H6���r���(��RD#�~�A�jM|�9L�B�J�]��O�W���_C_����al����y��3ˌ���|�Ҿ�^���G��5�*[��W
89�7�~�n�4F�;��.s��1{�c$F48�!�VeX���M�F��hJ!�c�g����m�͹��O�(J�ˀ�Q�QO����(i#�"GU?K���1�<�K�Q��h�4ET���VA�_X�'t<���Mlom�9�0G�;��ٙ�%k�c�'p�X���Idi�K�4�RQ+=M�c���X���&9�jF?07��YM�m�b��g��2	�g{����M�7�,���*��Ma�NYYж�	:�g���1��Gu��@��9l:vxG�umy��o��>�W�kXm�P��*U�(�M`��)������hŬ\�y��R���Fq%k����M���2"*9�9B����Q��aF�����օ�k������ӆ�_�S篏���\��~S�O��ɉ<��Y����(�7�rS����0|�|��+�wd=��%3��:���v����ogmd��pȜ��.]_�D�,��<J�w�y��� �S#��C��V���g3���TG��4�G�mV���j��+�J=:���"?���c�r"�.r���\�;�w�&Z�mo`���D�X���h�zP=���E�EZӨ�|��NVO�.�(0��/�D���G��qo�ZG������T���w�Pkv�J�O@�l�?����%��P���E�k�}��?ML�q}�VZ{��W����Q��ﻢ���idg������a6U�����+�P[]!��ܳ����mլm�yDPY�XO��F�PĈpLa�}��w�� ��`gS�$��O�[��3�Ҁ�`�U�6��]�F��ы"���'�������E�P�|]���%,?~ww�q��U�[˺���`_<�p.��O���sx����+�+W���)�
,?��)\��>�{��C��K�R$��ZZ:��r���*��y������#��Z�ܼ��{�����a��T$�,R�k�z���C�����^�O:��M�O�w;u�ζ�2UՈ��,���������<A���2��[��Z����K��O�i�wy�D��S'�?�Zp��X4��*����l ��A�ā�tSSS��i��6U����0�����`��S'&��.�h0�AL�ϑ&`A�o�3�Hg�g0�J�}c����+�9�����'|�e�ſ��q�m�eh�����]ܽ�~M�[�M,�?ۉ�y<��#���k�������,��3^��U��߰����ժ5��	�S�@��!��a:Ap����H�\k�kt����K1�pn��� �X_��f�����p�j	���ȑ�B�tX�V�g&��T�v/��6����6�/�#��U�
*�� i$Þ��T�o�5�w1������q��k�p����Y��;�{%���'#�p�7�Trޤ�B���_1��}�S��'''2��l�bo���R	ub/� d2�g����T�K�[�A�&���a��q?�M��q[��������CY9\�}�<e��GV�g}8�����v�b��͠�X���nn�'�NY��2#F�M�Q��E.��Z���A7��/~��	��6��߻�(,,L����`e���,�+�*�s�.&rA|��X��d�535O{&J�� ����6��^��t�HUin9%e�c�s=J�5�E�J��Д�J��g�Z��+3 �p��Z0*9�q^VF��4�iMW���[�;H�s���!G$�����B?Jp��D�p�?���d"բ��2�\��*f���_z�q��Gx k�L�9�׮���<���,ff�h䢘���St�����H��j<�%���ލ�.����[v*����'xp+w>�)���?Z�|����>ٕ���;������:��:����G<ͨ���Qn$��A�Ý�.�mTz�ӘϦ�#�.�r��(��t��!M ��l\D4$A�{TI�Ibvw�5��Qb�W�tv��?Gi���E�����0#��?�ԧ7F�j]�����܌�Mu�5�%�����p��c*E���`e��:NI��h@�<K���5	�z�q@��H�m~`b\�U��M<q.K��H�Է��ηz��tN~D���X%��(b|cXw��2B@�J�����YB�¼�p;���cS��8u�"*u�Q��je�&q���K{�7��k�����./$
�W��r@ܸ��E�}���tc�M8�4��sb�����e���
����o�4�g�M�Ã|�3sx����n��pk!��Y:��^�`��sS8�8�/|��]8���y^��4n5k8x�����l*�2�g�c ����]	a��v��k��/ F'�?6�!�B� pc:�M:䟼}#�1�h8ͳ�׋D�%��ER�/=���7��WǞ����~��isy�Rʬv��yt��v���Xʥ1{rݥ4i"�!R��#^���.`��s���E�"m�w�s\��[n?���K���3O=����oi�5	��/������9l����C��u�25��D��F�Nrr��=ɟ�]xc�>W��ĉ��>� E�4���5R1��1s��)��bk[�qŴ���I���*�3�{T<�:�H����6.^ ���g�O�\�����>תK�F��� ��}��3�"M�ʇ$�m�������t�;���(��X���feѶ�@e��)W,D:��Q��\���iL�lk$�9L��*�����i<9�@@�E��Y|n�>���k��v��w�� �,z��o��k��N٩F{��7N-��B0�������0r�R�ڌ��>�Q�=Q�?��`�@��+�FP}�́���ܟr��B���A^���vFx�e�{U<��>��M˂$;���o�q�f�A�z)�|�1hZV -S;O�p�wJ\�ݲ��z9���f�����Oar�8f&f�1����d��6�) u��Z��_��|/�r��iP�Y� C?�a�>?{�[�L��tF�S/��3���7�Z
�q���+wP�:4]�8/����,>����n����{|��c�wG���+�Z�J��Ѩ�[����&gެgƸ�Do�qa�A�od�r@CM~��ܫUbI�l}��g�9�1ӟƅi?��6�4}7T�L{���ʸ���Dl��.�9�n5J�X���	^�e�A����/>;�Xt����sFQ�^�/��b�M}�����=�~�^�ԤǪ��UH�Bѥ4dݎ�cK:G��MW$#��V�N��PiWM�b\bT=���O�591_�J#�䥔�8�"���Ӻl���Fŝ#q �8��� @�)��<|��D��M��0i�XT��l9k��;�V����\���?�b��8ň&H#��k�+Ep�B���"��/�
����Өk��^����� %��hh�(1r���2`ʶx6d�v�����#��(�3W9��
��m���Ϝ�\�Y���Ԭ��X���> �X����;[e�:��'��IQ�/�������y��5���q�F堁�ե��!ʽ������}�Y�>��Q (虶����P�}hA�44��c�s��c��KU� ���Ky�db��t%^�4}��������̘"�֣KN/�ް��Hڨ����z�zG����z����&��P"�r��a�i`�B:���T��UX�18:Z�#)1���v%�!�J�db�v��&&
)<���t��x���.q���z�qD&Rx�U���_a��{F[q����X������Q��>ϱhL4par�4�EF�%�_K���w�?2�c�8���>V��ߧ#��D<�5�Ͽ��Ŀ�y�����LG3����D�;4��k�k������8AǢ�{�>21�{����X40!z'�V�A�����7�%p���n_������=�'�X�>��?�+��^bP���$N_����߶ra<����plj���ыX�i��j�N�ş����qg��|8��/.�C� ��p2���[8�|���?@4?�`4���r�T�/��&�˗pP:�i����{��"lK��go���� ��215�r� �A-�����#9��7�����,|�����bo^��>�����U5�n�8���gIe���^A��=T�=vW�`_Y:`��k�B�@�R��W�(�b�F�Ap�N���;5 ض�J6:�Z�Y�w���PKis�f��i�aS�w�T�"�/`ba��ح5��m��lU�S%�&��� &4�2Ǡ~��N����k����!�:/1�_]��l8�O?���R4N�@�p��Y��K:1p�n�L6�Ӿ�ci�m|�_�o�F����ھ&AP�뷰_��s<_3�Z��5̍�W^Ǉ�
��x��jz���`^�P��v�*3�梽����GQ��-թ5!����CгM@/����,�8�:A1��N�=\����wcx�)�˓Ce�!�y,� ��
�����F�羰� �lAD�:�\|:�c�]�����`"��O��{��s-Kx�E��$B�r[�/Ó��t�����+�\����N[�?�_nI�`�8$D �4"�/UFlȔXi�P ��Җ�x�S����	$S��m��λtk}�̉X ���,�	����=�^}��<?q�����6e ��@[C\�1�_J^)!��Me�>⡏���?3��H��pT�JcA@��^�bJ����02& �i�`u��F�w�$:x���q�(p������a�*�ǿZ��gf���^\C�� 1� �oȊ������z/<9O��|�����%M�IRj�jW����_qg���dB�at�]�d����.��z���5�TIC$X+��%L=pb�}Nh�`dl�4
����U���C���e�Eg��<~lYF�]:���s�n���"��֚8�׉�����nּ�������(��4/|�F"�U^����֪Ȫ�|�F���M�'��EC��P���[�^�J��ǜ2��#�0Zǖ�ߺ�+\�"�?��p)*X�K��FA��<th�N~�}��z=;��v�g�y���	h�gQ��e\��g�RzO��F�<r����u<u�#�,�}q��=�v�pg�i^��oq+ �Gak���T�XՄ�rG��IT"=5	�B&>�#��g\d�]=5�A�\�t�.n�0Ňvg�/M�hd߯K�;�3�LߔA`�yq::�d��,<d6����F����z�¨ֻh�JL���,:m3J69�q9��- #:
��7_4����Q�d�3��ʖģt*����d�ZnrY|h�
H�W"���XY��9�Å��KH��lZ�R�y\7SB�'�(�Nc�֠�����ukA��ē�2
�w:�R��B>�]x^�C����/��\��ƙ��;��ŕ۷��Y`��BP�|ſ?'!�67��Щ������Ѥ"�7��u��8j� ����}3�8�wdSs�	hOG�q�IW��7��0��콍2��s	����M�	Zz�SF��5{֘�ַ���;�^���'Na6����"ʷ���]��(�#��,����&~����N4�?�	R����c/ 3�c��w��ܿ|��ck{7.��H?�|6��"�Tܡ��X�c'h����G$Z���x}�����������&ї�,�M:���^{�.FkC��b9�:2�#��W׭�O�,��l[�Ð6e�@B���t�{�f��-ʞ��Xb@����i�3�Ndl.�,�\��ԗF���{�E��6�u���=ލ"��6��NY��y�B1�z~}j��*M}}m���*LӁgy�v�E��v���Dk���P�O\*'�š��n�`˂���<�H��VĂ߀������������m#����6������D��v��l��5y|���e��FJ��%��1�Ĉ���¤���̗ą-$ә� ��"�g�H�6􃨽�>�"�M�v�����cϦw5M,#��3�}�=A��ss��j��*� ��mp����޲`�=p���q_pO}�#׆��*s�u��f��49�t�USB���&�{��i��{����uL--b�0I$\¨��\*���$����._�U�����d0?��g.�0����?�����$_���k�����ŃX^�bqN>+��+\�����7����-l��À�vn�k��;UTvob��Y|��������:����8@���s΢EPM��_�z�4�{�����e_��v��������g,�q�m�|���g�!�c&��S�x�@�po�+{�z��ܷ�B�W�HuV�*)AFS�t~�]U.����'%,�
Ǥm��Ҍ������N�5�FS|��'�L�s�	>������4*�v��A:5�#�L%����j{���4�h4�қ��-��N��S��pEX�}�7Z�}o��wk�f6P�("��`n�`�n���+]\_m�>������m��a����MȌ5}�X�����ﱞ �ЌB�H�D��"\4���pL��s�c�#���D.��������8�4�!:��C]S�-��X��%/nC�#Ǖ/��Q���T�t�ϗ0zeP���t[&����j�i�K�ƃ^������Fp]|����h���l"V�|��)�����	D�]jWP\A����?�g�����{�L�>\���	Xfg�8�ƙ;M7*
ՐA�
��{��e�=�p�Q:��^�/O��s���J�������w�˷LV�U�˞e�<��x�xEݿ)8Q�!1���B_)~�nwRT�"=�M_�+�%����C��qN��(]�1�w]���M�9r�иi��@�/pD"�]/���y�!�������'n8�d�P��=Q*hJ��;��M=h�K٬�PG��|?�A�������.���*ml�q��"�H[�6駒��5I��H���_�*���I`�� �\zp4]��\����JٙI�׷Q]Y�S�)�,����^�)��a�lO��{� ޗ&	��<�4�~}~8�he|���i����C��Z7�baħA�Ŋ�58�v��~?��K��g!�x�4�g��⩥Yx�4j����qS���Hq?���<���@����x�'Y>o���=������2��9��t(�/�M�nRQ|�������ϝ@�G�t�Q���`��,J0�JD��+��h����Q���v��A����E�*��&�|x:�X���^�Ak��E5������A��+���g�YR�(�y�5�F@9��0��!/�|��l�Z���e���M�VJ�ܼI óvwUtU�G��,a:UPb�P
�'h�ÓX>q�T����n2���4�hYPv��)���1��N�A_t_��<�K|�F�	S}�m�&C���v˘[��g��@�z��.d�sW�-1����ȏ�s��e.B`�q��HI�vM�Y|�g�x�|�a��vo\<��K��I���l� ��as͆t
������)$�yd�)K:؝�����Q&Lw�L`����}��$�j8G"�7�:U%tO���'�*"�W�7rj*'�����9�r�E��$�HU��*>�a�@v�@�����-g4Z�.l�Cټ���؛[v^�a��s���7��zn ��$@� �g��刢��*R�������JU~8v9�d˪J��Z�$J�D�N 1O��F�Û�;���Z�;��!Q��ѯ߽���|��k���. ��hU�0i|�x��z��Ξ~ �o���a�Ft��V�*ı03��|�/.�g?�@�����1�ڗ�⾅q���������/���bf锘h'0k}̧�qr�C.޲��{�q\����y���zٞA��T���=n`�����Uٕ=�:�����x�|�f�w8O;��	_��sc������@8�sq~�@�����Dnܼ�� b�vd��,'�f� ��1�M��H�b�I�&j��Pj��>����k������&,�NW*Qa��jT��Hu[�P4%���i<|��j�nv1EC�ب0�Kaaj[<��Hn�J�2n��B���a�楓������x�]��8��� �M2ҋ32WK�Jv��v�F>:f$�H���Ft/�Y��p+
xɝ�E�7���H�j�R4�l̨{T`rN ��jZg���	e,$b�P�˃���L�3����.:����}�:fs	�"+i������p�⍄����p�3N���f���qK��-�p�6ec:\Þ��d�������Q�:����u$�>\�J!�wݻ�*����g!�>��Im=ҿ��s$�}�m�a��̟"Q:��KUY&s�^�N˅�4CP2��+�iR�[�-E�[� ն�X��t��I{�][X�c*!i\ͩ�i�W$Ig:f%rǙ�ln�5�x������xR�]�� �5�;҉�+���\2��Ct5}�n�3��`x�7�����G��aw�kV�I6��7�N׭L�K��'L4d��R M�rq�I_��Ic9  �.U��cĿK'��1������`��F+���� i�D���ЄGh�6P���U<t|�Κwՠ=��A�N �~W<2ܣ8j����@�3���̾e���$���qmm��b���b��}ZZn�^���/�o�-F�-�;=�����~*����v��՝N��{�w�|���ƘIޥ!�#>V��y�c*�z��p�R��R�P�/x�pm��/�{��&�:��+��O|g��AEɦY��h��[�V哙�9������ϱ���=S7�elr�h7��ħ��yܞ�@݈K9���0{��Eܸ��z����6n5�������'������w���$9	RM�PV�i]ư���K�۵��	��i*�Y(�/<�#S��%����)>c����
���/��k?���"t���e�GOO��?�S�/`||�,�<c�S�\?�f����_~���+�|V	׈%�v}����i��Eڋ�G��j�_��M����a������Z�����?��I����۸�b��-�Լ@���s��i�guq������g��j��e�{�c�����O~�L�Z����i���m�,����C:�IU�5�ҾSuG�=�>������� 7���&�XX����+����L��b� �PATZMG�H�L�0=���	�=^�;m7�b�v���mӻ�[.���>��ɠޣ�$���l�ao��}���OE���kYk	Q���k�M7���c���5�e��F۲V	��Ilw,8T�W�� fbͦB�JZ�S�AzW�EMc�MU���v����ny'��1���=�rG��`�H��&.o�p�A����{UͦN��o����I|�s�~?å[%��@��F67�d$���E�׬�*j�v7bغ}���'�q߉���n�A]��o'�Ah��)~Nm���O&1�L����� ���d�l�.(�?���9X3Aq�u�LMO.�:
ք��{[<o�6�Qg�i��$M׃'�p�x��f�[(�?�5�c R%��D����`�����̓8:�O|+�KL�ml ���Df�D�6S��*��C�?�����?�޹��K+��$��HM���{�9�|��(���Z�����=T�u+���#�k5bV�V��E�F�h�T����wc�IB0�mT�V'�u���4B��wMR�����$L)����G��F�u`�]mZ���m'���.:�I��t���]:$�+�5�ūQ˼$h��1�"���<.eN�0껷E]�*����Q7A�K \oz:l-�g����PS}�K0�1��秇�Dy�&�=AOS�p�O��T��2Ջ!C�4�缒Lb��@^�>��l���GÛ�9!�w?#�[`�6��y�d�h6���f����}&РqF�(��
�Py��аV��4i��D�5�2m�̝��N񟀶v6�Z�A�d�j@�6�+z&+�I����'Y�a^�	�4-E��:����)>�7�}�0+�k�������O��:�^����õ)�z���I��:�K
��-ܢ'���u�8�L����$��ae��*�"e��4�(q:_Ј9�嶲Qq5�m0�=]aĕ�u5��(�W���u�'��*e%(�4��*������Qq�xwB���jK�T4}@]�5�h�:-���ss(,�O:����ȟ%Қfѵ�{���Xr�4�f{�N��t`������0��h:*X��آ�zU�����iF����&��.j��9�g{>�XI�n��N<£�C*]��v���e�D���m��⯾�WVz���$�qF�4t�~�f���t�QWꗌ�fV����o\���k�x衇������}w�\�Laى	����]�X_w��"pVeh�������ʛ&�!���s��_��_Ň���ȥ2n<�>_<����mZ�h{c�_}�z��8�q�4O�<��~�,�~���8��8Y4۝e��0=���^ďn��3�����Jq:o½'�5��:�՝�
������Ǟؕ�#��M�[�_���<5���#��C�ظ��1��v��m��{��5��r��*��
���þu��������|�&T�����vy;{�>���E&Ҙ�ӷ1:���F&��Gy��^~[�ⱊ��������7^����E�gJִ�)Π���^>�ڵ>�ϟC�`9�ɇσv�!N��\'P��v�R*��s����f��$�{�g*˚�WkF�@ԨIeݬ��w[�.���|ݟ��:�)�NtV���-7vN�8�}ޫ�`�0p6P������U�6�V�E�Yb���6�]m�ͽ-LY�Q�%>����$�s�*}ʆ�'�<{�[M<����� _�峘_��g>�1ܿ{���m\�v`�7�F��u������^���eB`�e�/N��?{s�q�����+��47pP�P�Ǒ/4�<��N`�v���ڨSM�ir���g�� ��� �r����=��o���$��X:jMv���8)��5D���E	b5>��h�4������nt��￝��� o��[|&mt��4d�~��H|�~����c��!Y�A񙧑��ƥ�=��,��<?��SO�n������:r>�gS�H>�K�cs)�iM7G�����l>§�$�u~.�q{`=����4mZB'h����d�zg36�����i?7����Pm���ְ#~U��=�Ӗ�}��o���kD�NY��mx�n�&G�̥�UNf���pшGh�w��x��t��p�t�:��0�C����̩hM\7� 
�KH �!A0W�V��+����[@q~K�Nc���g*�$��o��$��no�����&��zw%~&�����2�tӁg'l�T���+���O���m,����D�N�Ļ��0�WQ&CC�;�rjnjK����j1���ڡ�I�=I��63���D�D�U&��:�yk�R{��F<m%�U�4T��%ʰ���S���s�x6��rѮe�R���(���$W�9�RR��N�Q��d�w]�<Xrp�g�c��' ��-�" �ƒ���8w����3�^�vD/ǱqA����Y���]�w��+lIN"n����M/p��
h }��V,׬�Jam�Q&M��礹ʞ�K�qW~�F��ݍ�d�b�n����eF���~��NC'�"����ٶJ; Ĭ��Ƌ�
�6�$��升A�>���Q$�������ٹ������?F����qs��Թ�����u��i�b�L]�x�)>�a��������+�C�:�ݰϜz$�SI'�?5~*M`>˽�óV�e�^Z���_��;�X9�l�����\�=>>���w��70�J��'��D��v�b��^�_�.�&�Z����(�Q鞏��&�<f�n���)����7����l����އk ��$�G��+W���;t<L��^�!B[�oIo���A�_r��|�P5�^��#'qxk�h+Ss�uҙ��p��>�,b�x�{�{����T��D4c�>���+(�j��j�F�P�G������S?����y��|��w7��i6n�>a�zyq�cX�ۻ6�@��ࠃ?��o�;?z��v�w��3*B�T���S'�n�G�,�-�ũ$��>&ǋ�|���qcc��r�FۨQo��dM�--'0?>�=�M���[\:~���������H��o���"�����1?����y�����'�M��m��V�f�e{Dl��S�N�I|:��F�1��1�a�g���5���}�ý;��x,E0��}��fsD����R�ΚV�%J�Q�bDF�\�,;.a����6U�g�- ( <�SN�X����A�lJ(ɆF��5��i�y�|a%GTj+��2]��lb��T�Ua�n
]>���v�y�s����N`��af�f��^�Qپ�ܗ�9h+�nU�5��>}e�"$��'>����1��չo����ʕm���2����5v�k�qt/а@X7��an|	+��y�������˷4���a-�t��U՚����d��<L�s��-��C�މC��"6&O�c	i�j$�Ɵi�HgQ��f���(6�a�;A���j�ʨ���mL.Oc�7�[����`�ó��O����_{��.z���X[C��<�;��I,���G�r������Z�N��D9M̓��=�{tz%����~y�FY��7lO['kV�XC~i=��Tޓ��&��	�����I_X�D�mF�O�G+�6$[<��+Ҹ�{2���x��.SV(Ńݯ7�,�aq���I_O )b���i���{�ݽY<WN}?7QN����b�̓97��Na鑳�X\B�Q��"\{���i�����'P;�1��!�����>?^L�ge3w�݋�����er�_�P�g�����U���]�������-��\�iF��D�ՠ�
��\���[�v׷Q�9>������ ��F��`�/(�Y���"���X�/b,��X�D��/eL�t�@O��1Ꚗ���ܔ /:4���C}@�6"�A�+�G�Ycv\IZ3Y���ͶE`�����u,lNY��2L)m"R���	��*,Vό��I)���톍�(����J{�/�y�2>�j� NCÇI���k�A^���J5�;Cl6�Z�cX�[�J<p�a�)j���T�ٷ6���"�i��L��G���p -�Ѫ��GsGY#9��=ݣ��'2�3G���ٿ�+����y�C?��4>65�e�s�g�����ߏ/��W޳Ⴛ��IAY�c��x\�x����K��k������.�qp�2:��3���\�;���x��/�8��@r>��x�HGQ�4@��zq�(R�ǝ�6#�
H���Gzr�8��v�*������=��V-a��TZ������F*�A�|�	��67����)��������9�^���r��r��6NJ���1�l�^yHer�η����2�?j;�I�P=��q��s�}�2�[�X����6�$�|<��R������^y	����vP�<���v�g�6��lZo�cyӂ�`@��ޮUpzjTH��\����^	Mejwwx=��С���R8w�:��dhww闊�4f�܇.Aû{�����Q����V�	zÈ�7�9׉��/b��5��R��"�\�4�����B*o���s��՜t=����W>��v�gI������*/.�������Ƴ�z.�ګ�2׿��X;|�x"�w�{ۇ;f���5��o��R
H�͖e5*Sk֦��0hH�x6~��[wg�~HP1=�CaB�LMa�p�}q�i��Ryԏ۞׾Ѭ�XH�E�=Xwϗe{i�:�w?v�;N���X�5��駤������r��FL�.�*�K�"�N����0ǘJ'	�`Ҏ2����H�J��7�o��=��w.��>@:7�����l��'�B���"2\M�ZE��M��Ɩ&v�K�ȃ9L�v��3'���4�嘕���5~�@m�6e�M*>n�=õV9��g��rXj���M���[�?��jZq�2�c�~g�>艹L�<�޻���UL������o"w���o|Pi�j�MEdx��K`=�R�tW�i42rd��ί{]��|�:z�]D*{n�xeaz��U�Nj���gQڸ�^��n�*bܜ"��U�ύ#���]�m�DV�9�ET�)*u#ç�7���Fil&
�����h{Vv�/��5^S߬�7t
�*fun��g���)�I�}h���V�|���q��Q�-�)a%�47��4%B47n��(Jd�v�ƛQ�u��Y�f���O/΋�B��=��rrj8軲�����H��Jze�8�<�Q�|�,��3V��r�	|$�(������<�����,�� q��'p��o���hHC����֭'�&��sp˦��dJ(c�':��p3��a�ɘ�ڈ���e]���%́��/��vD}F=�J!^�R|����5�4Z}5��ۖ�R�P<�\�-�y� Q,M�2;NCO��t��4�$��V�����v�������Jߓx�$5Rtv�0�ڦ�,��NE�wdJ�J#�r��t�
:T�VT����9�'a��зk�9�4���14���kk�Ҧ�nnπ|����eN�;��*FP�aD?l�x�9}a�G���vj(�x���U�������g�{=�^X"��9� 0�T	����VnЈ����Z� �22&������6����6�q�s"��M�P�v�}�2xI�pMg��I�K�1��`��n��g|��T���ܛ�U0#}��d�:|]S�k4q"�ʙ���P�>�Ȇ&���y���.2t�	���߯Q��xg�ޏ��N@��Uf��c���I���}�=�s�L7��F})X�8���
�Ⱥ��J�q��d`��ɜQNp������E�F0�/�ho�غR�هD� ���kv6���}��^~�v�f�N�A0�c�mqM��W����/��Xǎ��7Z�`>���i����*���EMR	&��3��ﯾ��n��*�8����9�\��=�}Bg��4�6!ۨi#$��[G�`����^�DF4�a��Z�3^6O?�5�Ͱ).V�>�nS4]$3�E��B�q�*�}s���/��'>���U�������9���~k��y��:n�{�	&[�qF���Q�S�����Ѓg-I�i�J�=��6���ͷ,{;����^8��F�8�`d���cܵ,�Be}��Ҫ2��]�ǹO{q��<�����hzJ���" �[\0���az��5�l��llX��m�6�I��3�n�\:��>\l)��U�f�������RU���3T����J�jvӗ:�Ah����9l��o�/��:
�s���d�D{Q2&p���ǧnԁ �M�#�]�PIW�*�o�0E����϶�#��p�ǍիX��s���ҁ�h޽��+������N_xr�v���=��Y�9ڕRM3��X�~�%F�9| :�����&�L<� ��x�ǹkQ�b��Gr8�lZ �z{�������t���������X�9z�0���2������>��u�ڽh9��]L6m�[#a/pX�#깾 �v_�k�p1��9 ����{��.h5�4)aGo�	#\��;�}+��}����U�G��F��͡�mX��y/�:([Hr3g{��7��s�`�\���I�8yԕ�i�x�KF$h���!�[Cie���-7��D�������IZcCހ�V�P�jġ�n6.^��P>��dz̄��6Y��Z���y�ؒhX��5,;3��G���?�Ng�����o ǚ�|�+v�M�ȍ����3��?A��1T��v-f"�MY`�,�ĝ5&�{����)�c����S8y��������`ZQ9���\��7�B6����N����]99�v�#��]�� �RC��\����uu1:�Z�����uU��ج��.Z�?���eĭH������O�8���x�8��&�҈�웉!��[����E �U�3�a*M��։ ��3O��9�\�ԇ���:0##���L�f�K�����Or�[�m�x`��!%Hie��n�ʵ���9VMVПƇ�HZ��2����z��|��d5��G�P��PSQ�SGЬZ	��)~k��T?��b��6#�f���m��?��[\�a�^�D�8~��D�''aQw⺪K����wxk4��'`�^p��~��A����ɢ�xqo�۽���+�`e5z��{���Dq���Ag���4(]�[R8��~Nb'M`���){FE����V�	ռUnV����P//�K�z�Eh�m"�M�r�fK����`vvy�����6�T*�-���/<����?q�+�ޅ.�\���_2�*C���1�0隁�w����i����K�5NO>˽���N�}�q�|�7�ؑ������m����ݭV��_�6��U�XM̨T�0�Y�T�X}nߺb<��1���nlD179���[��F�������G[��,�l��2�?_T�>}@�kK�b����oq:���N�}�e���Mp���4si`����r�"���d��˝j��Ui�����]i�k�1u�^{{{�s�J�6�\��qq�l���{7�$�=�~u�hc�p">䥭+�q�&�����G��[�p����	k4l�z4w9-[A;��%Lx����� O�f�z�u+�k>��N�kQ��e���]��B��@�{�>Fz���8{�>,��q���X]���ڴ{|v�o^��W�̷
����=��򠤗�T1!�&��`>"YC�
5�D"!/�qua�gT�j6k�I�h���(�`6�v�D��h��Ц�(;g�$՝�w͇ҵ���qe��W�k8M�PBh|z�g7�v�JPXc�?ĭ��nLĸv��|.V��`��s��o�����̑�h���N���x�'��E�FǗ=��q��)T�M�no������*g����o�����ݵ�K}SGpu��y^C��z,>���c�&Z��<���k�T��*9��µ<��Mj'ǵT�ܳ@{�H�RXW]г���1�ϛ�j����,��@�h��+uoQ��i�����JG��Θ���,�|`ͷ�!�'��اpm�j�,"��	&�&�ƨ���ぱ�4g&���^�8miq��=�J��a�ňm@T���&���E�"�Hf:��g��2��)�;��	�7���\d���ԁ�$�W��F����4���Dsq��;� U����ωY��U�+o��M��cQ7kq�Ni�4e�F�"^��;P%����x@��^���<LG�M�{�a<�˿����r�ԉ��f����, �����M��F�Jh�d��=$��x�~��cx������~J�i`r���dRܥp�.�1ͬ$c�(Ҿ�
�us�P4�$�2��*Ŀ�A�P�ݧ��k��j'mE���wf婨�����k�0Kt��� �}P'��O��v�dB�EΌ��xgOM���4��|��P�Y+��J�Qe��h$��n5�cհi�N �09��"<��h����wKˮl%�������s�"�Be��\2��(�YW��t/��{FPdl}��17@��/_�s�G���F� ��v��^b�X��5gX�+���a0��^��LLo�*�d�n�R��|�1�j4�� �!&<,�U��.���[�7�Y��j�O۵&�'��T����ǵ5�6�1b�ݲba�Ýp�@�oYݽ����(\�'�v�îqy��,�^�yi|zv	G$�KФ�2�h=���OYͨV��T�y=����VVФnO?<cDհ8=?����avhL́�)�W�7�^2���)�����ȹ%&4�����>o3�������X���8r47�i>�N�f �-|^qc�:V�X�\ٔ+�j�к|	 �q�[�3��x�6�3�8�ll����ի����P.W�& A���}��:�+ N�fܮ��Ӊ�3��j���ni��Z���rio��H�z����Γ���>�~��E�Ӡ�֐9�+�q�$��,o�����C��$֬���N�+G�8tԅr>��r�"^��A����S0�q�ju��rH4\,}�?j�&Թ~~1���9�?�.^}�U���Yd�ٮ�u/�M:n׮zX5!nq��3����O��m霶z����ؚM����:Xs�i�hτ��*�ݗ�\�W�:��Y���gZ����F�%����v�*	s����f�v�������.�����,#ȣ�<���9�w���}������c�?�[pIЛ̸�H޻u�
ת
@ ��ךL+PZ�I�%KԄ�"H6ʎ&^�&j�K��8�J�͑��J����OcogS3����]gT��O:��$��*���d�ġ���2���ɁK�2��@ET!裺�iM,�����Ck��Ls]E!�8w�'����^qO�ow�R ��w��c�K���C��3�fW7�h�P�X!�q�X�c���<��6�a��ꭷM��;h��O�X\� sz�<3�*��ȼG �����6�iv�u�=B�!�+�+�'�v�'Zf.S�Gzf�b�Y�y�*��6��˛����l� '/�И��<?؋ǭ�*�2�����m$ol��\m���O`pm7^}cS�x����2n�{��x��x��O N#Ҽ����-쭯��{�3Ԙ)/�{�Q9�-���B�$h�GC� 0C�! T�eih�Ւ����I3"�9z�#u:�,�C�g�h�~�!�{�w��i�̑&E�W	F	���"�$J��-�7��������-$x���t�#���N=�V��W1�У��2��9Z�Dei��Pu���N�L2+���HJ�_�4T[mn��x|�K������QjWl��$�ҨƓ�{6|���0���ᤊHx�ሷ8�߳�� ĸ��	�����y.y��ɰ�2��4*NK������$����E0�*��8�R��Ըu��H{a�Ek �."/$�:zf6�0f����HYJ�	!'# 5y�p��2F�7�}����iJ)DK�Ģ��r���_�{�ul�P&��j@�*�ڣk�����*������c8[W�oK���@���Fve�rm��3�7eiЃ8
~��٣Q��{��	]t��	:on��5p���Ԉ=s�v���=�w���2�z6�x`��5�8�:�4�(L�\�E��iz��������[[�p(.�2�4�.��"�䞞�ͨ��юX�F�m���_���N�˪��/��$b��kx���Uy��:{�>�#9�rK� ��11]�fv{	$�.�ݶ��e�(-�w���~��^���S�'����oz�.���`�  ��IDAT9��Gb�hNHgVYG'�5G���t&��"��XCC"�F�Y���̃�����>��ڪj @�q�:�o��vp�3t��d=:�l>�|�aR6���bI���]��kϮV������ѣx���H��D��j�.6޵i=⿵�\��q�lr��#�эhdL��N�#�EGԐ��-�~�q/љ�x�⇙
B�@{߸���Y
b����j��afi������?�,�z�)\�r��A�Nۣ�����A��#1V��W���m8-�OP�������Xu��/� ��{��1�Ҏ��!hV�`�Q�Y1�ܘ����VP��nz'�дVeo���|�z����ג�T�|���.��8v�4._��w�_�d&k��CuJG���MKRp���[�Zπ�����=�v}��Ě,Pg (N�\��E�S	�ͦ=T�~fr��~6>1�*�~�}X2�Z-�x:\���.�3���%-�;<tKv �_�8�b�p�S�s�tH������֡�K\^ӧ���-��YⅈMzh��D�eڕ]M��U����������_��m�hJ�"�6m"�4�J[�Ȇ͘�S�O����iX�o4�\<i�?u�9>��uV���Ho1�IC�~V��qՕ9�Uܓd�=['�4d#mV�+�(]ȇ)K�n8Z�X�R���= ox�W**!�PAgV*�DݚY!�-0�0띸���4����6�Q�~�~Az�Q�$�\��یD	��J�ƦgB�"��s	R���CY�����g��U3�B��e2Fĝ"����Ē�(�)>U�3�"9J�T4f�uE����=�;$���.�4����9!� )�P��	(ǂQ�.�	צ�;�+�qQ�l�����V���t����N]��8��O`�SX��@HF^ire��=,��ʹ�]6�����t1u��C_i���bcؤ}�0?��g>�̕�X�yL�
�r���ȠH�=������RRi,����5j]ǑP�3>�<d:zwhG�L.�*�$G���R���<���Wi?���u���J�"��(�YI�3�8�4��G��������V����u����[� J����W�N���;4!��/�ukJ��"�TĚk���nшqL`
�N���b�%�@`���,�Ѧ�S�� ���������#A��o��*a�!	���n��No�}�
�v��}��hhiX���L����n1
�ƌ�Ф�Z$�H�Ñ#I�sȖ�(�X��`���Tr׶�n;AC����E��=���x�ʘKHu�ī���±grr�Җ���A���逿QY�&�҇"�y���|jb+�~	���#���A��q#:�����tk%	FF�eܝq�54)`�Z��F��5��1fYY�;4���v��4bs�&�ׯ�Ѧ���;��KXY^�?��_�̍�i��.����ui~qod����eZd�7��B��U���'�Ȼ#�#	��e�~��iT���*�r�Hװ�i�駟�W~�K�|�2���r�8>����{��?�~}|�C��f��� �C�P��a�Ο7��];{�V9M6D��q^_��3>�\*��M�0� ����
n���+�c��T1�'9�H]����ű8Z��^��Y=��~��mV�L��4#jP<H;:�*
9]ɞ��#F�6A�,�W��@��4@s��
�����ams�<�	���>��X����,�`LY*���'8+�]�A��h���q��i�I�ƭ[(L��j@*�NP&j,�,�!��B&�c1�K�Z����>�H]�2�r��E�<�h���z���������6����2��n���mM�q^��e���]@-~v4�-�Q*��t�=�6�Q�'<�b ��Y��h6�eϓ����>�!2�C��ʽ��&-S��|T���k�����#@>�KW�D�D�ʑ�r�_�H&J]��2|]�u_�%��a�J՚�Q3�~
��,"A�kY!ȣ�hzH�����h~+��mI�7&���%t�	�Ʈ��:m������$R��n��vbCA���]���{��&�)r���q5�)�8�r̽�kFAp'y�*Vu�5�@�+s]�V�F��{�0f#���ûk�j<��/�	�:��*�<�Q|�Q!Y"h�u�2�'V�;�@D��G�]��@e���t��G�d16/�ǐFhA�)\��!ߚ�D;�����lm��hTs��@<�~r��>���YM_`"u#>���!������ZܣKf#���n�[K,Ԗ�����h\�B��{�P߷A�d�G)JG���F3Q]ס1�{ks���G1y�A��j�+�X���h�Kp��e�ܔ%�8O2�:~�(��w�K�)���H"�[ۻ8B���~�m������{�LmĲ�nB�֪��IX�+G"I.²9�a��?�ל�="��>��c1z�H���W�w[�R$��LWS%�D'�M���1,LM!�LZ�ֲnC������]�Dax(F���e�F�P�4�ʵ��E�N�O׭=�N�?U*h�\�fw�4���g--��v�eT�P�6*Ah�WI��w"�=4=>�~*A������Y@�ѫÀ���޹L�4��P��`m��2�
n���\/�k�7'ڐ��)p��לe�M��2%�j��x �C��<�@��A�+���j"��zI���-��΋���U\�=���2��y�^_\-	��?�Ǔs���P+��`͋i�I�$^d�W������}3��s��O���N睿�N�Ѥ��~�v��S� Q:�R�G�/�f,:�6��P`�Q��=���(S���I�$m����M\!xU��ĉNb�EXa0��`��N�Jk�!v���L�ķ,^$�w��Y�����������2�}mo�f[_e��.f�9&i��z����+���B�Q�Ji�qڍ�zo�T��yڊ�j  ��'��$�9��3�/e�U߯I�M�`�T���*��u6���5���uV�>���h)�U�G3��*���YN*��������[x�����
C:�6�w�z^Q��x��^��Їk��[�gs�K|�˼��~gϞ��e��{��?A�l���1��}��
(�5��R���Lз����:����	k���/�#|��_�A� oi�(}��r��|?:r�S�ײh0���P���o�w��W�����T��X"�� ���Hw�����#x����s��ƛ������̬���V����j�gV�Ͳ�\o5 (	\6L@&N���9֤���Z�e���j��7o�S�Bٯ��~�s���EW��x�7�^ϸ���'��U�r�8|�_ђ��?��:���K���p	СrC���D���T]���tJ��F�ҀϦ]F,"o9�c����hk����4C^�:Uhocև̳��1J.ؔ���;���L��v��{�p�����6
5���K-*�X(�e��Y#o`�'ǝ���.�0��`B��I[A�y�=Q�� t�^�%O���@6`��O��
�LGR"|pQ:���f�?���#�=q��W��Y��cb�n_|1F���M$._2ܠ���NF�WQ��N}1�	��^D% �f�B���y�He�1UܢA��k���rD]����Vi<f$d("�nj�iK5ZV��,�� �� "�(��s��ꦩ�&�F9m+�nR������=���r������ʑA$��ߕى8x���6�����ԃ[��,�?�a4�pʕ�����h0��Ԅ9��_?{�E�cO3w��q�vp������x��=�!3X��m�X$#��c���ă���/<�7�ݠ�+�0P/��i�ѽ��UZC���JV3�8j�P�@�ɥ�F������!�C6��)�1g�=�&�L�[U����+}X63ģ��4����&�^�O����R��u�dMC�[	��i��fiG39}F�Q��=fs��+2�z(QES��t�4q�h�ڣI���]�a}��a�-#�s�αF�9�4�H��u��=��H���1>a� Bb�~ǳ���5�G(���1'�"c�o��\<8�6��T�cQ�WE���@kߍ(��6V-�(-��v���΁�g�޶��"_��'��_���JZ����{p�3�'�����7�5�[疀iH���{:3����?D"�� c�A��AC�q��0�
h��?�~�5��5<�"|k3nڈFiY���A�2e�S�����o�r�l�����ieV[Ve�Gi���@j*=)�A�������<��0�y��V�����n��8�*�3�B]A��3��F]�v��&_I���i/�\^���a�@l&���1���z�ş���q~a��� ���sh�2P����yl�O����6�;�@���l"��`*E�D Ю{�H��m\:��~�L
��w?ݬZ}C����*N�N��bI�VK�-��q��9���S��{%K ���5���:^^[E����po��V�~��5��!!�4
�Q��:�mDa�`�I:����tc}5��\�~���ۻ��,�ߧ�eycǺ�3}�\ѤI*����fm�n�W�k����J�\���}k�и+ii�(��r�Eܸ�����������̓!��ʌ��ơ�}h6���f�7����}$���>�S��v�*&h�?�ϸ�%׮16��x���I����SH�?O+ߋY*����g tze�fb���'&Q��1��,1 �{�޸N,����4>��g�fpP*ar��k�]ƫ/�l�T23�������77p��M�xz�۫���ivɲ��L���Gt �vZ+�ϑ��o�D���kO��M�.VD�=��b����C5�%0L&��$�3P�. ��UG/�9R���M�8��'��!�Kh|���?��`�� �[���ĥ��*���%�wM�D���8��c�\���+��U���~�w�nԡo���Ϥݬ��U��h1^��8���$a�([d
��)�ͫ��7��[{(h��`fj�J�t!.�aw����"Z��!��C@�����Bh�+�G?�D��k��&nh���I��u���hF����r��<����a'阒'�HF-Ke`�Z��aR�nF(2����"���8E�G[4�G�d��ߜ�O�:���r����$#1�A�{K�] Іև�R)�!�a�в����c�n�ܱ!�C̜} ���qs�L��f�?��ME��~�}�Y��A\��+sh6$���́��vw��w�g��S��E�)ݧQ���4|Z�f��+?�A�Ca���*�A���QD�,�"i��ӅM��	[�G%&�ю{��"q7-0�	��H�D5�����-�]�:�NO��<��?��,#_��jv1�����]�XRM)�Y�&F��>�-'�-�. �){���T�u%)Ӧ�:m{f�v���lD���Q��E�6ngҿ�d�ƭ�aoE�M=T�P��Գ,��8�~S4��8��YÀ���v�M$��	�:M��p��)j4�������*�͜��e
l�@*R���DՄ10QU??n���!��Iiuu���Q�A�����kLH�n��K��Jk���\v7j+���0�x}�ml�[x��Q� K �s�9|(����t�b*�z�1�r��i*H>E�IQ�n���n�/�!H}�2���MS�c|�Sc��{��k�V���2��+_�e���*Ddo/�hi:eM���?���n�\�g_3��1{��t� �A���X�d�j�g���l�2>#�AXʳ�}ǝ��iv���9��sS8��<rFr�*�N~��_7R�&>$�i�>y�33��\��O 11�[�%���Xn�h-�f��rro6�n'�;�.k ������mQ%�yl7P!�H<�k�'ҡ�Y������e+�S����,.�l �~�>�����v�:ӏ?���v�`L��ʉ�T)�Y͔�����y��"�!б.E�ƥS'��3����}�I%��}�+_Ƴ���|V��mRYL����-1peԤ��H�k��r���y��u�����jT��ݱ츸][ۼ���e��-���V4�	��TI@%�Y�W��B� N�C���:��x���XYY��K�����4Y�2�)��f�4]�;Π�������V:c����v���U}P����<~�W�
/�7��:��ӧO�E����o��������kU����{;����u�{����׌���������0��O�#<��o��~���l�O���}��<m�	�y#�w���NMH`���V�OMiN�i�_߂ψ�ax����:�D����d�ES��#3�b�qra"D�n ^�t$��^i��n�� ��$�l{�C,�0/��s�Y�	�����J,H5'.�$T���{,�i���.�H�jF��&�~������>��{��lD����<�Zeg�&�1���먽�24j�rK�j�T��7�B�{[�w}�������z�h�A��L�ҋ�ܽ�a�4�I2f-bG��vh��ZUg`�$I?c�&��<oj���,��Td`��M,n䐛��n��Y�xp�~F�����j(6�n��;���7i�Nd�It"qb)��-}=��FR"��|�u��:�bwH���89>��A~�� Lp��xՆĎ,�Ǉ)9u�����q�i�	���[�W^��u�u�	�VmX��P(��ɓXY^��˗p��E�:}G��;#N����qPo��n!�����Ө��H?�1<4��ޛ�b��3���M�[��ސ΄w����O*;X��t�|[/�!:��и�6����t[F4�gI��!���M���mќ�Z�G�ȃ�x��<���a]0rm�W���Pg�N��,���j�'��P�zCS!4h\綦�D�SN��>�X-�r2p��$?pe�������Yv@��Qĉ����2�7*�91c��I�q�4�B���	�w^�ؕ_㞛���B�լ�ƻ�q�J���3[��8�L*�(.����ٔo ?�ʘVU.ýG��;7d�C?Ip���n�u��QH��<V�`.K��~���D?�d$�q�g��u\c���uR��(#+i��S���W/���v��:)��I��S�y|yf�j	�F&C3���$��?t]g�az>VZ	B����'��������*��Q���(���7`��Y�;�2�]��w{uhd�����~�,�iw����q������f�f3�����븴�߻X�6��������f�F����������K��Id	r��T	��:�L&>�fa*�'�@ˇ�>�{�a���/����~�8�t?�̧��'>ac|�f�,-��� �ka���\��̓O��b��m�d������k��S|h���#܃C����>�q,Ο�s��FuP��N��b �lV���5��'5��a{U^�r� 7h�~���]��v��׉���b�s�x��_G�୷_���o=�aP�$E�2��J	�g���=�?�Y7֐#PTc�k�Lң�>�'?�6S� ��-�ÝL�lV�|?���(f3��}~?�'����J����K��1��t5���xݸ��59=������_�^�s-��&	��V�#�u�qm�='R/�|Uo�1�q��٣� �����|������;����U�}�98��Ą��,�|j6�/��װ~�&^��,{��.�F����{����Ҟ�{6�`��b��q<��k��������G�y_�'���?�^[��g���������Z9{��뿊�������u{�Q<�����ό�+��O�x��l޺� �7��@6�7xw�H���r��2z��A.�����Ѵ>�N���B\`{��݉;p�a�]�g��Z�pLǤ��Vf�ԙI��%nB���>�����~�a��\Qk�P?�'�G�����@��]�`�!�bD�K��늷�[`��
��F��ߪ��7���@VzV�/b O|H�)�nٺ��z�|bv�F�Lt�����@�C���Q:���
#���&vW��0bX��������<�A�H�"�w�y4�;D�$Q��1-$�S�%�+�Ӄ�S����iL�ݕ0�)�%CQ����I�Д��b��к�pw ��w3R������kx/G phY嫦�`�x�YBˤA�iG�Ϣˢ�d����-t����R��$� �jЯZtP��F��SG
cH�/��	����z{�[�秐���q(�ψ.�JZ�H݋��^�U|�?�Q�`�Q��A�\`s�����պ���"_�v�n�Ʊ3GM�4�t`טTJ��	��]��p�S�22�.A�Ʃ�y�U�ݞ���a�u�N�(�f"σQ�3�W���S�U6����x/ޞ��u5�a����g�'-�6N�<�>��9�V��R�������L��SY�6V�v��TF���aɓԒI]�)#աS��Sk�2�*��M�����f-;�]dyW٭�IFJ��6�G;D���f���!��v%���O���]��e���k�1���	�Lq�M|��<#��۵���	9:��\¸Vri���b��t^9�z�b�Ě4P�t!ˠ��pR q2���b���(�aŇqkuˎ��NC�����wA���xe�)��x��{�޺V�AF�������,~��q,q����9=�'9e��M����-<3�6N��e+{C�U��w���r��x���d��X�5�m^��N�����t��4�S��	:{�l_9���kx��?�m�)H���X����soڳ�v��e������a��n{h���ߏ�I���x�_'�r���zɺ���M[Mg�*�E���������ɕ�I�4	uFJ�?h���_��m$���j������mS	t�j���w~�w��H�pS��}fK'�1���d�u��M[{�kWW��O�"x,�):���cx��gyo=�RE�L�9�(qrbތ���y����=+=��~�%L>�A,������S=�O�X����|��J��������0�1�p�d	��v�}�x�s��k＋�o���F6�^���|�[8���(2�V%���A�������v}�� �W�ߟ[c�d5����m�no�����CYZ��#t�5��d.�'��8��e��w�VU����Uڞ�u=�i��鴫.q���>9�ua`�5Y<z��i��t�?M��\|���>.^~Ӆ	��9��zyӓS�r�g�������<^��x��/�����*yy��jø��� ����W�#�|?~��x�M��^����W��c�O�M����ş������l�ͽ���=��(�����&^��q@༳u'N����%��-�ڕ���$.hO�ڡ�p�2&R"Fٹ3�@4
�)�Q����]��wwj	�|�܁ӉV�^�H�]�l,�/�C�ʾ�
�h�.�;������2���=e��"B�b2Uє��g��u;9]gk1��݁kS�M�.b�h��4�s�.&�/*����<��	&*��jE�TJ�S�*(�F5`1����=@OvH�Y�ywGo9��G���sS���^�m�9�CB����;q��ţ��B�	g�!�r4)�2U��>l5��\6�;�DN�E��sn�lq�1���^�� ���$b"�kV�fG$��")V�0�;tu�Ƚꨒe�i1�G8P��5&J%�EzrD'$�YE�N��U������N����o���42 �g���8�� �����n��n���On�η.�M��?������ҝ*r'�̎�☙^�4y�jH�r�D&�>C�Cae��8�CD��2;�"g�m]_E�Q�X1��j�&DD�)�x5E�D���tq
9�b����^�������)�8���E�A022p'uteM�Ł=/L��s5�^<�N�=iS�-�m`�B���}"��]:���,~�8�<t>x��A��1vsԶ�ʠ�L��a��!v+�T���*��[m���_V�bi>p�xF�U��8����>,���4J����Y�u�!�Da��3h;�~G��W?4|"�����}�j��뺲�DtG�o���È��D�2}R��s�'��-F�0�(�,Nbv��ٙ�i���J�&<�<ۘ�Y�и֏O����P�>ă�d���6uL�Ƹ���T�K����u>��.��7��h�I�K�o�g�?7��9���۫�Ѵ����&�aYT�����Q�i�8ϴ(]�;K�#%�Y�yLj��M��+*�IWb��o��o޸��`�ydi�������KI�tr���C�����o�hi@��D�����'������>�,�[6�����L����q��u��u�ӈ��Iq����&�pd��q���	kK�mw{������{�]6~k��5�Vs�у'��|��obuu�d�٥�Cڕ���.����<>�jW�rUk,<� >�����8���,��D�p��=<��J�[x��[XۮbqQ�&��ro��Z~�ԯ�2����7q�u��
�qd��\ۊ#��-����g�e�u��}9��U�]�s��0��@R�(�aY$�D.�6������c��ey-ɲ$Z�l�&)K�@� B �f0���ӹ:T/�����绯��g Q~X���޽���s�I{�7�X�y��+��E|�W���.��r���^�l�,Ӧ=�2�ة�c��;r��S
z��Ch�ZA���<������mS�&)FP�"�z��	<y�<6���^�}���=sdb�vr����w�vٸQ��ؙ�	�ҮLF�u��<f̡�i��YT6���-��uppg?�����3=g�p�6�?�{()��`�N��+�A��΢vi	w����3g��_�y���n�!���Ћ"ь�F3Y��[}��?�k����������`Ij)A�Sk7,�ؒ�i)M�X�M�ِa����>m�d=�ϧ?�,R�������7��F�~$wlGΞ���3X����7���<L?��5��Ų-\�F�����7�iuQJ��6Tiz���4$�˔�|�il�63�I�z!��&�[����J�M�nH��h��׸�X��*o�yʸI����606Z[����1Q��S,y�M�;��85���|��0y���hʂ���hh�#zvS�ns0n�QS��� ZI/e���Դ�G/�a����
�DW�s��V�g�ؚو�r�w�;(�J�X�z&x.ґ�i�O+u���2y����f3�4 6&/j	�d��>�ē8��h[頋Q}`>I �#-OF�^��U��QF��ASW�f�ξc5lM5f�#��9�.C�^�c�U�ȑ�*`��p���I���H���RhFw���w��FO"|��o֫�d�gd��(��J*���xn�!�z7�U��F��{��?r�����x;"���N��N�����2#�J�I�;S�8�-0΢,�c"]���aG��mT��ѧ�T6�������ǝe��ҽm�tTȦh`}:q 9����15ݡ�A4,�3�^[=j�R.o��A� Q�ʯ��΄���� ��%�MF�p}=�[ƙ:'��z���Q��)�n6O��Mv���ʒ����hq]k[=l���PF>=��F�+[�X�a�:��v5����5I�)�L:�KD�Ѷ�S�����`�c��8��܋�����?>�w�_�.�{�9��[o��S�ZZj>� |o`��e���h�(��Fh�'ؽ���T>�SG�h<	4���@�G�d9)ál��tg������A��l
�t��;m�k�t��r	�\����ܻj5׾��g�09�OLϠ�nb{}�>S%��9e���eZ�+M�/�@xQ��ы��xn_I�P��5	'�Aq}x��39k��0�����ΰo}�Mڋ-f>}���8�/�9�����k��ԗng�ػG�c{{O��?�Ǿ��z�i��u\���I����5��#���������o۔cZ��<���y|��?�g?�)�<�$�����WB�ە��y~�[�ǿ�{��;8Yxؾ�,�&H�������S�a�@si������k��\���/� �Fw�6�7Ͷ��9ڕ1}��H�;��)���>ߢ�\g�hQ�	�&����\��Un>�ݡ2�q�o1�ڸ�SgC�kѡ�\o!���JPf���5�ο�=<��S����L'�5��Q ,-T�+7n��^�m>��L���}k��6fRY|�c��_����|�(��Wt����"�������a�w�7��P�����#ϘsV)6�������s��0A����k��ͯ�
X������s>x�<�C��BYN���Z<f�k|��o_E��}bXDV���:�f�X�����g��� &�s��Bc�fI�R^\�I��+k<7w޼��_~��S��.ۤ��b9�-��Ϊ ��N坢���lNj���9<}�<>K�-:���.}����"��Uܢgyꓟ����8y�(�޺�?��?B��q�\{w���pvg>�穩Ix��i�?��VrT+H��4_�2�>?7���m�̅���C�{~��E+^��m�rm�NG��m�����a�GNR|梐Q���R]���g�E��e�UfVI����q��sZd���z��1�FF4%�?�>17i����\WQF%D#��䩚�P�G��[�NYԸq�������;ٯAtv��{]��X/�&��q�I��r�'����1}[x����:b�6r�)EW%Ӱ��:ecf��ړgY�����Hn+j.�fR:Uc�!��,��爚{֛�S;w�H�4�ˉ�{}4��˞U]H��ƹ=�]ɸ�,5�K�:-��/�����#���+M*}:rJ�Oڼ������c��2�rT����:�*r�S�90o�z�����jc�Vh[&�������R��R�fO^��yOJ��h N�q[��3�h/3����2�t�5:�8#�
��=,<x1F-a�� 78��~g���G��OW��ҭ��-#2n���8vG�l6���8��'��O�}���X:�3�t��j�eY0�?��l�Z���~90�1���}@�ۇl��^$k�h�ynJ�w|5�J �W/a �I���T/��3�x&;�m�P]�ߪ(�٪�$�~�R�`m��m"����hD���g�� +��~=5���}�t�Q{�sS����e��ş�ƥ������/����G��f=��a�_�)qo`=����r[�-��>AU�N[���1+-x�$ivx��~�������(k�+�(H���3��y�nob�w!���]�6Ȅр����r_�/[�V�|�������4����u�׌�,�������
�C�襕����ݔ�[0��8l\y~���=j�ġg`5Ϳ%(Y'�|�ļt��s�M�~��6m�!��g'�`����K���e�4G�>>�h���R
[�D���⧞՜)f�������8����{���W����^���4���G'%��ܤ��4�l�w5|�>��^�٢c*�9x�>[)��|�;M����s����|�v"m��	I��Gf�T�P&w��#���������sK9^699���M�*�$`@^oV�MS�*�5z-�x����7�����o��iߩ����7�kH%�.����z����~�@�%��&1 � n�Q��\���_>uʀ�����'G�P�����`���^zw^��2A�t��:�-=�'����q��<�y�Z�$����ݗ��/�͗^ķ��E���eRH�RhZX^[�)�A�����	��'y��Ss�o����CG������8��N.�y�Z�[]8���C���\�J�����z�!�����7�d�3-��mY4P&�o6���D��K�d�������MZ�G��m�2H���K�,�-! ��N�a�Cg2%<3u����VE+�>}[�7G4������b� ����Z���¯�=�<�,~8���S��G��o���W�`����V�s�!J�Gqf���b=ÓP]�g���?y)���V~�`���Q!���-\����#���[(�'	V�i��	�cG�^[<7����h�c����U��)ђ���a<o�B֗(×���_-)x!��Բ���*��Uҏ(�6um���tÕ��e�]�4�* K\�\��4z-+úJ���ޫ���Y��H��,�/��]">��ϝ�9�q-xK���޻���H��s"�B!�^:f��s�� ϋ���>G� )� 2��Qj���o�1�d9���vw��"7d
7�6�(-e��p�&�w��fG$�Yސ&NF�Q�w�������|�����~��\_������q�$��p�Τ��Œu��U�r���L���AT�Ξ8��x�:�E��=n�nh��J�zcZR  @��\�����ɟ`d#���J ���i����F��NM8e���VSo0��<�bد�����o�����/}�*<��|�F��+4�I<��I+��n���-��d��ZZ<IK�䓏W���z�*G�Ĉ�QH�R)~O� ?������p�+9����'����2���1���p����f|'͓�d��\�����[�K��D���zu��	Z��ܡc�V���
�EG���܅Zý�G��Uу�@G��aT܃V㽢�SU�7����D^�ӿ�y���O��hً��}Sj�J����Y�w#����m䆊��wK�t�&�.�p���ؑ�|���h��T�x�[�7�_f3$]䚕!c�U���,44Ȗ���b� >����z��5m0��%��:P�US�ɋ	P�9hߟ�)$"^��v{(c��T�+Ä�ÎRq3�x��)4hDW�'Ē�dP�tq�T�<��W�b���������a����gZ=�5���{���l61���s5�F��"�ͷ߶�da��i�
(�J�Z�����B�cET 3�� �PP���~��{�b��e��SFJ�M��G��d��J�䈧�z�D/d����N�J��t�&A�F���	r|��l4*��pjR���y�7-K���Q(������W���W�������`P��]2Z���5T�-�<��5�	@��)�ٙ�j�,�^1	D����)�)diߕe;S8���2�^zٔ�b3�L�����O�;/b���:�Q��T'�.�@�*4�>Š�^ma�P��*�\/--�O��5x�)�L�X�Gӊ��U�����KXz�
<�����t�6�'Jn��w�^�h�@f�<�&��\�0���"���z��W%����	�������N�J����W��w^�*�Z3���*.\��I�7��f)(�Z8�}�<���"�P�|m�d����k�ں��������s����۬��gq�˟��f/�������2y�:���!���x���,fGE��&�D���o|��87Kb����@�r�����H�;�w._��K�~2�R�/�l��P��͞�.5u����wcO��j�P�&1nT�mxB@OD�J(�ޮ�6�ݲ?Ӝ�^�㑊�hE��L;}�y?O��\ ��TG�Fdj��7œ�����l�`�KƊ���sдrn�$`14<Jp��zTi�&�%��b�s��f�=d�hTN�d�q�#��y� i�?�!w������5&��(�8�ʼ�[˛�d�Ȟ��pby���w��"���HS��jƌ�Rٓ8�Z�<F���D����$і��� �w�v�LnGK#00"�Xl/�1L$�"��۽4z=:��|��l�n�㋟W�L1R`�ʃ5dd��)��ƨ��@����Y�Z��)Q��`�ʡ#+���7�P�������{�M�{�r���@NΗ�l2;�4��a������)?>썝�Mp�&R(�/abO?r��3��M�F[�`G6Ý���t�Hd��ۈ�n�_�S�C�W��N�c�V�������"�߻(��O������(�ܹo|�[�6�oS����7&w�M���Kz�������~/�)2�K��z�a�k�m���{}����ֶ�\��傜F�q[�x�&����9҉�eS�F���C�K�����$�������N�ە��~r�_AT�y��%�7�f��m����&K��qe�ɗNZc�~�� @���+���9�ہz����j�Z��튲�}��4榺��D���n� K�o�{O����Hs�"��0ʹ�4��k6#ﳩ2~v�$�466Wx�vO"�x4���roɪ�2kIw��7{3����6I�6I`�	�"�d�q�i�>n�|���i\KD��r#��-z�+�M�	���Г�7���"�A�d�2j
U�~(�_��m�ݿ�wPg 5畐�����pĻ&0 �[���6�)O�Fn�������z�=,�A�4mļ^��A;0djm}Ǜw��"�\�ͨ�1��c�N����?���W^�L`D`N�!"TImlmb�@h1uh��&.����{,��:bu^c�`os��?���a�ח�{��lx�eeZ��b\b��hz\*�:�\�S�OX/�N�b|v;�p�Л��i���`j~+�[\��9Qm3RHOp�fzHM�`kFo�?3�t\H���c�׉,zI^�\	�Q��"^��c\��X�Y�d��J�E��F�6��"����s�4��Ԥ�ɔy�oݸ���|x���̹�>*�w�p� T}�0�~�o��G�1�(��b0��	vt�Okg7I`S�Y<z
��,��]��y���J<��L��7�G��r�(�N=�4������nk9��T��<k�2�Q���4M����c�Sx*O\k �tӴw����	�|��G��|������8���!vj/�=z�@��m�fb���zx�����
xqe	'<��3���7p��E{���n��^G�@z+64_�nUm�=e��m�ݺ���l��>�I̋'W>Z�S^�+���2v�wdbV&m($QԄ.h�@�ίZ0 9BQMynZ�8<���5����>��|�x���nF!��]�A�6����8�H��#��(m�~	�{�1�����J�^�uo5��Q=�Ҵ���:�"�r�}�u���c[d�#��Y�v��|qۚ@�(�_y�<g{�4��|Q�#��H�X�m�ʗ~]��:�K#Z��.b��{|��D���+X2�P#j��ŀNa��+�y3�؞��u�Q��T�pƓvz8����������m{����$ѢG$<��4TaN6�LhdqZ��C	:1��V�'�):(Z�g�!�"Z�{�.׫��e�q���H� d�����-2�T�2��+�W	�f1u�,��l������M=N��͖��U:U`ҨW��31��x�׮��_}	�1�]<>i��G@��B��X�Q��qD�ѣqz:�����v����ßV��w����R8W��������xc�	BZ��v՚NLr� ln��P4]�)�>�t��A�iJNM�D�IT���<�0k��g�p�_��]�_��M��e2�����.�w�3����G����Q/���Ic2�&��r�{V��-�;y95ak�wG��X,���t!�*n/��]�n�ݔY;t�r�g`�5$�[�f���G
��I�<uM� �~τ�����^*��b�SG���@� ��a�Y3���?m���]LY�.{4Z"#.����3q�b@�A����r���j`aL m�ғg�����g)�鈯0�t��u7VP�XjT1��a��D�Y�R����N�d�/��x�����D�~�8��G�_GsuٸDS�)+D��>$�=�u�)N��/}�^���-��BlY:�O|�|������������7tm%�0�;4�SN��ѣ�����hlMJ6����4�;�]��?�Gwf�#GL���v�|�6mL��e��T7	����������GbnK�:N񱩺����i�D��5��*9���jb�f�b�`��_���;o^��vT
���6@��LbemӼ���|�J/~�ǖ�ɋ�T�D���}�Ә�x��͡���K�'	���� I�C/X?�72|�3��`{��mn�6y4l�&�������E�N?��M)^~�]��Z[E��w��	<�?���x�G�`ueӞ��%��PYA>���S�E`�=�F�Ԓ>/qeu�z�SY�PLCB:rao��=,�np],��I��W6X��F��>��cH�<��߽��b������zC��>��g��#��K?»�\6"|�뙢�:��Ĺt	��D����92_=����/5�771���%���+W��_�9L�M!n��6����=�[z;�!��o���~�\�y^��mո~|vWV��w��C�J�璚eT��/.Bf���ʪ*yUL&3�{k�+��{?�s0�m��w�qO���,mMɎ�ƹ'���v��o��8�዆-t�$�7܏�0��I?����c�Y� ٣�"Z��<l<�aD�$���A�Z���q�Ј&�E�6��5`�	��m���>���$Ů`������3��^�y��P��Y��!4�XTR��(���9�����*�h�|�<�VJ?$�
eLA�MCb���3�]7i3lؓ���r��*w7�}D��w[�X��G�8�����i0p�*u�i�c��L��X��	����g�c1��SO�ݨ�}���qY��&����*�C���w��v��E�7��[��}v�0L�p�|s��#U��rń��Zc\�FG�7�6%T�A�����TF��e+5G���[x��7�vp�����wz����nc��v=w��O�g����1�k���o���_���1�#>�E�"������� �T}m[L�tR3�@�#%�^q�Ep��S�����N@:ze�tOƏ�)&�Q_"�K�ϡ�5����<���>�r<k����ѽz���9���P���#����?�A��"`�4kǂx���h��L��r����.a���鈆F"�L�=��fZC���!>��J�:�d&a�-�ST�M���AISC<KY+;>H�3�-t��U:D�>Ig��Z�a���<��O�<�p3xuF���_���e:�;#qa�  Μ[%���h�V[�Iͺ�NTV�pQ��@���+)Û��Y~ԕ�]��F"��7d E;Fc�����V���Sx�@/Ȗ�>��^��w���������ӿ�;͊5��,)���ɩI=q�R��_���,�����Z����U�T>��/�S_���?��H�F�zn���3�p�m����a�,oce�6n_��n���>�����'�vk���z�u��WQ�Kv���E�"��9C�z
�\�{��n�i$�1�;w?�������ױ-�l�����:��M����8G������E[�oo#�@+W�������+�_6=�/i��gb�gc��a<��#x�K���_#h��!/����M�Ġ���������l��gq����e�^�ǰ�C��,#<�$��䓘{�,rm^����U4+8�GQ�;t����3_�"��?�����D�x|�{�ӸU��O_��P,���^�x�&'�>�>��=�������A)��kx��8\Lcb�^���bj� x�	t����uI�u��)�g&	�*����5��J/�qݠ�g��:} ��:�DT�K�991�G���#G���#�������w�v.����b�k}$]�>��+�*��\�n��d� b�,���Ńgѝ~ÞY�{��d:o�7�� �w��&�����O�x�k_E��W���:z��ux�=�g��Ǎw����2�V�1�v�9h�������%C�����2=M�들a�FBD�}>ξ�4Z#�
�F���S`����r��9�,�e�T��������ߧc��Z��!tU�%V�rڲa�0��?iqRN^-bu�������<��:��yQ/�ѩ�=�ZE�*�4��?4>^U�x	�Ud��8J�^g<+ՋWo��'��FD�j+������o�BL͞I�8�VI:��������&��iX���I�$5!� ���d�̑j��kT���ȱ�T��RZC ]��0J�wm��q�(� }���9G�="Ds��=�u𘼓vF<~�f� �z�,���#����L��e��ĵ�1��t���'�V'��O�e�5tn����E�(S��*"W�f$����A��̖�H��,O#�H��f
W^�Əw R���wAM��U��������2#?�44kU[7ExՍ-��=��pMX_���"�j�(���w����t~�� �}_�}����^�8Js=y��^�_.<Wb��mI���K�m���Xw�]�D�5���o����#*q�N�I6:�\��;	3�M��ȹ��D�����˄M(�=Hw��cR��˺Ab.�1��Q`Ri�_�2�Oz�����WI���c{�?�$Dڦ��x�Lǳc�LQ@$�"S�����IR��G~�����5�,p�r(�[g���ӳƹ���Ș����"V��/|W��u�@�j�k�I�>��s���>m��`P+��vm�R��np_���ow6Q�;��x��cĘ45:�a�mݾ�MQ�8��6�}c�ϫ䛳���h�H�iP�	-�<�����ֆ�����U÷�^�?g�<��]�Q�I�[����w�Ʃ�a��gB�6��G��~wk�H�'�<�)���W�����?�s|�S���ӧ��������b�'@Q�>�X	J�cǎ����~�@��^()&3�=��o۝�|�ĩ�7��,��o���cg{���#���=����~�S�B�s��?�'�mec	�+��[�o�Џ�"p����"���X7f�=v� �4}�Q�V��Jp�șG���!�������?�u�n'@�5 �\�3!��_��_Źg���P�|kۛ�J�k��_D�*����k_S`k����O�^��[W�Cq���Ǐ��1^<Q�֍;u�y����4f����a���^\y�]ܺ~S3�VJ_�q�<�׹�y������߳l���=�{~�A���F�� �ݻ+�q=_x��ӯ�~����el�Ҹ����]c��&���������E"�[6M�7�w4QZ(�Ѧoh�d9�5��U��w� ���ᆀ��22|����N�l���^y���6n^z�x S�)�?"�!�V۬��?�ڃ�R�2
��➯�ܽ���Qy��},LLctx��?_xmU�j-�&8,���F����k�%g�澈7;8�x�wڸ��;��hmW���^�(�.�p���r�@�:��,�O"�GJ6)��JdL�A�t��8������ʔ%5���$�+�ʧ	�#�E/bk5���,��
"�*T����N���U���$�>�T����q���$�Y�Q�e�q��w�`G���K�ы�0�Z��a5��ke��g��NI�1TX�:�zu��Rj�pH�xC*>�aݕ�55�esf�+��R��/)�	;�LI��P�.Jz�"Ե~:�t�?����!#wI�d`�.��D?�hWL�!��x��D<��J8&&��R��nX����13=PM��	*�f�}W37O6��jP�2'�٘���v�RR��E�~�W��%��@ʽ���4�ЍxW���G�6�]�g?VĈ�9�&~�'�f��w��T,ك� ]�R<=���B/]f��3G�m��&�Kۑ�-�*X��+�O��� 5\���^!�n�-Z`�C5�hdC�e���-�8}�:���kwpR ��[c�!�&�ћ;�6�2�>Q��^�9����t�kr�8b�"}=�G�mx����̒$���4Y��9끺��$����ɱb�ں�����QuT*�v�]kE%ј#2�Gq_�꽰G8r�1*_Õ�XD����z���m8�,K(���Ѿi�1K�d�4�˞����R�$��t��#�h9n8��v�D��T����ZW���_ε�U�z ǃ��v���{&�f�[�Ҫ*OD���8v{����{��ӕU�w�I����e��X��\Q]:������&9��*���׺H�� �lJ�L��n�+
$�64J�R:�d�D9�7�����s3x��w��ǫ<��l�aP`�Be;�q3fi��dj��Eū��Qi+3�c���iɬ(Hh����5�V*6V4��$�LK�/����S�ֻ���V��3�޼j*7��#�7�]| 7��E+]�ج3��٥�:|vG� 333�)�:},�{�ߺ�g��+��>���o��_�}��s��ĹE|�3ET�;��ŉȥҘNܪ ?=;B�O��/���m��o�W�x����Bh�K���b��2v�l+����x��y�����N��~�����SHM�crq�fo�w��Aa2�O�{m����:�>bܘ��1�Eӭ���@��	����������D�P�+��|��GX���O���W��y����" �}���p`~�1Z<��|	�._12��̄M�*��y)/�:�J�x�O��{,g�n�����&���[[<����A)����!<�|}�P�~�S���������/~˔"�ޡ����~Ӓ�b��ŧ��i���9�z{��Z�7�s\|�P<�W����Sؼ�d��O]$�M�0M�h�k����G�ި�俆gʅ2Ξ?���~6���rw�(k4�2}|��b&k�0�]4�\P�����8B�;� i�]�����Jz-��m�>p��?BU�=�v��]��v�C��	���W��2�1Q��ԃ)�9�[&���/NϘm>��U"nD�j�H��KBmj�1�����ꦜ٥�~��g�9�U"�-
�gy��(;wY4_��]���Lg�V�S�S��i\d�G�~���1ADJKʦŜ���j�R�T�d��
��E�M�-?���&�G���/�%L�-D�@��3�����L*3i>�*�q�&JYWY���l^&�ڡbN�a���]������\F�C>ς�u������v�|��F	c��	�e���qO�O���a��#95e����V-b�t�F���O
ˮV�h'pRV\�]$.G: %*M��q
".E�������y��˅�h5�����#�g�#��&Jn\))�08+�/ML8l�|�8k�=��?J�x91�D׬H�.�ҹ��ݽ�DPJ�DNK��H'�A�����ԛu�6�p-j�LYdiD��9�'�	|'ܴ���3�1��a�#���$7:�-�@�]M��f�7x�[\�����6�Xߩbcc#�����eXa�Т!������+��|�X� �����!�C��2�DE�X^=t���&ۋ�����zI]j��/�s\ѐѨ��6�n9N�����~�{]���5,�,��}?k�Gh�>�t��C���ȷ�q����ad�\�1v�@���K>��a,���C��+ZBc1{oX�`Ci����o�p7��$̆��k�-p��O������Y��FY��9Z�=��>G�ZI����m��4���Z�ɭ�xK"4p3uC}��|��Gl�Q響h�(�Q�8����o6v0AG��)i��*U;�ʂdrY\#�Ӹ��x� �S�yM�3�j����Jm��-`��lY/� �գ����w��cO�̉�v6���5��kg�j��\Μ� �kڿ�gk�J�,fP'0�5L�����amu��=���B� I�f��d%�&�S�A����f����C�g�NBZ��~hA��ֆ���$�4��>�<N��+:����sGp�+�f����fm?`@�5��N=@RV=i	7{�7B8�n:���*.�?�K��v��j�jNF����c�����Z��z��k~�(�#sX�v;������ɃG1�u�ec��U��4�юI�OO���ɨ���^h�H\��TL������yi�����"�J��Q�<y�14�Ms�z^:�*mm_��jl�?��o��[�&�H�=�<?�v:"���;?[��֖M��;?@j���ӳ8]�7��Fk^mG��	�~m��A� ,��d�`!�(�x��:��O�� E��-��A�`� s:�b�7�)����^ `}����+��j�R���:��4�ss�>z��/�ڵ˸�*�ҳ��l��n������G��Ҍ� ��6
���=$j	��j3�u��Cb��<�j�������W�M������<r��/<���[\���1<�䬵)�[�s�P��]뺆aTyW��eӤˤ�Ab8��b��mp*P��F���v1tɠ������
��*�~��n�d-��E�J��E/�dg�^h�ǹ��ȗM�B�̓A����Z�����Y��e�\Do�":0�ą���j��^�=q������D'�=��)^���7G^����TD�f�Q�tvKHr|��S��F�=s��~��Cz�q� ���Ư�zk�p�D�.��b �s N�JE�~����t�)Gu�.��-�H������	k������������"=\�<��.`]�9�}�eI�ᇮ����@]�����K$'��hd��;ds�!Y��i� ��x۸}eF���b�#F�x1��I�cT�6e��N��N����G.>�R�&l��|5gY�C��l�����Xk�p}�i2Wx��_E�ױ�^�`��.�-yG���j;>D����|��PhG5*s�5I<��� �'l1�NlZs<��E��q,L��=N5�jOH ^�MZ�(�nǕg����J����,����h��>�:�wM�P�����U]��tl"�ʭ�O�W�9�6�l�^������,[������rn,Zc�Z-�H�׀����h��+	�ڐ���T���t���A1����$���	D$)���k��_�\v5�àaM�|��~"=�`��K��x���'U���2�C�~i��j�hAuM�:��m􇮇���c�����V�D+�������}���6dG���m�6��M�s��4�/���7�m�1��� ���Ǌ�\U������ŋLL�U*y~���*[Uӌ�����l��AJ.�Qh5X��2�i�*����˳�E���,b*�A��#���|��8����M'�x���ۣ���[�K��z��ꑓL��brV^�/����_8��b�\�Π��|(��^����.@��Ti��2t�"����|a��c}c�u�x[:ȧNA�W�7m�G��v�m�̧P�8�I�mon�)�3x�^}�-l({���K��Ze�x)�5j���	htz]��E:ҩ��G�����ոSTJ���Xh/1�����:�|&e�[��q��@L�QD�q�G5��{~8�'�*�찏o_� ��,�<�j7����y(�_ʕ,�����;;���nh�6}��͛x������9k?8*08е���{��dI��ӌ�T��.yI�I߸�`K��`Ka��%:�]������oa���ѕ�P>�&����ڱ�9R�p��"	W��M��M;VٮF�g��SJ�����x��W��?�n��m��?rY�!��k/��a�I��;��R %��,AP*�Ա[p�9���Q���x�*z.1��o��Q����[D��)Y�/L�;���Yj���a}ae� ��A���[�_���(iԨ����!��hn���$���-�2�]}p��,����.���4�����V�I �A������ڋ�E��D�H��I�.	�8�� 爄�y�9��#q.)p�:j�9���U7&R�M�PX(�nv���W�Y��{W�z�l�%���l�o`��Q����5z6Z�M&�:�_'2*QqS7��n���u��eS��\��18v���&J�g4F��(�`(.��	R�Q���]G�S�؝Б�Sz0���{�NY#iBxC�Y�7��)=��1��5���o��=ll�,���5\�"���x������Pj*�1� s���d_D� �5����$���S62�����!���Ч���m�s��ЪU��v��R4r�H��2o����e㲦[�p� E�	���1����pr.}>�z���p��m䀝5��7Xa=u�뿲�Iqy���"��޹�ea�&
�0Æ�+-Y6m,�$ݛ���̳ˆY�ep?ȋ��ꍇm��,���{�O"�ʽA��Vȷ�@�/�a�{������2Ѷ��=��h�7#�V�u脼։����~_�uc���(xVY|�R9����Z�t�VUiP[�1"�����GWn�ҁ�K��p����o��w��\y�Z�?�e�3�N�p{��K/�I�,i���V��^r,a"@j"c��,*[��T�&��������ѵGW�Yh��{Nem<5=a��?XY1~*�m���g:�3�({��e�\�jk�ipʨ#����������zb��9���;�c�Ģz�C�� ��x��x����]@J�м������z������JpOБ>t�y�a+�}���k Hd�ڤ�ݝ?�_8t�����m�|�kW��/�M�-����f� ��j�9]�9~}��ƹ�c8���$|co��@� 1�eL�K����E�&��6�\,��?�CR������o��	|3�2z&K%{�w$s'἞���M�5��j��oZ>B ���zw��Wq��%�|  �@㴻&q0��ɸT��q�i�"���D�4�c��
�LN�\.�COl��	���B'�7�_H������ɡ��">�T��#�<��@�e���%$��m���v²6 ������C�5=�Ȏ(�M��g��k�J2:�
\z�ŘN��V�<}�z��ow��y�
����9L^<�Օ��ϥ��e$:VV�x�*	�m��� ,�}��Yݬak���������>w����}�ǖ�Ϣd������K��ĸ�bȤ$�V�Ld���2y6�s�X�Jvm��������?�:���'�6s�
�tAV��g`�Y���ҏi��-�"����eR4?��b?Q�u7�X�{�͏���ZVo��S�q�gFYA�(����U�4������]g�|"%/WarYQ���:����:�Ͷ%����}��S�u�z2oc��{@���q3����C��'%��1��HH��_��lָc�F�W4w��ɞ��X4�s���-��1>'T���Eld�_�}����ۨ,����5`k9�=����h�ɉﮢ�������.��-���BM��<�C�?�s�vs|C��&��:�f{e~��S��(�P�*t�qB���~Mh �ke����=t=*�����,x�~�wK���P�vtj�(�<,�I���K'��ךƣ�D�1�Ky������$�]�&,+��<\Y�F� wce�4��V�ʥ:��r����(�)�Q8ޜ�d:n�����˭��`��M���_6���c� �ŷ�����%�o��&�Vg�E!M݄��(`(��t:=��AL��Eg`S���rƽh AR A�5N�^xt?=�����%��ǉ=�nÁ<������9P�F�mPC��k����K��Y�\���Aԯ�(��}���v;�ݽ�l�o�j�}��A����g�U����J���s�n �ёe)�B�+'D`Q�)j�@�m������h�{1$�h�x����|o��NJ�J��~��Y�%@m�g�F5c ����x	����9���+_#"��ٲLiN`�ڡ1/��a��֓6kH�1����<5�@g��ז���!%�w��d��f}N�n)�0�*��4��� �f?���Z{�Ԃ��9��MɞG=�*��e4�!/�M.�4�j��"%���YS\�֎��%b�$�M�]�9I��S�©E;s�v%��6~����[H�Kx�����%��|n� �t.k��l��Qx����k��Wl/�tF�E�����x-V2���X�"2�vw��7���R���Ӵu�%��.k,��k������=� (�����L#u�����˴���P���#� U�����4�r�$�N� ��$G��C�J0&~���^`�'�>Ī�=K$�3���tn`��Aw`�ZU������
�}K���jz��- �l�'耓�&	��0-���-�Y:�Do�|��W��6��D�H��=�4;������	�GgݪQ�`3u����ĸ&��*��x�.=��W?y@ۙ?|�Z����'��|3����-�9�K�D"c��w�h�
Y�,׳mlf7�l��liNj 9�_k7�c8U0�V�����l�2���*��X�n�Tom��k���gZ�e�M�9�Z�G�Gޫ����Bd�㮬k�n��E`� �#յ�Eu#�{� ��D��g\����K��$�n 3�����NMbnn�l���$XkV�[�?��C��ڬV,��rv���s^�c�[v����Y�ou�;2G���8����x���[e�=^_��["t�j�S�Cz�N۴����}��)�cQ�-@~o&/��Pu��$�JO~l�,We(&bNk֍3�w�H&���2&����R-Q�Z4#g�i�s<��ڹg��i�a�:��쬽�`�m>�����<J�)�>|�l�"ӌL޽�._��i���/¯�����;��ƛ��ؖ�m'����:��|������+���
�C�y�}����f�a�%�
��4z8��$�m�!ٔ0�w^g�$MI�_k�K}3	ˬ8������c�l@ƭ���u�iQ��&s����>͝*�U�6L��9����v�#I��\�dU6֚�^]A���D�Z��.}T�)����q��>��qVH/�����d�E%[�yMU&-�������+Q��ϡ{8��F�R/#A��.���Z��j�`Y�E�W s?p���=��_��A���a4�d �Ͻ�����X����w9*��k������<|����1���6*�$� ��}���{jؽm�,H����=ϽI��K9&�vm'q+{�y>y萁�o������KܑA���~��_8t'ʮ]cl�G�<�Ly��1g�\�������BN�=_�� ����E��ҹjE��(�dֽ6|�$)S���G&g08z/�ޡc�#IД��0}S��y:t����2K��D�N������M��>)�@����(�wCS�H�H������f��Q+�=�Au���J;
��=��*/�w~�T.��z�ղ9O�N"8y߹{o7ū�G���{�w�&�������L�+����᷾�<mK�{�SA�%���o �YkZ�q>~	�6��^6Sj
hb�����6E9�v]�CY���Ѡǻ!��k�|.�y^S��.�E���z��`t=�t�z�ڍ�BS�s#���T�`�*��V�v�םRP�YˏU�0UO$!����y�N��Z�T��Ԝ�)���e��g{t�)^e�VU��L�Jo����r����Y���1�Z��$�#�9�q��ْ���{Af�6gG�F�R��ċ��9h����iJ���XEBM�2�{x����L����6�3U���˸����W��NC�_SO�ZJ$Ԋ���i�G1�Lh.���W����6��w��O�'M񳋩��ש����QDH�e���?S9X�@�)1�G��d9����<�������|'�	W����X����$�;h\~P�k��٣8}�(�x��JX�y��fi��A~�����=ז���]�k��.ˮ=����e�ۡ2��%��pYJ�^�0znfϽ�E�w�[��)͌Y F�8S�T�&���V��ET0?�ed���}ڜ��>��	>��+0�CW��̊�zf���*
Smٜs�R�h�2t����\�ǋ��?��>�d� �clT���+/��@c�28en������ًX8p�R��)ON K�T<XF����s�q��14[�|<qa����|����==�sc�QĽ���i�0�H{=��j�A�uNF# ��)�[Zc�}�0mw���vo>��J��x�8tn���i�D�,��f'�M���̦�o1�ঔ�zl$靁}/������Z[TW�0���A����![Y7��6ͼ!��"�AA�e�NM�Ꙏ����\�v��8D�%�J�pO��۷�v���}D������ވ�J-&3+�������m�V������(��']yw䦝��JQcЧ�Yd5&��Wp��-K�S���އ�DZ�֘��v���O�Fw6���?���~P�yQd�1x����z>�%�դḻ@�`�A��ȷi�񰄩�(c'�ˤ8�����~�Mp4��������G��M���@�_��~�+6qK�@(�%��|��I\1x��Z��}P�_��{t�[�p��m5:n_�s3�r��s���,ϗ3�
Bգ7�H�N�#M�5��/L4�~�ν��g�tP�>�Q���������v�7��\Y�uj1�R�X%���1�w��r=V��0���kU�|S�P�Q�g�5魲Bu~�@��=���S}�4I{�Nml�Y6:�|�E;Y{x.;�X� �s�Q�<Ck�����9o��L隷h�O/b'����&ztL};{0*M�E�2�r�e�� ����uʷ���:mi��9�\�O��q� ����M�����i��s]5A���c8�O�;���u��Z��\���v�t��|F#�����jq=	W%j�OI3|����9�L���p����)��1R���ԣ�	u~H`�	{����X�M�˽���K�(�7�Dc�}G,�e<��Öe���)i�Y�nm_�lac����A/i����gJ�:��*"cS��s`<���l.��%C������9�(������ٰ�ID�E|�#'�&�u��w^��Kj�����CeF��0A�j��AM��B��,e�X ��h8�%��V�J�w�e���/Ugszz�Ϝ��#�m��XH�P���ॡ2{��5��7vyF���'=�WV�����t�D���9^:�N6JN�]�)�$�AED%=<t��뗀[x�:y�$>��3X�$H����w��ӄ_F�gObz!��'�Lr�c��qs/��|��o�&�dI�L��;h.]�s�@i���XD�ќ��}/��0�U6:U��ٳ�o{���e�/b�����S�!v�?}����,���ak�L�g�2y1Ӟ�-x��ˠ��~j\?j�JU��Y ��\FV��g}��jX���U"��.��p��1<��S8s��5wi$� þ�v;�܀M�;qG�-��[o�nZ�S���֯� �p��G�eg���Ec��G�<7�hm}'6�YS�&���z�&�Ƌe��� h��&Je'E�+j4ZF������d��FX�s&f���HN/D�kl)��/Q�J��Q�zŹ:�)sރ�F]Ek� ��)�	+�E����Y��T�R^{Y��gg{a��h=\{�j/��7Ɗ$�_{-�k��>�TR�OO��H���keY���ݳ�G$�g��Ȉ�c:rtD��)��9\3E��x"����qf�C/���3y�ϟ|�T��#��Z��Y����C?�Ơ4��*�?o�26�x��?��4	�}���zƬ�\g#�����S�;b���|X�gQ�h2�=.F��<��+�ƭk�v���ш�<Y��q��g����;+hT�tSH.Fef
?��>hV�uڦ��l\���z�Q_�(v����*c�&�J���"�ިGX�2I=]+C>���}�!,�|��5�N��ѓX�9ټs�N��$m�&w+���K32�/ӎ��݀T2n{5�\?����Ǫ V�Z&FT^Q&UIО���$��Ж�O�u� rj����&�Xno��o�yݚ�qbqw�>��Dz�l�đ:�y�|{��~�@[ר���Ý�	<� �s�����M� V��M9X;A��Bs)�\���)����|vA覮��-b�g�u|���Ʊ4~�� �~_��fx`�k5>� N���V��l��SEy"�zC	64=���]kV�q2��|	��~6�.��Ov	�ڦ�S�G�U�^�}St���U����Z�}:Nu�+�/��E6ۂj%�V.H֮�w�(�a��:A�"V�45�X��6e��!@N`4��Z��o�;�ң$�Q�9��e�-��H=,�ٻX)T��D�(Xt�4�(9QD�o�S:��wF-4�G[ݮ~j7p<m=�0�ux������ꏰ|k��e�����T����y�:Kj��bp�>���l��]Ȼ����{�~�aۭf���ꍛX� @򿶄����Ӈ��؛Z�4X�1Hфh_�S��\&��T�h�����؝�m����xĸ�3�WF
o��O�@1A�����w��y�:.\8�/|�S[�q�nmo��T+���Tir�*x��$���<��	��Ub�;/����^5�Ӥ�
b��g�/aa�)�8�[������2�4�6�dMʕ���w�/4��,�Zl���s���'M?��Ƒ�Wu���g���m�S�� E����*� 5w�AF	�,2>�^�"i:mϏ�k����BW�&�Q4>��87���:+�P��'@�������~�yLq��w{��5T��j�GJ�}�j���l��I�چ>�*��l����/��*Ns�P���.*d�'�z��*���~ޥM}>������GFFx��iƑ��̔��>#����S�U"��4��zĆ\#��ۤ����'F��Sw�)�a�8t�١êw�!����|�~V�Ng~�<�|�Amc���sY�����M�4��@ԑ��+I�:o�͚�������[�Q66��="z�i�:�]}?"��Trp�S����9mF?�ި�{˽���D�)�9ei����.���z�54�v,S'���l7�v���T8�w�Ε�ԤiL��({"���T<'Sݫ��/a�3��&ieĦ��f�252�*��_v���� �y�4�`�������k_���ƥsg�J��Rz��0F2l���*�`��5h�CF���!��:=����~R�;����t��M�֌�d@5/ ���S���Ii:��(ѿ7�����o\}��̀��혆�'��y�	̶���٬WV�O�0u�����{�Iv^Wb�U�U]�9�tO�� �"H�	�`R�Z�W+RZK�-}��my�L���+-EK��$.A�  �� �<�3�q:Vu�}��_�4@j�M�7�鮪������{���8�'�/�dz%��x�Ϗj����CQ����4�4�ej�3˲$��r�3�D:��+���A$�ľ�}��Xp�q��a�Jt@>��U�|��&�&��؊��2��F���V	���f,cG�DG�=����]}�������[WE�����Y�̀�c薅������Ӳ���C����IP�TT����k���,�m8�5'�񶫉}��(*���;u�xVyO-������/��t�G��jf�����õc��N�/^�Zu������$�ƍ���P;��@���!+6,S* y>�`X@� �B&� Ue*Ď;���WJ�Db�}H^��v���j��3�V.�ħ�,��u��8������5k���n��KS�����7��׋������ԃ�+�u�C�Gl�a��8�+������Hf�p%�;2��� ���?�72��8��K��c�E�tN�'��05aወ?���&���d_��e,5�������.�F����]D�Q��{�kWR�������Nt'�=%`�4z�mm�d_{��Gh��L8ر�ٴ>�<�r�ٱm�,�:�I�H��_!��MG�,�W��ro��z�����w��SO /�"DQnN��8I��n��r���:Ά����a����\Ք�K^>3����g����ubque�SAl�؁���ۂ��xx]Z��:z�ZI���ak%�d����M�q�4�:���W�[�����..{X\ki�m�0^v��H��4{Q^���#Gq�M{�s:LYւ�e��' �T^�y�N	L���s��Y]�*'�{��~�w`5_�-]���*�ky��1�o�z�,��8B�yU��k��.]�Z�=�+����ʥ��1`^}CNj�5�>沪��WC�Pl��l�7;���t�k#fu$�6[?7���6�!X>S>W�4%0��t��*.��%��T�<��|�y/rPd1��H,G�<�+Ө^zE@WX��x�]���C{uF������5� ���)��d���*'����^4*�1���L��g��આ��9�c�l;�q�֚l��$��e�¬��%w��gS����4m��H�3����[��%�:t�T�\]@㏨
;�U	��!��t��"��.�I`W�:qzC/í�a���@l�l�D"�b���tc��c��߮�-��!̡�T�X���~i�IkZv�AW����_���ݻ����!�b�:����)�⍄�ّ�SSR�W��E}�	q~��PΕ�1���	�Jb�'�yX�6Y��G�Y��N]�9���nWl�.U3�g�t��ݨ[�)xm47��G�X퍬��c������+��VW���"@�1�FI����B�XuG�����v��W2}�Gpf|-���*[v���t��*vNHCJ����S�'�t�ޝ�5=<K�r�!�����?�pO�	y�Μ��V	ã;���ǌ�ޏWp�ZF-Q���i�� K�;�,��i�!h'S�E���b�-�K�rp�¸���#���=��q��f ��)�TH#. 2荫(4��z�'(	@|��Y�_[��_�{l����;j�X�NqzbCh}rMq�M����:>%a�z��V� '�`�^��zFg/69�܇���Djuo��|��]x}uo�u%<N�_���`���Y�e:���ؾ1�9;VVp��9�IY��>8v>�˿���nEI[����:�_��(�˿��=!@ׯ�*���?�~���_@��8r��q����N�z_��?D����6e9���}����[�۵��{�LF�Y��ɿ�:�}�Q�_8�I��gG�$��<��]�stG�ǭn«?xO|�����ܿm'�~�����1w��|�,����гw��K/��X��}ٻ���X������[�V3�Wֳ�B���wA1�~��Yjf�I?"� >yv��i��3��Y>#^O�YS1kĘ��&N�=�~>����o�TY��(���%p��z�Loy7��`���f>:�~�dI�R��0MV侫�e�d#�g�P���n��Z�:
�x�,������wh�J6WT�(�O���)�6U���ڨ����i^ ;���өN�Ex��[O�16گ������_Ä�f�l�l��F�h��v�+��ݲ����fv���7�y�{$e�Ro�:���6��ffřTq�Y%�E�͚p�D��D=!$V�;�IQ��EO$d�d�f�sX9`�G�ş)3t=�L!�ˡ�}�q�B!t2*9S�����=�t�b����L`@�����t�D!��f&Z���j.L�7��B����VG�������r�6}����n��.���굴��s)�:vI��3�m:[J�v�]FJ��.�w����n�u&�e�]mR�&:��okg��|X[�q�C�G:�����Ɔ��b����"�q���}��Q1�f�^�k."~��e,�%�0"����9�f���nF������ظa��qV�r��N�e�F���"NdܸJUIE�ME�EZ�rxYFѬ��r�#��'P�7�k��#r1JFt�!�ې�_�(ћr�"A�$�V��Y>��C����*PY[�J,*`8"�E�qC�E��LBjze���p���FU�}�]�c�D ���q��Yz�M��X[���}d��D�9T�ο�����ItC��0jne�b0{{00؋t��:R��y�kٚ=i�2F�sI��L����t��d;nӘa�EK��v�,��|���.�Y>7������yM����E�m@�mfj��Zcr����6	��D�i���ں��w:oؖoyo6o�po~*�:�w��K��/�]�:�l~� ��=�"� �V�&�~��-�����NƥѹӀoq
#�>�Q�V�4��w����R������_GQ�g�7l�*$`�	8�����䍤8�D8�K���I , �X1M�e����3�>��R$��U���C��v�q��8# &�O�uf
w��p�w_�r�Ky{� �!��X)���t�&��K���X�LN���#1��8�h�O�ETlI@�I]Τ�JP�74� ҥ���ﾁ�#�Ctr+�=	�ݶG��B������zǇ�e�$v��}��x��ӈad�V�t�vNN�}w߁��(��*�t��;1�����o�C����{�ͦ�G^�
�L�
�o�W1�u;��?��geA�N�s����n\�:�?$&�K�Q�\Pn�j.���yy9����/���?� �l'*Q��K�iI����/#/뱘Z���,.�s\�<o���]QΊ�u�>�F�Ω˸p��H�X�M�m(`��Ӯ#� �9����$X��pez	oΞ�3.�5=��>����5�Z�ד&[���dN�V�P�Pl��v���m����2����[�@P �Ubύ���ξҔ=R� u*���X�gp�)7�@��m��l��_�AH�@H&<8��+��$�eʎ_�YjU:�!{;&���QlJ�Kw[7���q3T�3:Ї���:a�{�T��z_�
m��N���U�]��f�5���U)�e��d���G�r�իS��`��ɋ����@׸��+�d���8oǅ2��4�a2������[��F����.����E*(M���Jnm��4#�sb�[0�D]�b=�*o[î-��{U�̴{b��UA�gx�##*����B�rhC�
@9�r��:w��uV��l y�S����C(�;�|߹b��� ��U�A��2c��]�����uS�C�ݲ-�Bj�f^���;������R7jۖ[��ٵ|�-{vm�K�mP���f�f�b5���{����Uh�,T���f��k�9�63NA�^?#�H��� ��.�(,�+�CG�#�F���'�C��6�� \l떍�t/��Ė�$�T�zm�*�fft�얭�H�z�^N��$�x�n�%v]�9�Q�x�>�Bڋ�S�i�y+WڀY��t�dVNm`:���,���]F�W1�F���!�\'��m�W7��~pfd�D��h�B���]z����4;�Zb�!?|rX����\B4(����-� 26lZ�
iR<�ڔ��ȶm�K�d����(�2�KJ���U7�c��B��Z�FsFw��6�sΠ�G�)�(J����c�`T^P����5���L��! �ii~NgS�,�vh�;﫮&�7����h��f�6����@Y*4�� ym��E��X�۰эt�_�W3oo�*a>��;ۦ��`�;�F����p�^�}]�z?���\�I���h��{������̟����}�g�٥(�Nv�]e �����/Z�9c�n
)�6����\-䑈� �3�¶?�>�+�i��H�a����` U��ণ7��q<��+(�K�!2�+���R���5������q~vN3 5�60˒H��T-����(JD�`ߎ����O��i�,Fb!��?��O���`�`E?y�RY�u$���E�J���L�w�%�Oe��u��O0�ϔ����O;�#ˌ�勨���q☼>���_��#X9q+"����}㈥P,��_�>�zƶ�w�#��Ϗ|�<���z��I��Y�,
�*.?�~���8q��رcB�8��%<���#��$�_^P�G^����WA�=�vߴ�������S�����
	��$��;߃�/��L��+o��_}�[p-�
 �E=�E8@hxsKKx���p����[�c�n�;u
�~�����9<���f�~��O�BA������'u؟�ٟ��g��vY���-�3XZX¿���F��?�-�r�V�]�ţ�5	 +��SQf����ǳ��f��`�|�F!�������c� �U@��+����(\�����f�Iu�2]^�t5�?�� W�+�����3r�l$c�j�
��NiP�E>�R\����jД)��bC��j�*&��,�&0�ۇ��ߨǺ{�^���fJ��C�V���Q�p$dʰ�$v�����M�d�&�T	#���j��"O6���P@3`L��
�۵{�$X)7�-b]|�[=�ٵ�>�]u�Z���Mg1�&uN�{���6gbK�V/�,J�ޖ`�b�p�Ů�6IШ 1�l�ё5��m�8�wRl���7�y<����[�+1د"��hRG�~�,�r}5�嵴-+i\�����I���	8v�g$�\��=�*.N�MU9˭b���w@9�Z�R	+�r/��A=��N��<�RL�C���F��t�VC�(��$�\���xu��Xt��>�vK��;U����r]tt��ew;c��芕�f�ӽ�F�?��D�Nm�Ȯ�>�)��T��� 3�"�<���&(��4KnxRU�!|3ܝ#�q�G�܃{w�q����whH�Y}����O��ߋ����Ϡ=��a�z��$�Um�L��l��+���kV��T�j�a�̴�C3�mE��rq=%�T[�0\�!�*ǉ��Z�u���#08dXΖ�FZm�N�o���]m�L[F����,�D��NXcEC��9H�����GRm�+�T����M�{G]ڱʑi���6�n��ck�ul��z=�S�&���d��c\lh`��f`�020Y���t�X�tk�ES#���A4�AO�34�r��2r`yi�����:�Y��|�����b��n9��2�Yn���R#����m|肧\[��`j��23�{w�,�z�n~p��n��V�.���{b�������f�L殡� ם��]����J���n�F�ksv���7�*6i���I���4 �߻�T� v)���J�hj%���E�Q-8�Ji����gq1��f��.���iGj*�`����Z7��)J�����Q���@$�e�����L3)�w1	l�	KY-��  �,[))/���\�"�	P(���0�D,�rz�%�y�9�ݧ��:"�E�u$�t���y�1T�~V�G����[w�DU�eEC���r�{�.�ęz��:\��� )���	`ddL3(��.�O����߆[o�YA���".�����P�i��E]@|C�^�ø 7N���_I�#+�&>1����R�c�����ǟ����l\K:��x/_��)	�h�7?���>����#{��KO��'�@�$ξ�A8<���5�v���q|�o9�����W���
Cs�*�+��糺8������{���8�cw�$goO~�lqS�ĖT�&��<���}�3p�3����O���|�v��j��g𝓵8~�M��C��d�b<�ݯcim	[BbBb�[e,_?��-<�;?��(���8���}�	�c\�dt���S���>�셢ؓӯ��sO|�JCr�(5��j���f�
���erp� R��/���74=Z�$'�����%���pV,��޻�\
$��U�� ����g-��xM(�~R�uP����E��j:�]焗�LR�dOP(Y}X�%������Pk)7{a)�h��jlT��/���������k��7�Iw�<H��ė�o[˦�Vd�Yx3��R[[U��N�4'�9b�m��ee�s6I�x�|�,�Ҹ4� O�K���knf(��9Z�l���d8�Q�Y-(��-��]K����=V������et��j���ݡݱ-���B�C>M~4�9x\L��?��Q��#.�R/�S��Ȟb����@}?	��
�a�z	g�N��Ki?B�U������c�ǰm�_%r
ՌN~�%��=��m�|R��aYq��fs9L�K��o�ҴrŻ�;�F��&Ӓ ��҆W�6�Tf��Z��϶�j�7X6�<n�����xw����i[v��$��Ta�R�(�ѥ�)!j�z�kÉ`�Tk0\!ِ���5	�g����� n>qG���3��&��
��37�b(�_EU��B>+�'���~�9nF�S�)�9O�7��11Č��X��`�P�]G-}����Q�T��'q���vH�$��ѐ�@"��N�`Ư���bG'*�����ju�F̟�e�v�4����D�>��N���@���W�De�rc�����ق�� Լѡr)�y�[qt쾥���vz�RN��_A1�I�Cn� ��8�Ȇ��?4��m7Q8:��.��2ٽ�\�9\ؤ����`�eF�mp�6��WF�fQ��2�-���g5W�ϧ^��Ҫ��'F�1$�.�]C6�Q�˥.s�,+J�a���l���r�K:��u3~]0�1�o�M�e�LĻ��=`�n�
t�6�4�I�x�٩"[#:~ifO˸?{}���w��5/���:v��>��S��2C�R�,0��-����1�%R�������{�w�)F̭�0e�LNǦ�m��6r,f�@A��j4��zdI=#?�i�d/��l�fѦD��ĲbP+5���WQy�5D�}z4{���q-�4'���!�O^΀rj�>�ine�%ٷM�檖5������(�l{L�S�߿o|;�D���@Q��{`^���8���V\�����-سsw؏��͢���{p�Λ����xgu>	4}rF���9q;Zl$;�6����~��V��D	������=7�08MF%�ZGN �+�S[B�2f��Q&�`��Yl�FQ�ϡ�n��2���R�6J�"}�N�5�`�,:�ѣ�?����LL�U9W�Hc<3�D~�ЖIT�sj�)���$��T9�n?z{�(����L+���yt�����f����|6�l>��PD�jJeD�z�}��K�*�T�SK�E��x��G�1#���u`Vo��<�k�Ȭ'�'�uϮ��66����f��{���M^�X)�p�,ܲ����cw(,k��@�<*�8����ߌd����W)��Z�Z��^��
���y,	(�����
(��}HH�08<*`"���\y�,�W$)��Ŏ�Qۘ���eʌ1��q|�ßDGl�5��'ߐ���=�NoR]�Y����)޲��� �ӏ	��Y	�a=�ڼB��W8�Q?F83ۥ}.�fR\m>&&<�5\p73�Ě"===��`iY9f]
+cc��-5�.�gm����())̈- �9�+��U=X\���Ip�[3��V��CK:%ZZ�u�)1�ƙ�@Dp���V����}��:=#�7�ײ"g��/��������,���%�i��ˋ�v���F���q�^��?�_:����J��UҦ�v+dw�z�m�u������HP-��i(�50��6�R'���;ovi4ժ�;x��k�kꂼ�anr���Ȉ���\Sf�և7���߱	�݆��|�S�()�˩Ζ&UL>�UX�+.�l��Btp;�S���'����tސK�	$�T�� �
�[���E��pЯm��<���N7�?���������I�`|�V�]=�jvA"�ڂ�ٵiF�p�f֎٘ںl�%94)d��C���]�j��v�5j*�l���e�	��&�P��4F����B�2L�#�&�l[U���j��E��i�[:S��a7�9I�:N-��3ITr9�Hr#x�~5���D?��
w;;��B��kaf�9U&ƥ��U����V�T�^N��ɢ�ȡ-C<����vf:PQ�Y�M��J"40�!���3��]���naq���v�`L�ף!����-�Đ�[J`.Q��e��.���&�v�w�d�U�U�e�΍�YK�G�7l��-��k��t�6�72���������"��lg���9K�:o�3�[��@���>�ͥ�.�t��|�
���[�3U������7��(���F�g�:t�9�{/9O��Xu�Ŋ[��mxݿw	|W/9z�_�}�d�nhf���AGq��]�U��l� 8g�2�e���@4�� �� ��m;�ƩӪ���q����r��O� �3 ��P#�?g���t�:���/~J�k�@�")�zՒ�`����:�rޭJC�c��론n�W���h���\
[GGp�s�޽�p��Wq��<�/<���th��x�����L����N]Fjib}�18ِ���3W�7�W��6�R��F��:���h8g�V,fe�q�"F�zqR��|59�M97��uU��,�U�#�I`~��wu�A]���K���}h��LϬ"��tę8����~�G���D![ Ч�Ƶ���l
5�	�ɕ�4u�~�{��3=;#�XJ�i�|�=�
��U
��q�%���3�[[� ��ID��%����gyl�s���S8�֔v�^gܖ�$�{mi��˲�WY���εi|����ܵ��v.���>�c(Cj�L�� ����DÚ�U���;0�������0z`���(����RM�E ����T�?}��~]�,~���µ��Pd����Y�m�6Z�n�Mn�=��s�s���,�����C
��z���O���:���~�>�|�ߒ}qI����w'�~��ַC]<:w���|�SS@̍HB|���Ml�'�a�)�p��e� �K�w��W�S(��0|dr���asF	�,cW�t2��m�Vײ4��K��|�Ďz��'%�D�򫭢Cuى�ߑ ��r�t���,�&�,sމ'���T)@�J��B:��s"J�窂_gc�������.{&,'���j�vL���_ g؏��[$�s"]�#�V@)SՁ
r� C:�f���w`x�_��V�b�(�����Lt����o���˯�B>���$ϡ��X]-�v����8����=A�G����A[M� �<��M�o��췅�h��^��Z�au�6�^�+�Ff�貴�\��=�nvr�]�ͶiC׋0��~��6j��94]���3m���|�% ���#. ��87q�"��j���dQ ���:�m�����ʈ��1<:�z1'Ѽc[&��[�p��1�{1s�����"ሊ5��y5����*\A��5�nJ����NM huF�ނ Ĭ�F��;ܘ�
��� �U/�~���*��K����j����2ህO����=��FZ^YA4���j��x��*JD��6Ё��K	�ë���|��Cg����������fJD=�f6�v2�~Ղ��[��MٴZ]��l�e.��+��=C�,[1����:��q�]s��\JX��� ���3���z�nۆ@8���i905��\�.+v�Hz($Qṽ�>/IN-�Q��J��`G���Vw��F	�fx���(� ��ݶ������0Mٞ<�M�t.�2h�K&ƍN��C��k���rx`8~�s�Rͨg�_�$ޘ�a��\:���ٖni��]���HT�}�~q".m ��!�_dٰ���݄��fvT#�\KP���L�s�k
[���Ы�,��z��k�3y_:��rE���0��BH�,k��ܧ��&P�.:8��UU�'�'���OAr�j�8U���Jf/+ٜZ�@z��(��(ׇeO�n��9L�,��dJUw�E�}V�s)�AKUU�\.��z	���s��X�����ؾon?�+o��+6���w��X��Zy�����f�_y���Y4�iD�嗖����Cp�_'4��͉��E@]E�W�R�W ���Y���*YN�9\������y�"��#�\�QW�L[��׏����ٵ%��YNs<��򪨧�p]33�q�����{`?��/ama�n��%����c߲+��-����/cnqY9NW�Laiq�n��x�Hj���,ݣ�Ϟǵ�%-ASQ������η��j(�hLi9�N���ً	И ��U[	GQf镁���+��9�C��FV@�p.�8�J��(�1��c��]:��ҫo`���o�߇�c��迶����������0u�z�Y�(}% -KJ�� �?��SXYZ��rHZU�Q.� ik��t���i<��H|�^8q|�����?�)d/}�������q˵�|�?�r"�%��R��o��~�װm�|����_{����|�Ch�q;�I�a��Й�G� _�������&���x�7��f~q^y�B��?�4�X�G�B���F�8�<��	�-!�=*�<�J�����!���5��Ւ��u�qy&	D��58�^�h*�Ō�c2DeN����3�k�TP�B����f0�	�dj�r$��\O	9Y�t���t�����F����x��y��5M�D�a�޹K��6���X�#�d�U�'���4'�̒J�y��	��ϒ��5jq��b���S?\e���WާG|Z�C�1'��~��I�`��j��a�x�օ��rr��& �
�%8��VG4� �-�Cj����e|�K��`����5��~!)�x"�(�rh��%1��f�7��ZN���J�t��D>(/��F�);��F�P�x��<է�����:�f����3b�>��E�S�&'�����=�J��y#X�Pc�{�vY
G6�?�/��5�Z�Ƿ���,�(3y����8jv���a@�|2�v)���{��Q<�;&�(/���f�Y�)8�)�c��G��Ѩ�N��q�L6����.�vW3ΞM�{�=�t�Y�UY,��3�!-���A�p�Cpu�q���
�4����F1/k�U��_�d^5�:��|�jQ XAn[63c����Cf>����	0a��?�C@�l�.�c���a[da�T4�ۈ-���R��c�أ<�.����@��Lc���ԑw�X�$��@{�u�Ԛ%�0C$�El��L�N��� W�cQ�жm[����1�\��^ɔUIf�� �����-wV��L��1��U�d�Ƀ���#�	#P
����]�?){t_[G�5Tؒ#��.����l�<�d�a�++yc�u[B�c�Qk(q����F*���@�t��zv�>9A�Q��\-h�9@�v�U�@�w�f�^&W�}i�JP���T�h���m$zڪ[e2wa9�*= ϰRk���'-}�5%;3|�DJQ�z�w����Jۣ>�p0L]4��Cp�R5�l�]6P��2¸$
G�%�g�%�*�^����A�,���N���k.[�ҫ+,v� ���Y0�n;Jє�%�>v�}.��*�@��Q-C�J�8��D�:7��2b��S��)�f�=��i��4�^X��_�����ⴊLIm����K�$ϹZ���9l�)?/��
�}�O���o��:�K���`�ݼٝrף1����EG@������?�54��@��<�����%�����˯�){�"A�U�h���x:kUv�˙�y�IJm��Hd6==W����M
��7^&[@E�{hrB���e$����c1���g�RՔ��Y���
�s�&g�!{)���"�Ba����+�Y���`,A �LcZl��� 2�Il�@9���5�J�������'�M�"^��z��̴�S�pQ�Җ��`4 gȇ���C}h�H%���J�$@PΥ� ����Q�s ��o *gۿ�G?w�̒l�j����ZkI�~I0ݾ���"7=��+b������e�8E�C~�����s�-&��@`�ӇR�2��àc��o$0n�:�\]:�9����z	}�8�_	M��$�zꇸ�#�����;�q�H�8*o�ыP���m���ҏ=������F5��obf��=�{�%��Љ���_�5��Y���feͲ*��r��T9�Ai>���e׋v���\�B���=8o� V�x����8����^,|_(�x�:*�:|�#�׽�i%�X/d`�:y�TC�*Ӥ"�7޲����}��*nM�-�x�Zz�5;=�Kʪ^���C��;P�?�B����
�+|Ȋ�p3S�`߭7k6����w�G�1���T*��oLcmmE}��`Y�}Oă��(���ީ�-.{ٱ>�S�av.iD��NQ̓8��C�owQ�	������Q�/����S�r�{�9�}��aY-S�_d�U<[�P���G5f0�Isy��^�Q�U�3���=��{��'��r���M�(�v�6w�����s�����a�.� w/o���BZ�T%`��8�� �N�{��(64���&��ufui�ѐv�Q��W108�-c[Q-�U85�Q>��D��h%@�tM�qV�V��;%W$�e�SZE�mv�aAy(�H
) �i���"S���Ʃ��n���TM��iF����f:�͜'K@D�*>�}E²�9|䆇������� U�/i�"j�u��`����&_S���E����,bY œ�e��\M,,.!$���F���A֡ߛg�j?��de6��ٳvyA����I]#��5�\F�v�R��7��N��?ׇ���� ���8\F�m9T����ǁݣ��Vt�h��Rb����A1�-�F��	K�9�A�ΐ@��� tM[�˗S!�i{S}"N��I&[�[n*���������d�.NGG���c&�^2���r9�,L&q�eF����}K���ك�����S.��'Wb;�s�:/dnA"�r\�:�����8dո��M��uV�v�r2�X0���T��ҹ2-`���̺EZFo��$��,������9� �	%��`w��b���^���ct*��O��5�{9��s�W�R��YJI0�r����Z����py��W^�^'�٫�c�	�1]�r[''�s�G?~JGO���������z��XֽQ��Ț�tX<�Y���SW�
�p�	.bqSԸ8:��S�2�S��T"
��=�GR'_ǀ�������������>�+������:#Ю���7KN��S����,{fl˸؂<JEb��;&������_C�(k���cq._@Y�kp���ݦ��-#�RI̜�BTքAw�za`�u!�|go;��և�JRm=��KWQ��L5�\Eٛ���c瞝��}�|��W��_���(�\�,~���G�������=�:
��3�@@@� �*� G ){�6���=��SwF��K�����I��';�B��@�wL��j��Qe+�I�91Ci�\WjB�c�^��Z0[����� �X�O�ΐ��
�+���Ѯ��j���8m�9wuJ����P$�`�rW5�(�oE��!5<�驫�������Mt�MbD�y���&1��D�G��� ʋkhع�jۭ/��xy�U�o�u���(UF|�_��Gc�B�-�t(���@�). �<{���0��.$d��gֱ�`�D���-gk��6ݭ�&G���8Gi�oF��>�Nr�5�d�e|	u���޵�3��'k=
ٌ�.b��i���?���w �@B~/aHלo��D�U]r6���QYf���`֯V�%`j��-�	�k�jj
�%�y�w#.��M��g������������#ܘ]���g	�H������>}��]���,�#��Yk9����us?�9ه�7GJ��ƥrx�.C�h��)R�T�������5�uh���d}��E�2o�|��_�5S����&�k˅s�ST9FmGv�%����=�ycѹ]A��('ϱ��gY���{n�ݨa�L
7l��w���m�,4�\���v���\�謁 �P�j9����etj'�F�ݲ�1�HA�3�O!��R�0�Q����z6�� ��J�(�g��S��sx=+G��.���gIHTZZN���>nzQ�r3��z���{�����C˞��(>L�%J����JA�� ���"���J�7b���=����M�� S\@����1�ޏ|��`"�Pz�t}��u��]-��լ�fn�֢�`��8�cD	R��Ӣ*:LFQ�u��rv�Y�LdU6nN,D���e&%4�Td]�-���w���2X��P0�T�ꊉ��>�1s;F|��'Qaj��rV �)��P;� Y"����ܚuS7uB���ev��6eU�ҩe�u��϶���S�v���1��L4A][���0�v�����弱$�@�M�aK��8�T4rj��P��P����Qɔ�䛝�Z2�TqT��Eb�������q�O7K�Ee��[�ƣ\���/��^�XU�.��*���>$B�;f�C�L�=�,��]�v0,{c���}�,R���`!�qP�`�q~o7?�?�5?�o����j�%��s�jV���s\]YCD��#أ�+�ELD)x��AMێݎl���%1LV7�{�Y���%�H�=K�C������ƸK�.�@x��[ey`F9�2��t��x��Y^����h$�W�,��ͮ��y	�'q��q��+��k�`W_ @��n�����K(��^�:�-{b��c���<�w��ȑ�HD��R��s���'�$�zN����n��^�c��]9��_��Ҋ����yyr�r��M�Љ��鉫��！h�G�S�'qX-[����<罇�C���\����˘&�k�"�sw��Xo#/����!=vT�L_���^{]���>�Yq���~��}VΑ��ƫ��D%��g:Վ�:�3�ܳ�?����"�B���>�e��Y棽�}C{���8~�m*9ŀ��g^A�҂q&+�՚��
�>t����T�!���o��:~�RĘ��%�Ͼch�����	�@{E�]c~j��3�tT1#�)p	(���4���@)ԋ�_9�[dM+��M��x4��|�6��,#u�,�DN3����5޲���_�����p��?��?~F�Y�J���~�۵N��PX��| ��s�K�Q	w0�s+��J+��QN��m��΢M'�T�� ��6��3s�\sW��4�5o��m�X��/����i���X�m��r�����7�o�8m��o%vl�&�%i$��c��؉Z�2��jϜ�6,��A4|�ϼc�[����2u��޵>1��ʋ�|�Y������$x���mj=��뾾>����G����\�;�eXul߹�5�N�x��E$�I�Id�<�hL_��l�ߣu �6ҏQ{W�]����t���+*Ap��T+9�+N�rJ�k�|ڠf�b	�SWw�)�ɋ͛��{y�U�AZa��U�C�eo��e�7'��yd�&��1���-vK�qr̋iX��~�W�HF�̜4����t� 4(�t���,Y*u�#1�e�U����"�,�O�~���$r���}Q7��={�I�c}uM�oM+���aR��іd9� �(f
�|��*�Z�N����B�L���L��g�e2`]^A����t��K����Ё8	��T��Z���+��-���bGRS�!����M�g��r(#ޠ7�����
��#R���&_ţQ8Y�B�v�K�]��vؒ1m#	cv�ݠ`�{�����Zjۙ<nn�T���&�U%ZqZMՠh{0���"y4Z������+N���p5t"�P" �xL������D�9p HR�I��Ȑ$�
���BeMX6f���fڹe�!��_ʸh��){U�:X�PЖ7��ʆ�dɕ��x�v��ED���L�ې��e��r��ڔ����B�MN�Z�3�+���R��\��#��L��<)_՞�J�xY�D�CÃr�h���m
P��3XXX�,b�Ұ��M���2To� �et�T��t�d����|%�串V�d�� 0Qij���O�n�P��6��YF{�$�-��N�:Zr�2'��>Ћk��R�(�ڸz�
X�A�&�*�0[�>q���2c#����%�݂�>�T�9�2�#�9�A�����z�WЃF��!S��z;H�^�d�����e�x�UW��Y���:094���C��מyO?�4�(�ȷ��kJ�a����sx���x��:��;��zP5��?y
�-����n{ࣸob��p������Na]E�����~l�>|��Ϣ�2F�����_
ъS*Ukz���}r�;�.�xӑzNg�͠#{���ch�������z�*+s��	9v\����$Ӕ$�����k�^)0�+@>"p�M��c�=�*�kw��ɗc�a)i�G'w�����_"�~���^��m�3,�5��9,ۅe�:x��SBDf��r��hY	�x>�����`�\����_�_�j6���p]W�d5�߆d��p� n��N�On�@)���$��U	,"��P��Ob��8���p�F0v�	4�Y�߿����/�	a`b�	s���k/��<�ځ�������_�gp���h�Ǳ�w!#Ϫ���=F�9~;UU�W�0j��x,*���L���w��bf�<򵯡-6$�� �o�QF�k,A��g��`����"�>'���v�V2/��4�Q��J�R#jڽ�
8�"m�V��FѬc8ʔL���Օl������-l�]��}z	��l�il�lٶWE���~�k�iv�2^�!��wH�Ƙ�,��j��p�r���xGda�nv�n���S8<���E��$��ᮻoš�����Q�����0��7�}u�S_�w�=�^���%��A����r��M�P��V9C�f�4�u�|�|:k�y�X����3�1Ħ����Ѩ3 �����MU��B��%���s�J�.�/x�Aw�	'����� �JR�ˡJ���0��F�Cn�����͌!q���P�~; �NE����9x���ж�_��x��/t�+����h�������F(��襯w@Z�G۞sW��C<g����%������7��(w|xA��23閖�kk4Ǔ��Z��Q7\�['R��	6�0ت�0+�2�E���v��e�L�6J�N�_���NN`��72�N{S+�c���Х���^�UY��s��SE��rm�.���#�1�`�j(�F"r��k"���(fy,KU�[�G0.����)Y�Y�x�>��o���z	9�Kbl*j�vY�mY���ZFĒ���-���Aۻ
0�igOM�;H�J����k����f��Z��k�"�r�4'�al��>�./��D0��� v�E�m��Q'�ñk�\Y�r�e1�5%������?���F��zG3He��8�;�,�@"�k�Y���qq���rUC�R��0�$�mr�6��}wj��ɓ:�zpdP)\/�kX�����c����!�9�3��K j����a\���k=w��t�$A�[�u�,�P*�Ӄ=�L�9�J����0v�ة����~�� �)Y�6B̧q\�؞�ӯt����̎8������qS�[@O��z8"�jo�	_�(`�����`�:Ԗ� ����t�6��(N��
�~ێބ� ���|SW�~�\YM��s7>��/`m|i�'-59�O��	<�7�->�e;z�Y��v�'cᅯ>��SS��Ϭ� ��-Ϥ`�*XQ[Ay�ΎԪ�3�S�%FKS�Дg�?À��3���Z�~�3�������a]H����Ȟ�#���M6r��: ����pڎ+�\G��N���B��Ob~5�G})q�#�8����A��Ν��L���9i��`��y��'^8�*�.�a�o�=�1-�Td_�8~��=ңg�Ru+��ʩ�H���%�B��ٜ:ƫ�ty��LQΪ��'ܯc�PZ��U��d�n�ړr�9�h��!9Q�bD���琖s�,gEl4M�rg2Y)�/���t
Z[�Ј���֦��S�W(�cU���䈼�2$����r�����r�����T. �L��+�R�w�s`�e3�r�b�9m�͋�p��7>K��<>$`޿����G���*����{�	Yym��5�ɕ6��va5��X�>� ��u[wO�z��Nȇ_�W����=�8r��z���x�<oV��)g�gW��w��s1(�`��v���Jj�T!vW�zT|�7�"{Ѝ쳯ʺ�Q�����!AQH�@��TN��mgM�ب���*�JN��N߶ڜ�	�*gt}�9���a�n����ҷ~ޗv��#P�&3��f�py��2EV���č���ɫk0���#����첬YG�Z�dTl:1�K��U��V�s�sx1w=�WN��m;�_�E6�T^��e栏o�І���o�T�jP���r)�Go�Y|m	шOy|1&MdS[��n��
JM�y��?�h�w��CNr�>���t�&�g[�	�Q�1�oʜQ7�\2 ���9�^y!��y�U7��ƨ�cL�CZ���pY�!�ײXpm��o<�v�XM�&�nɶ)sutV�]��nJ�6��,i����m��n��A����WW���{���i~��Ѯ�\v�kI�މ��֖�5���ʧ�6��;�ˁ#u}U7�Dc9��f���r�ʬ  �?�'׵��\/���*'a��?8b�H,���h��昢A��[Qn$��.	`0���H��3c����	�2�ܨ��mF�m{�(������W��u1&�|]�;����It'�&�]gS��r�Dh�Q`���C��֜v;�ƣU=�V����
�.#t�m�,Q"	�W`M��E-K#L��,[�*LG�����g�9;�{TEHd��ai��E��Iu�\Of=��8��%[�WF�z�0؟"�nG=�Ge��r���b�ӥ�i"E1* ��#�4���[�A����Ʉ<�9bؓN�?y���l"f��$���>˛��K��nF�s8xI@ bO|P�j�T
1��j\e��X��y��_*U�HnݺMŕ�U�Th��8��ۇ'�����-#Z�9 ��CB�ޘ_@�O���a��$��=k�S�4�� p 7[e9МY9&�m�U�щa).	>(`�;�E�#�@ɯ�C�x�A���82�{+�Q|Qw^���^Cmpp4�p�@\��A	&��T伡g_��t��n�67/���R�p���>|�~u��3�^GMݱ�ߏ�Ǐ�~�	�>zۿ�E��:��W�����<<2��맱��v���Fd-����������m��>��x�rVG,2���FvF�eK99m�=��L%�܈!���ޣ�Xq�߽[&���?�%xB���s�Z�h|��s���q�Z��G��M|��_�/�����-�Q9ٟa|�׿ �&�K'�_|�Ő������[��j&���WQhִ���&1�Ӌ��������Pƛo��@��
��(��T���qe����
��r�"�g07?�DB΀lV��ג�;T���ǟ@&+`U��s�(G�aTQ���A�xX�F3��y��~%��S?BR�Ҏm;���`v��Yu����+�7������7��P�y�c8�M���3�{�{�GF>3,��u��='1I����ٸ�
�RJl�_��W�⫯I��9��$y��s�m3��\?V��/���K�����<�S�."�7�,3�p"^���!�+�0�ݨ�^9�[�����xZ���/����E��˕2�}�����s�����&��
��M���Gz��5�c'����Ƽؠ����ؐ��SKBb'�%�O��N��ױ��U|�W�1�"{k�Kb������~��M��~���������.D|a���3�h	PgC�4���D�*���ͪ���n9�sC����^]Ѯ>h��:����rLl,��Ym
@�K�6T�*b�P��	��h����.�I��%��CM>�ռ�Lk�?y�l����;Jm����8���'V׫�^�;q��U��)	�waU�˥�z�e?�>�:=��v�15u��~�sD̇BN��s���\P�,
P۱������4��j`O�P�V�7&�<ʳ���Yf��σ�FS�M�ikmMiCe��Z)*��5���#_�3A��x4�䂧��u���DHP�ӕЖj���l�{?�S��X]Ko���-=����c��ڌ뮬��Ch+��x�Z�T>�<d��k׮���]��0%�c��қ�Ţ��{�p��L8<<���hx���<�|}A�����Vj�SČ]�P�����ؘ!T׌����U���ր�](�\(e����������I�0�İ�pǌ����i�f����-JQI�8):pI�ٛo_ ��ի����.���s�#�t�2���s�T��Y,٘^���h�y}��値� >�>�ey��9���G����dX9ftL��!�mC6gs��VpÀ���"�~.G[�G�eR9ttF�J��>R�/˒���ȡOV�L�����i�+�9)d*��c���#�òRi���ܴ%��D�<q.��ҬW`�~zZ ��҆�q�<��ր����-�uWT;TD��-�����C>2���[��Ss�/��^&`A�w
EF����_T���&p���*n�L�n��О=���QX��F��#	M�o�:�R�D�=��eK�K҅��W��[�v�����D�<�B�6�qL^ģ>E*� �*�(����N��!	�un)��[W#~qt��r�N��l�,c�B7�b��Ʈ�U�1��3�2j�g=�A��e$
�)r�a���rm�*��MN��Q��`����p����8�_�u4�����+ز}/�������'O��Y���������܇��p��b�ŀ��6�篼��wߎ��������������hs�,��nr���M{б�k�Iw��Zp4��"���{q��	<�� q9����G�}��R83��;��*�vr/8���e��~��x��Gp����?�Y��������/�k�u��Y��f�f�06��z�~|�#��/��ϱ|�ܭ�F��0���¹�����	����%	|�����[\�gQ���{�}?}��(JFJB>/	�P���3_P�D9*_��7�ď�B&�E�sGsFd��.{�Qm#܎�!窹���o���s=~�^^Z2��\���5�	0<��;Z���Y�T��a��Eui͚�՟��O�̋���8ĝ@�"�tl��}���Vg��c�i��,������1���v�ו�:Ý�7x f Ap�(RM���v[�[�ǲ�vwG)Ǖ��I���J��q�;q,��Ғ\�(Y�HQ)��<�o��<�sN��߹ %ک��K=x�=�;߷���Z�U�r��|��T�������jĞ�b�j�Cb$����`0�؍�KKX|�M\:s{{M�ӗ�fl߶NK씬����p�]Ƒ/~�t��:6�� ���?�z�����/�y)��BQ{>;Q��r�^C�?�����F���M���`hϴ��+x�ěx����~�A���i|�3���m
����`����*"�El��>8��rw�؁ꫯ���+�*�h�j!�,�,"6��+��d}c���@\�����'v�\��L�'�8�z}9˛�`ㇽa�ߩG� �-�5�:��(�]��]3��=���'t��++��DX�%W)�\b��iaR�H��Z++%	�Gq�<ߋ�jY����M�=\p�J̘`�A�����<�t�\0��˧Ω�������`���J��8�%X�G'���'`L#����[}ф�qK޶�A��9ז	��c5�r	r��(��Q����O��);K�� �0su������f��4�I��HBTS@N[˕}��NH+�^/����E��w�Ę4�5�-Zf��g��w�ұ����,͓�_��09>���(�:uW���`~P)`J�T|�N��3ʤe1�wG�I,/TqQ"N�)�'� ��,Ȝ�+,@�=NCfद��QY��'�p�	q�)Gh�B"[�L��\	(UX�}#	x!O��0&�4�Q����GPH�	�-��-��+����e-W�P�3�E��N����n,�w��g�jT<K>ŵ%$Y6ȣ&����$WRd�#��[�p.	z}#�bk6��=�-q��߂��!;>�����8 ��p�\�������o�`6��Y9��^D	��H�: _�IH�\Q*��nm3l&.��bm0�����X%�n���,��c!\���:�-N&'��h�2,/��,ה�f��]�c�&?���m[w
�ۤ����#yt��\�9�p�S�)�\޳uw�ىmۦ�%���cH�g�k�aO^���)��y80E�%�������T�2��e�?���\WI�Q�1���`0#�Y[ YЬ�^��:>8��Dtlvwű6�9DZ �$���]$b�8�:v���u�EO�53
�Y�TB�O쾛_�ay��N3���
Jծ���HmG�W�]R,}V�SG�E[�[:��x��� �]/�����}��8t�x�ٯ�~��ۚM\���M���Cu��'��\�	ٯ���� 9ϓr��
	�+E<w�"����[�bp�ڲS���7Y����I��� g���~X�*��|�I<��O��[��D���SO"?�e�vM@��Y��k��X~O��#q��{K �	_y�iD�2���o0������}��ǿ�;���x�����g�g�*6��_ӧU��M�b�Z����]1�v��%�>RK�N����Fy��^�\�LZ�T�X��)BRDR9�X��-f�e�����YaX��Ѡ�<|	�pydq�h���l6�ޓڒB&�&׀��H�cm��=]0"�[J�m��o>J����l�6�?'�
�ʛ�V�!����)@���m6�R�wi�ȧHIƮ�2�)�Ttڣ���I��S�Jp��A��rz�W��2a�Z����;0�e+~�7~�wm�q�(����~�!l��n|<��X,�����y;7M��מ���i�ɱ��O}
)�+�v���'?��W����q�F����dM^�<��M���/����A�y�L�������ru�����_� :��]<
������L�������I��9���o`��1����(���Z�;4��0�A9�d������-�z�g�gd��x#����|����3u��Y �cd���F��:��=CA���}By�ve^�����	L8Q}Ji\��BWU{�P\�Q	(��E����B5��F��f�C_�����'���a�)P��ϟ3�'bs����b��ZUܸ��t&#g3)��\�#@9KI�@1f�\��!E�Cp��nJ�M\\'Vr�^@N'�m�
ȉ��5���'v��*�جJ�6�S����ǳ-���k�w�5&Q�:�
B��TURJ��Q�a���i���M��lu���ԯ�.#��c���������{Ӳ��� �.��W�F���p��u�~�<�k'�d�صko�uNˮ)w�8B��Tڈ���٫:X�m�6,�ސ�9�c9|�X������z��+���9�:�������F�j�rS����٦,x/%Ni�tc�U��׏�nE�,�����l�"G-U;��0;U�쬁��3�̞u��""�fI�Η��]�d31*V�_�E�u��A�����Sə��5	:��(�K�nR6DzA.���F���-8+�x�2��#��n6�=-���x���CQ��E���_>��qY��LO�%F*�y3Fz ��[P��LKtY��KT}��I\:z�'Oc�Q��؁#9#k��h�"}�3`o@��������|W���%lY����;���1��8ߤ�I�=m�����������7���7��.D198!Nv����"���[Ap��S���.`rr�c���hjޖ��#'g%YǸơ�46E����aF	�sK3x$_�+�㖨�=sH���T\9���D�-O�f�N���RIq�d�;\�W���5�#�y��ς���QZ�O�RQ.����b�l�xxy-A��cʲo��,��B�� �lpo%�i��aIxl(���&R��.5��R��ʒ�.S�{�E\�9Hg$�wISa��>�!S�bGs~��.%����py�}�kCm-����VBY��#=x���%l{���_����g_��jM���3�����g��!���UE��--�&����g��ג{��M3Mm䓔�30��NS,��ȹ��R'63<����P2�we�*�0���N���:���`ғg���}�W�������'�+i�o݇�3�h	�������N	q�����1���U������Ɩ�	�������_�?[Sέj�����Su��J��jW���Em�<�f�4�#�"��g���*�;��(� �{FiF���W{�M�=#mG�̆�(E�X�ӊ�����]*W�1�=�l!'%����E�g��u����=fC�¤ �¢aO��m��~hO;b���Q�M�H��!y8���T8,�� Ƶ�3�D$�)��%8
T9bߣ�!::����� Q�Л���m˳K*POh�W�k�H���?�,���[1$�����Gdx���������hH nի:PU������^	�-'��r9��0V+=��l�܂O������e\�qW��FJ�}:7
Kl .�� `t{��s����Xĥ�}'���j����8����DM�SSz_g��+���&bغe3��K�|�_Z�XB���Zc�)ˬ,X�dڅ�PZ���L ���U�M�F���2�"]�o����-ǋjP�|o:a��>C:f�5��d�	.��[��\���K��IE��@QK�*P툏���C38sm�g��r��%`��������YhR�c[|13��b�X��U�СTV]}q~N�r�lV ��N �K/�0#��8`	t��߼5v@��J�Hr��#[?�UO�E���Q�]�W��$AfD�p!?�)V<Vɺ�ə����͒�9~s`���n,�*%F���u�M������A�ਵ	�o���\��m��h�먃��fxǫE�� �	`|pmV~�M�����g�Î�)|�>�W���ocǎ�'���=�r���d��s� W� �ѧϊq��Xm`�D���$^�z^�)��d��[�������5'V,u��|�Ć�b��:�*Ջ�f<3�ҍ(��	�ӟ@36�s(�%
��ۦi]��R���9����D�Aac��"	F<�=��dT��T�OQ��]3�7�\b�!���*8�S��8UL/˚�6�b|k:���:�t�Дڗf��@��{�(�b�0�Օe4Sb��L�ٱ���mٜC�X�&��r�TiR6���;��w�8�z⃨�����q��+(�X��9���\y�F�B����S`�Kd�dLO��'���b5��+5YL�N�auU��@�1$�N
q�t<%����5�F�W��*F�2�q�������s�%��L��8W�l6cI9P���8��frm�q ��\�N�AJ�ch��e��[Pz���
Z��<s��氫ΰ�5��	�d&�����	lzf"o�[Ufc�?����5�8�Q��gk����TZu�G�8E�s�ֹ�l�pbiX@�۳��uY��������_Y���87�wG �Fwec 9Уq]C�γޑ�I�D��\R�o��!�Z��� K���ݿ�q&�:㱈^��ʼ�g��د���{�7���}So�Ɛ8�*^XY�5Y�nT�L@��sq��q��y,^�,�&��3�����e���q]r��_������Z5�tm��_�ϔj�RMC�h:��M*�D"60O��f�&N����r��8v��y�˪{Kq���S��un���#��w���s|����XYq�i�6��ڲr�:�%!#%�\G{tu2�0KB��b"r�9F��U�K=��:���X_c�n��Bk�f���Ǣ���3m&v��x���Z5Ӗ��s��+�R�� �ֿ���t�Ɨ��t�d����q%X��[N�B�f7�Ew����[��y�ڏ~�C�R�ր��=�Ξ� ;*{gflL���=lj8�59gQ\ ?�e������ F�lǶP�<�����|����*���){g:��7�r���PC�k�Dg�ֆ��"�p��E~��e�ʬ����N���`ȍᡩ}��눋�OI�ؒ�k�M�!��h�+���""�2.g�7�i�]g��_*}�si�o�WzX[�������'~E[9����pe˒��V.i��?��'|g)��g�ş���a�Ƀw'
c���L��enE�Q>��3�`<��˰r��,�ͽk���y���GVΜXh+��ѳ.v��Gpi����*���r��166�Aa�i�f^�Y"N���5KUq�oII�&A^<j�3�g(
P����^�7��<.]bt"�/�dr'2[H�7�v5콳*�������c;C,��c�IAz��a�|����]nj{˾$��dΘ&�<p�u�nջ�,��ei�u[3��6�"����iu��
'yCL��L`�������{�奨�(N"���|��,��!�Z��ma�����}[���T�4v��-`9;���ʕ���Cbp#��؊�ksJ�I��� (n���{�߅#�.��_�ʋ�`ǆ�&QZaZ'�|���(0��uCNG�ђ4�N|�6~h	3�cK�P��Ґ~N C��I��>_ y�T��5b����@h�Ni�]�wu��lTțڱ��6���jS&}G�1"���끎mW[�)Gu�P �U*寮�ڕ%��\Cd�J�Ӎ�аh�G�o�3{J@�N�e����&4���f]�N�B*�H�-0�Z!1"+�j �_��GO*��Gn�>L��rz7ν�:'O��t�иߘi�+h���{�(ѦD��@y0��8�����$�I4P(E�X���	�%��Tu4="F��-��|
�TWI��Q��f0!�p �(w���\٦{�&����F� ֛M�gT�)ό�\�
3�=K���L'h�=�WK�]�&��:�� �}b�8O�ɻ�L-Dri��Z��,�V�F���\ՂT^%�I{�ב�^'�)��ļ��n��Q �CL�N��2p�U(���/[�i�e���5%�&[�������_�I�3�K^+�K�$O{����:�֩	�����1���a�-x��2k�$Uk�����UB�x��e�\[^@p`���_�	,����ӇP8}ZV��벧�q�ޔ�$;��L�28,.����3J8�I�A6@7m7Љ_꽆�zF���<�bl)֑���_�� s�����m��/� �>��%����j�{ͪ�*��VK�
��͞�/=�y|�_����[C��&�;�޲��O��)�s:E�n�&;��7;�`��C"G��li+���N>k�+~MK�l�	k��[��۔�==���o�& S����"��Xi9�d@^� �pp������Ma�O����3�6|��������o(�n�/� �#ߓ��}0���>A%���Cw��K�����N�,�~��h�E�Ȕ|��o|';_W�����IP�e�ʾ�$u�Ym���n��a	\���T���4�.^C�ZR���L��-��4��$>(�S�{���_��3������~�%p��؋߇�����]�a�aj<�{��E��B�K�,~!h��=��k���?�~͠�ɲ<�V��W� ذժW��K_n�>�#���_������ra)T����V��j�g�`Bl�o��oc��}�l�y6Z��v33�e+�`�[|k�9
@����l|�jE*f䰇�6%�w�G�vQi�{N}�I:yzV��V��=��z	�U�fKXY���Z��U��	�k�ܰ�#j#%^4!�=�rPV�zȶ�ˎ�������7��̞;'�gA�M|s|��"?~�J�A�J��J��[{��r5�fT��*��dS��C���/m������m�J���i/� ��C�H��N�p8��(���o�����_���0za��
��}�R{"��.Q
e�R#[��~�ce��! Z R��@�������o�گ�q��H�J1��v��h�L����.h�Z1eY �JMLo�����7��o?���q�b�۱i�#X�Q�eEh��!�c�}c]-�:a������a�!l���K���`��UE�i���4���fn��;���� w���&a4{�����&�V�f�I't�Y"=-�3k�/�c��5�U�>���^�L���h�N�|r,@0
��'��{�";eX�G]�CcrC�>��ScX��e��Ib�~Jƕp��y,��*�L\������ˮN:�%��Ffhp�� �>�aX;w`��O�|�D��*3�e"<�;�L�{hHi�t 14�pt���6bb�,�]��X��� ���(�Mb�Ԩ ��b����'nJW�UBq<�GR"4}��l��Y�T��:HWG�)d5+�ϛ@�1ivr!N�2�F�h2j���-�:m[K��qG 5FH\�U
HΒ�8i���wIj�3`1��L���B��9}�Dؑ�=6j�$▽FI46�>LK�~Pe3�cGf�H.�A"f�8��ev��d!��K��+/R��k˪%���29��{�a��Q>	Ѵf��Z�Jx̞~'O�}O}��_�οu��3>�n���A���vNc���񹧿����?��Ț|��1~�|��pCn0Q�LN��Vʔ����1ո,W״	�N�4:ɡH�q�'��A&K��%#��$��X�k�̟�)�x�>������Cc����3r�=9��!g�Z+#.{Y� Js3X��������Z`P�*mΞ�],�4���lˎ�cg�ґ7�&�I"��m�dF'6m��^���<ߐ�F"���~&3����� �w˿Uw�������`K���f@��7��-�{@�������u��u�y����%��/��.~�}b�)%ҿP0�G$̀k����3N<gگ�L�k4X�k�T"򱸴���Sؿo�������:�ˣ(�&�r>�Cbh֥��v�2�+�X����/��D����SZ���JXX��,UR$ u!�5���kW������� �f.���|�����g��ctz�؃Ry��{�n`5zݴ��ܳ/��E��9c{��#� ��j������33-W!'=G*� ������_�5ꕒ�e�~�Se?�cu�@Ql��}T{����P_[�|C�`��%�W�Tf��q8��9]�|%O�!; TпQ4�V.X%dFx�����񎄔eh������F�׮\)���7�g��ԇ`r8����lʞS�.�$D��H@KY�j00\�t�����O��\P��	�����n�Z�A[��J�,���~�OU�^w�\�GUyG	/h��Z*}���:�J��t=�k�M�6�w��XEطC��/�j:�d���;
�hrR�<�;�N�j�ɍ���?�w�B�T��<�9���ܴ���g��k�MtU�Lq��A왞�ɷ��ŋط� _�~c��&�jC@]وF8��0j�}�0~��7�x�%��������MoCm���֞6-���f-�}�-�*W૳ղ׀e�4��LK:��Q�G�QGo8����v���j%��҅�Dr�(��y��
ذ�J���j��Ⱦј�,���"��2�
d���8	�l٤�6� /ע��vJ6RU��ڃ
�Y����C��S�(�d�x�8�`���{�޵��*�+Hn՞5�w�W�X�<���Y��lۺ[%�%b.���� �;�g�}n*��{� G~����Ls��p�a�D�2�Ѩ/�����r��r�qG�e��(��@��b��\d$�ʦ�����cu�y��c��_R��N�͗�%�zT��,�
�y�κ�OL�'?�vB�/k�P��!�D*������=��ٯl�������)�����}CX��-;R��0ϕO�a�Ĭ5'٫�AC�`��e+<��q�D��Б�$Ha�V'��1�coK�>#omL����o)�'�[M�Je��i�104�@�2���疊x56�����G���?�w���\�ܿ��2`-���^?�]��į��?g4�W_:�-��^�'N��G�΃��bd4��;����=��O<�SG��+k4���YA�VGvӘ �Պ(�	�^AgyAlO��U��`�6C�i�9mokK@C�b".z`�6�1���ZU��o�<����љ_��w�ס���6�4]#͖��3���h��s�i���O��NQ�|盈�C����$
�1 `��{��������q��C���<�3CG��k'�����FVm��}�u����j�f��#@�Q���
6ٙL]�G-�JT�fjt�j;D��xz7�~�׽����Iz}���	�x�!0d�n��tH�d��u�6%�g%0��=�=��z�/����?�u���(L�q�ǟ�{���(��
V$X@I�q�j��@�s�=�A�_]�g>��Q�P�6�6���?��`���+O�X���C�b,��ŷ��|�
"� ?y�vl۶p�U���Vs+3�o�^����ӛ���8����-��\  ��IDAT��f5kn�LwL-������m���4*9ͮ�m��N���b�ka�Y�}���DZlQ�S���C�������⅋���`;�Z���R���X,|�>��}��u�ځ��] @��;��y��N������ �H��	z�����7Xl�����{�=��γo��2�����p�H�M�$�LK
	�[��kD��:n��=X>[�3?8������q�=w ��!#�O�ݑ{��ό	�P"h�X�\���w��M�w7����Ml�=�~$���!�8'�C��˔hM��ψB�_韲��yv4X짔g�)vJ�����ǎj9��䤉s\3PfCX��;^�D���d�Ye�Ӄ8:f�ͮ&:bI"Nx��s�'�͏1k�QT���)`�]@���H�M{M����U D�yq���SX)5�Tj!��öS��5��qٜM�m\�vY���8~���7��728wׇ1���8��n�0(��]�6�:���� U��)ǰ{6���H�e$�c��̝^K'�����1r��hB�Fܐ1�����	q�b�ɴD>L�&�I%�vEY���w:�عY�<fz:�F)fh�r>�xhkf�|��19\�xD��2r@��Ҙr��&=	��w ��h�؁��|Βg8�J�p�_��! �%n�������{�/�Ǯ]�d=+hʵ<x�����o�ıcʪO���ލ�(��p�εA;P�i�oR�:#��t%H�@D*��� 2��웨lz9,I
�H�8��+���1K�C�1&	s�H�-'E{y`fu���1d�̊)Hc$��"nZ��vK��X�e�Kd�i����\��YZg��m-�29)�"�y���8��|� ���V�H��7�=S��X5�8H���x!	*3��������_"S:e���g���ђ8��<��|�*g�X,
ЈkDN�M>��J�+W�?u
��/?�/�(��0�(�f"����uóC���}�س���
r"�ܺ�8���8���`��)l�#�ߣ�p	[CX�[B2��,	�y�Z�^��x?F$�8��KԼ���؍M�z�eԴq?�@��T��������!�Y���È��45��Z:Ն��b���|�����i[������!�
A6���ero��g��XkT����Z��^��xA����Y+"�N��{>w�����n���4=��oJ_7{�֭���6g#H3��fyVm�-�GKH��|?۳���n��W7b�^�3Tx�}��Q����bs=7�n���w#إf��3���z������-�����{�{�a\]����T��59�u�~�c���rX+�p��$�!ޑ@q �f=�
5�����
6܇<��ʋ8:0&�ɒ@=��3H�zN�"m� ,RGy&��m�Bt|/��/|�ۘ�`y��Z	�(c�^���5|�W�������x|�~�v�t���H��
!�}(ɨ�pM��f&�Qq��<��G�˿�	��%KI�m�|�K�]�n.�itN�>i&��FA��W#懜{
�5��3��~/0�^�af����4�c�S��3<���u�f����;[%'m�Q�9��|��V0����Ƒ�>�^>�S���|�5�|�<�'�uS�&.�ߌaeus�%��@tvnsK8w�y�����c�~�.�C;�d�Ǐ�۬��m`��ƛ�m�Ę����}��d'��.	��JiD�5?̞sk���I�=��͵���lxY�͊��̞��f	�J ������y7���^�xroE��F5
�O�)�"��5zk�=�]�����?���>��������Ͻ��^>� ����n�j����YT$��q�2�.˯XPD�Y��:�ql}�Ku�ku}�U�C l�\/��s�����-mJ��Y�nq���&�M"/�DW�c�)\fa�O��>�y ѫ���l�Da�&�\�1p�BG(FO5���!�椩+ �47��5�� N���Xi����l(��/b6A}��[v"I�][�ۑ���kXYZEn2������޷��A$�t�<*�������)٬P��2 E�Y�:snF����Β��)�ϴ|dz<�����XfMʾȥ��z�bb<��D]������q�S�P�D&X��b&�����i&�};�܇�Q�=�TvI�&���!]#eF�a�:��9b@P3��p�<<1�43�u����SN��&5��Fn'fg������:iM<��c�F����l���l$� <���M��:q��*��av�/P�	}w�g�f5�aa���aeW.�����`�Hb,�(�,n.j˭8*�8�ϱA�R#o�oO��"��p��_���1�Ť��䀈��qt���⛟�Sl߹��a��iq�;�0)��;����;��g�S��Dp}���_(��w�	И8�{��/���u��k7Z:�G.5ϳ5���ѱZ���!��RI%/�XȲ��!vF����=1�#��]ZZB����⼀�r�b#Kգ�n2���l:��%e|����jC���L���L1{�@E�QQlTCl��-۴|���
5�-%sU~0f�"=%>�����v`d������������{~��Vgn�_�*��W�v���~�� P�Dz=-�j�]��TP����m�F��c�.�6
(6��
{����k(ͭ��k��^�a��Lm�F���JUl��9�+\]^�3G/��!5N��v%�	)�����!��]��ۿ�� P=���c�X�C~�6�94�������B>�Dr ��8H~�����"N�:��xL���4״c��n+utzh_ys�	t>*��]tʲA���k@��V���"�S�r���$~���x���?i�ɹI~C�H��vBy�]?9������V0�~�5ѽ�%+Z*e�i�6C�b��?�r���2��m4������<Gǐz��˿�O�]�� @��2C,����Lw��;�Q$Y�0^�?����>���X��|�LB@�؜zE�u+�h V�FNȜ<��Ͱ�[43�Nf��$*~�m1�gJ��?ӊ��(�i��q����*bGi�ZHpZX�i˱�a�3u���T��m��G� ��y�B��{Z^�W�����Z����ޣ��<km�7Բ���.�a�Z�[7/DK��:�@�YqĿXG�����G�P.s�dwUt��������Ľ�ڇ_��?BM6���uAګ:8�l��{(K�9�FD�}P���|�{���JG��Xb�{E�FC��_�a���B����zx���C`؟2���4Ξ��$����)Z�8��c��8G��Tv�.�������R]>J�j��Z@z�v	��@��}��c#~\OO֖�q�t��rX�e�l"/Mn��%rvɤ��e������a^�������F�u,�k�:�.���Md��laO!����'p���q��[(��i}p}~^3vQ/-��)H����I�i%?��,R\� 	Sʩ��k������$����=}Μ�����:�F2�#A�>��=�@9���+UB`���=m�cv��3�ʹ&�c
���>�i4����1��S��x��Q)x�'�\�{T�p����O��Y�J�aJ1u�����Ay|�ٓ!�����cOn��v\��� 'jU����ЉY�"3
j�������,��p���F�S�<����ԉ�-U=,P)
�^\)�t���y!�P�b	��}���O>������iq���5k��I�G��?��!�=��8<p� �����G
�_����!�/\�%��9�'�-�p$���ҫ+�D1�2� :s��T�#��>�WV ����xߣ��_R��ڏe�h����b�Fh	���j��Jgmݹ����#c������W�>��ь��Q���\��Վ���Ɠi�|�9 ������i�VU�h��
�d�oW�4����j����]5�:d�}��f^�� ������W�+���g��/�aY��/(�!
�	�6� 0��@�Z�U<b_�m=~�xm��c��@��3���px����RI-9]+��Oh�A�q�ٟ�	%�o�C�I�G��n���cJC�U��I��w(�}߇��`9_���\�Ё��͛0P���,�gfѪQ�tE�")��L߮ �|!���&��n\|�m�NQ� �!T�+Jó���W�8����J���a����O���D���������k�d#A�����c��S��Ȫp�V7�Jt�&��F�J}r��I�8yJ텥��\ð��rQ�E7��s��� 6l	���ąNC����:p�6J|2�b��mi��5��r��h���_�����Y�)jC��`�^�����X�NŚ��TM��7��m+��v���i4r����-c��2P] G�y�\��$������Q��.@q/#>6�j;�6ՙ�P	4r��m�e2�Zb�Z(�Jp�d?����f�*l[�e1	�c���F��#�r-��oK~��D�7_� O3KV��9�@��XY6�7#��f]���L4+�>#�Ql] D���I$�A�����C1>���T�b�j����:-�B��c-:��{>�Vv3������:�vo|o�_yI� l_�uZɭ��̂�J��9i����^����M�ڍ����4�r��ETB���4��1i��`>�8��\C]�̭��^b%���4�B�针�2��j���1_	q���x�mE�����?���7�H����.,�:d�/
 ��zh���Q��3b��I���+�}]irh <��-�w��W�ڗ�v �e��bG�1p̬,�h[�5�lcF��Û�'���b����@N��8A��QӲ���K��4@^i?�@��𲙙ʈH��T{+��%�H�����q��=(�PV��|aP������lG�+G�JrpH�L.�f��Y3�U�lj̒�'�$�m5H*�k(�d�7V,��?�Yw5��黦DlVo30��@�2����v���� *�N!�>�沀t3��5AH�C�p`�	4�������%pT�h&�l���(UŲ
���v}�|#�h�e���S�����Mώ�p}h�K��L�ȭȽ�	p�
�J���qj��$�u�[�����=��V0����p����=��U�7\1��v-�^��K��g�;��1����~lq1	 v��/ร� ����=���Ԫh��y���r[�n��^@Y�,��`�s�z�aك��1m�'1w���؉�Z�x~�	@��G�z
�S�1BG#g���ծ���-ȏ��)�{�������ZX^���W���;�4��1��=?`�Y��siv�˿�C9v_�[NL�W:*Na��Ƙ��J��'�_M�-�0Q��e��>�C�[2k�;�rnC}��^�
�uLi�<�J�L�I��k�&n��Ξ}C�k����~6���G2[�Qz�^8�a��)�2�rBa{~��X/l\'ٯRR�{C�k��8T�=�I���̖�|���jy�7���������_T����1�������K�22����_�!���u1*SC�Z��P��iaei��إ�Mr�Q�o��bc��ȩ��R���V��➶v8r���n��I����\1p�[b�f/_�3��"V�ϭ-j�I�i���V�%Td�gQ/�*
��y�ýe�=I���LBd��zb?YA���t1�A WiH@�Ԥ<����GT���J�O���6�*���1ߔ�Ɋ� �t�����9P�.X*�3��2��1�����t/�nd����ט{�d}�j?�V�A�J�q��wsÓ:F�iV=՞�*�L":���IyϚ�W�Yр=*7��X��	�
c��z# �����[��'N���[�(״[SVMD��8~B����H��u��Jr��L
��Y�3�����'�ͧ���eIR��g���⻖k���(z�k���k_�e�D�S8NȰQ�c��y����z4S��yX�22���ڵ��BQ�MK��+H6D�I!��~ĳ���'�X����%}�RA�F櫻�o���+�۳��+
��[�9'��nVL��tB6���'H���z�Z���z�o��1�o�|�'S�ck@mמi|�d�'��UU���Q]+;�m�9u[�<_^���R�M� U�	>��}��f/��ih�f��d���F��V���mLZ1�[I��1$�(t%B�Nn��i���"��8tJʬV�Gc�Ƶf\%�X���׺x��i6a�8�r׮�@�TB�ZSb׺{Th�8+QN%���a�ǒ�&Q��#?��*�10�Fv(�d�1̄nB�yR3�|.t��w���JQ�R�-R�ȶ��"9e�I%U��+
�jǍ��WM�N���'�ӌB`��8�@z���yUW�)�f���"`>���r��?G��D����UKҫ��'�=�:�g�8Sz��~r42 !��RJ4ڊ	��3n5e���:�I�"��f�������!y�2�:,��8��*1c��h�9�daM@:��#r&	.�IS�r���ȟ,4��!�:y�h��&z�5�¾B��{��#�d]�3+��ƙ�kp�	d��d&��N�zD�ro�F[�҅���I�l�\�C#HNg@�����߭%��3��H�;M�4ߔ�[���'��#���RzksK��kS-|d�aa�kԁE�)o��3�ǟ}�+�F�A �i��Yoi�~��]�"���f�����E�l�M�,[�T�"��i���/���*
����?���?��������"�c�����V��hT��ޙ����Y�[}|?3r'�߭w����������A�6�A��o� /|��wbz����"bR:`��pd��#�bo����ZH	X�4�;2�h2��'�b���w߃��-�>�Ƀ������4�^���9<k�FEK٤�)������0�c���Ⓒ%9�t�VR5h��$�6Cv�!b#��a�.�P�5$������r/r���,�4�涗T=���cE��h6�_�ŏc﮽���0cK�M�g��/�V�im�A�я|Ǐ������+�j�j���?����ك"�T9!~�C�
�6:	m���P2�Ȅ޺�5���n���#����j��r�͋��w�O�đ&F/���,Yo?��NnTWY���\�T��r�i��6���O��&�@-3Yl������
\b�ٚ�����f%�����zrn��޾�I.��S�zϞ�>�`�'�������׎f�z��#�ʇ�E�B�"M�2]����Y/e��4�`���/��j>��(�!oQM����)D�ӈ4�D��"`oX��,�M�س��x0���-����G�`�dQn�����Ke�L����w����ܽ��j����fSqZ���q�[&��p��/�|t��QM�
�Y��)��m&�,�љ�>c�C�ڈDli,&@`��A��C�Hv#�<��}K"��J~!����	q�����#��/ѻ��**=�fsN~U;������Z�eWmD��(��ƞ�^�-�e�L\��*n�%�&w/�Z��ĀUeR`�K
մl���ϩ[�HD)��B�n+[;{94BPҥdW�wT���j�����a �U��_L�HK@@5��*��L�1Z��*���i0,1�V��	� B͎��G�cf�B4@��J�e�.H<,`�l������DY�.t`���#d�Vk�" �&7^��1X3�hʮ�fw"hȽҙ1���9���_c��k�����n���R/����E��h@Cg���o�5�(�*uD�%�	uv�gL�iy:P2z�Nt�qq�]����j�A��ҍ1@����+��(�&���\��VW�|E6I]��`R"�bQ@,��6ך�2���8ٌ8�
�T��u��eD��fr*n�s�΢r|��;���75l�]�����=Q�` �C�Z�N��[��j3��WaK�Gǰ'��Iy�eP;������x�?~����ȣ:M�}`��!y��˗q��)̮���/��$��3%�*�4�U۽%�����M�җ�k K}�>�#�t�R����l�i��K�f�	L	h���,�3�)�!w��clk?)�q��&�����#mNf�H/�V��ͣǱ��Sػ�N-���Q�7��Zh�긼<�s�N�|/�Hf��*�/�c��O�*�'���2��(6�B�X�L�-��OX�;�{-�nل������D��1TJ8w�^z�0��=�W�}M�2��u��h2���玜��K�pgnf��H�k�r�-��C��۾r	�$�w%������l͑��ٟ�8��_�9\�YBU��?�� i�^U�#��Lj�;����~���)&�ܐDY�����X��ϊ�_m�Q��H$%�iY���%��c_*�y��TQJ��!�6=k?ʏ��0|���k��3)�V�~*�g���u�Dm����SG'�CN���̊:��l�!(m`U�c���`�h������������3Ҩ*���m@�ǂ<U��	�n����m3��i;�;�]��{��R�-fC�����C��p��N�C��ft�u3�n�Da������fd�mE,9�̐8��<�~ˋs��W�V>L��sc[`�G%�5����[�d�\��{Q���ԅ���p���8�o�"�/e��k�h���'��#eG��2%Zߜ2^+7a�Rw�7R�J6��#{���%;:!�~�����j���-�C^��d���|}�l������%\��!�e#3:��b��;r�P�2�^6��ΉdVK�];��Ţ֦��4K+�/K�+@4��fy�af���������[�q��e-T7��R=T/.(�����m����AI�������Dڜ�e����*��i]�T�<K �^���}�َF�,���'�Հ5���IP��N�˦&���A`/jWKI��A#�rϗ�j���3�g�Q����7������`o�+`�%@��P#�iǔT����~Ӹ�o�f�H��UzG#/�ڜ�%�Oh��=�1��Y�&�39��5���p�J�1I��1ky`��u��a����	$�Y��lyv��<(��`ٝ��A(���4[�6� �#��/�$)s���̪ �ֹ�h��6�/2z��hld�8������,��.;�O�쩳8q�$��Y�H�T�Lm��ro��J�=�B�ͥ���hy�"���1;� CgY*A'Q��of|��h6���%���Z��3�=43��Q9s	o����Z*[�}���$iW,*�t 1
��%�ơ-��.�2 ����vZ,:i>�~IQ��C ו���i�x
���[~��79θǝ���?J��y}��N�(X��A��N������	}���2~x��m�ONi�M �l,Y�x�t�D^�r)�G�338��������9<�����~��F6���Ө�+����5�X�^>�*�x��)x��G2y��.�����！5�s���~��WT[�����m������� &K���|m���9AR}�Y(�uY�^٥�T[O�L�P����'����8w����>�lF�K�$r,��뵆�,>��S��
�k�B7+[&9q5��ۄ�\O��I��C:a���ZP`o�,5�v�+'կ���b�iV!W�|�u+���o7'�#)We/��,�R�m�'���DϽ�v�_?�5�`���(n��Z�5����%���j'(� ֡h��YP���;[>"��3T��� ֒�!A��ޓ�c2yzp�m�8H`~�Q|?���:QSz�!%�'V؃���sI�u�51�V�Jtkn���ӯ�Q@�t��V�xIP���=<��.�O<�~xV�D^7� 䟈n�S#�H�l2�g���FTwS�E<6���z���;Yו��D��F�P;��oa��;2M2G3�f�9��D\6#Y������ r�1j������a�ģ���q�DK#G��r�J���ʡ��|F,�40�NH�AN9��U������c"�a@�U��a�����2��nݕ9�˫�ɵ�&�PO�,� '��� 3#���?42�}nss�XYY��M-_8]'��\�<�X�g��� =JV%d$YVf鏀F�oo>��
'����k��ß�M#�G�Na���|�`X"�ɚk($#�/� ?&7��dsy�t�Ֆ��	��\kJ�Y�uv�^8mj�i� [B?���oZ�D�!�n'�Ig+�߱W�%Q�H	��Z@E����(P��E�}ÛX-�#�療�P`�}�)��%ׯ�2<��D�rJ�FW��?n����n-6T��JpjX�AJ�:�'�r1u�$��@���_�i�TE��@$���3����$���uvK��ڵ��)QyC'���L
	z�uW{���yom��r��j�=%(H�OKaS	Q�䗎!�ʓ �H�Z����4���?t���}�}�'�����ػ{�&&p��%�D��w�U�6Z��}��H�H�CEf[����~+��s�2Q]XÂ8�اb�����"���9�4=.+�Q�h[��R:i٣Udd��R1TiS<�{�YJt����H�T��Ⱥ�����X�g4�0M�Z�l�pT�=�m�1��?�u;(�oK��������ˡ�'�rYζ!l�bKf�	 ��,�|1䅀��;�Z��:�f�oR��������ɏN�[�jsÞ1-�� ����C}94� Y����/��������� V�VUj�ǟ�� ��}�X��E�=�N����"M"n�T6��3Z!�ʵE�o�,b�'oTS�O��(�U4�ho=�"��ņ%�*36s�:�8rQWJ�46��|��h�{��Q�9Y+�h���*�f�ɗ��D��������V`��$B�ە ��b�/�-��S�,*�+du��s�����/˵,���SR���R�+���[��/�ԛG4�J����!e��{V���u=�b���`�=Up)��*C� �0��t�ᙍD��<�>��m�P��A�=U0
]�{���i��)�0�ܶ�C0j��N����3�`�����Z�7�b�F|4�a�����so��-�}��&�!d�(!s�욥k��d\������/�闛�;�)�쵞���F۰��^��:x[�3z���p��O��G���T�"2������R���U>��>0t�C�Ռ�D�%!���e�z�Z:Z��2�XX��5��0��Y��ZD�
�^��<�@)*L^H5����o�}o����N���a���S\Վ�sپ�%��o�]�0:숑�2=V:w$~e
����8N+G���.�~�3�%!5A'���$%�c"򜦔���y��4~�Nc%��~O[�tG>xX���~1�5eqy���q��8�P\Z��!��j�{�UC!�6�䜊"��1zY�mR�̤:1�_�		(JE�)�ǖX��_�b���D>�|L�~��/jbpn4WМY$]\,W<$R�������$�m	(a����
E*,'�ބ��cW�J[S�u�$�C�SsӛӒC��C�#WAA�Z<I=ڶ�n#�e���Qgf&A"f[5cP ����='piȁȽ�v���i#�9n`��	Rx�h�<r�y!a�e����ak��rB�d��xv�ګ�=��W�u�)Ԋ�>����g!$o6@3'�%�I`n��f]I"��r	i���?x�*QT5�5��r�
��=2g�8|#O��1&������)5�:Iͨ�7L��s��d����\kG�AO"�'O��k��{���\^�L���\9��,.(�LT։E�G&�s�NtrIćF��s�O���nOo�};�`�+�qm���>i��n�-kO�g�����?f58�0-�`��A������$�V�9f�	�[���a��=8|�4^$#@>e�me?�%����T�?��^���rB���3ri��{�h�6/W*��V��@�d�	��0c���ܣ�����{�W�n�ب���ya�l=��녓��>���9P�`C{<זU�~`h����sΝ>��s��<��%8�!M�����(�H��J��'�R�n�k����i�<�
���It��A�M`efV�ˊq	�#�&'�s��������5*�$p~@��$���J����:hEr�R2�U0��+{��\ZO(H�! $�FR %�!�fA_�LZ�w� U�؇�
���*φ�����	����x曳��x����A���M��P�M�ק�Ѳ��=�\s���f0�]�G����n�DXR5Ƌ�՗����:w�������W������~��9�Y��,CS�uM�Q��<2Hko����g�)^���ʫ(BT��y���u2Z���qC�rzz�
a:nG� �q���۷H�����8���'�1�dʶFʇ�����Yڨ�D��s���4~~���#��C�:y�b�w��� �cD�iC^Kp�~%��Y��l�jE8Kn��	��ST�7%=�����)����h�+�6"�L�=�o7�K�̒�8Y��W3�o�RR�m��ɟ�f�-E D[�a�\ �]�x�����X���X�{�����فaS��8:���פ\щ%������Q�B7̬�:`²i�7 <$�:.#��t��	��r�	�Y���}�E"մ9'ɘ���VJU�T�I���P�Wc�h������<l�%�gyY��f�X�,.�Ј��)X�uۚ�"*`�*�hU>\��B"%�L��U�ht�1oM,z�f;�
X�������ɟu164ppxa�U�TX
dc��]�V�~��:f.[]/���ƀ���@.0dI?��v
f����g&��N�U��磩v�4��
g��F��G�����?�щYoG��)Zt��YL��@��ټ\�Yf9�:��9I��~������7n�b*�v���?������p����n�, ��Į���,e��RՓh���P;�����Y��k6Y'�\��;����Ff^L�7f&Q!s($�f�� ҋ�:Q��Ɛ����a7ڨ��Z��1;0(F��v%�u-<���Q4Sy��=���bU�>!�7y�22'�[��Ȉ�H�q�
�o"͡�� T-!�3 ]�i���!������[M$��3n��-��i!o�m򥖬�]��̕�͖q�����r���B�M�/��� ��W��=�����1��й!��BU���=�,�3��5�%�L`?k�n�F+8Ӕ@��)����#�z}�k>�~9��q���l{�NE��[R�l*�|:�v�Ћ���k��7�bm��ØJ��
���!%�%�B�A`�M	����_��Ȳ�:��}9wN�1�A&�H� ���2%-��J��u(S%Yv��T��u�z�uY���U��%�Z%�ZRK1�"�$��`�L�tN/�{��w�_�i ���ݯ���O�����[�0��SeW�H�6�}��|B�hp���t�2}��R��R����X�Y���gpU�������y��9\��BK�~��T��"a(��MIī�Se�`�/c��aOa�;��>��u	�
x����cS�pX0f٫nl���*�gp�]�tU�Ė��������1���`�jk�5W����^��V����
{����?V_��m	�s���ܑ����lk�Ə�%��%U+��
"�a��E����@0�3<_ʭ]=yN�ŷ���)kɰ\�O!wB��Ԕ+7���1<Nq��m�R$A�+�T�XM�����{��v��eҕN��ĭ��;�526��R�)'i��(J�w��(��E�P�6$`�Uem�ȃ곌+���0�g���s4�J�#qp'�W��ZHҗ`$'�S��נ1l�������B'3T:e<c˿��n���$��R�&&sHE�Jǰ���v�k$uB&'w'��Of<CYH�lX����e����mD\��l6��/VΈ�CffO�N�[t�;
���/��P�?�������b�� ��EJ��&,J^��j���RF%�B_�%������H�%�����F]��pؕL�ӵ�iב�3/ԍL|�T���JHh�#'�h[[fM����*i���f��� ���syԺ=�c�zo�A�:� w ǣ���f{��p*���g��.��ֵ�CLX�!�$���{G�&׀by����ս�P��jrFf@�t�=s�3�j!���+d&�'��o��M��m]��
�\�̢��u�y��z�)�00���	j��lV]$p�qM�4V�T��e��@笰J&��Yn�RXq��Iʩ%ĸ�	�'`o�΃ �[�O���Lkƶ,�3E͋�"�F"p�U���R~֚#=H�IW�U�}t�,�s��-�'�X������4Q+�3���!�C%����g�� ���CSh�=&�s��Q��)f�ٽu<�kbO�mA����N���X���p��ިa����R,�d
*���=bPk�}�(ʷ����$���]Y�(NO]��t7ʓ���7
�y�K�M�j �ɰ�Cn���ڡ�3�
t��dTf.&A��'+�q[�����r��5���h���ףmV��*�8:��U::�^��)N�Z�J�@L��p\1�)a� w�|��|�Χˡ.%QF��@3 ��ǀ4�o��h�O-6�=��4�=�O>���Ⱦy����ob��d�-)�q��$?	}~��Ί��n�(�rD�k���ܴ&�ͮ�^>pbZ�(qq�9b����ђ{U��+��Bu{�=��i�$P����'��0N��]�
J�2~���r�L�ͣ_�i���v�|n������$f ��1UG9�u�����u��h�v����/�����z���:��e��1J����{7W�+e	�������������"���H5R�6�ar*�i�2~S\�X%8��{Y�����9o�AS��g��[��ܲ�a�;_�$xo@Z%�"���ӏ�~C�s�=3o��`��69}[����~��Z�LU����}��m`?��4xP���f����-��kWC�׵�ؚ��q��Q'��v���8�#+�����J�1�Kz�Q�qj��9Y��8�c~�Β���RBǤ����ClH��y%�S�6q����-�|��y@�A�p���P=��k�s��or�es��*�)��f��1�}��\h��)Y����:|��Mym�=����h�(�����������rQ_\�E�lE'�44��*%ZQ����=�t�NT�J��Q)M�^kJL�Eqf��۪��,���d�a*�Š ��2�2����L+R�I���~�ZM���z40� ��=��dʨ�0�+�
����=���8�^�iR�8�0�7�����N�(�v���*���b�8�Vk��#+�^��d����#���lgoJ`ڿ��[���R.�'Ǭ��aG��'�P��`cy�V��DWy.���R��Jqd���N\ߜ-�c�ack�"p������^�絢��b�0���N�``�į1ညrxK"�cǏ�Vmik���0��#
��X%;�-k5�EhKW�%��$��襼�z��2��*���.I#��_�F^+�T�1R	���A$96:�:�� 8Qf{�,���i�� �I��<�O��/`��	\Y_A�ڐ ���Hd-���K��
~K�r9��j+�t�I5[!2��ʩ���{�j����/�tS���ȹ�
E�Է�ȧt��YI
z��J��"(����$%�Ęv(AV�*URlnz3�$
a�n(Ͽ�H�)ʈ��D���K�XC�⫴ �ah��}O'S∊�	�>6%��d�=����on9�75���y1ab��3I���$�f�!iF9�s��eOM��B�����>p�,�S�%�F!-��K
�}���%��Sb�X�����M��Tu�)S,���b9������}�0�����mRո �Z���@�ti�*����Z�4K�ѧv4(I'LM�~5�=�|2xb�F�t��0YH�9��^��S��!���X�#��fc}e~h�^cpE��j��ItU�{V��N����?��?�/������{�O}���ٗ���6N�����;��<��vU���WW%)ɉ��$��%9��劬ӌث�Y�Ks�������v�R�'	�K/�O��\�_�V��CK���O|��l�W��IףǏai�0�*n��>�uK	�f�rȧ���{rӊe�eZLRfQ�×W���r�b��ݯ� �?-I��կ<�?��?R���E�`� ���Lwd/NLQ*�O�*�� @��]�l�y�5*��� !(Ċ��P���mb�a�z�����sWQM�����ժD�ϝY���+S1�����Y�Q�j"��PC\�I��nB����y-q��&�#[�<���d.�:����b�Cvv@�(,�������)��b	�BnS~.�Ω��D�fĪ�@ۮC��g��/��T�D1hJL�5�r��d�K"Ʉ����S�ߢr��To�X	�2!�w���,c�����=+7���$Œ5k%s4�<��4|�Y���M뫄��}�C	�H�<I	��#Pa�;9��jʧ4�۟�Q�)���\�Uq��%9M��K��s4�&� �Q��֥�y�ѱ7=��Ŏ��pj�g�l^�'��r-��m���ZHd$��EX*N�4�J��8��'�u����y*�c	%]U�WmIrӥ�mc��H־�{��6[t�	���<���f5)q:�fC+���M�*�MTw�6�� ��ժ|ã�Z�h���N�d�z���u���Ve���+�rv%:��;��ӷ��Z���"���+��������M,7v�)���mq�)���	�����aӥc�&�@�.�όA�U�±�m�)4z�q]���9��m���p:�-..IГ� �I��g�dqN0=%���V#Z�
���1��v�^"��^�0F0~����M;uÓ�%e����(n-������*��Z��~eURO}�c��?�,��E��,ƨ�����]{8Tǯ�W�G��&fH��h�4�0Zݏ�$\�#xH��X��k}i��K��z]�p�X�	���M�J���/K"�h��!���=ޏ���w60%N�'����s*�d������1����<�],?�},0�&�����Aΐ��U���l�=���:^Ա'�f95oA<�23����ܚ�p�\+�C	���瀂؁!#���YA�5��_˷ q�G�}�f�g�>C]?����p�7��s�:����|�W�F�Ŭȓ-�M)k+�}��tK}7ܠtN���P��NT�X,S��Pu�^���k0��C�;��sSL��wx��M��9�X�X=+lA�hT�`��1��NU�2!Ϡ�����0QF�^ӠseeE�Pq���8V��]]FR��ݍ)9�%q��o��M�*�f(6)j'0�b����$E	I�=Y��r�H�3=��<�+[[�|��T��w�m����=+caz5�r�-U7�	*�����g$�M�d����/���|v{{�*g}J�=��ϋ�U���TG)�2�b�[/^����-��) ��B`:M
	�N�y'>����Dy��ɱ�����a���umZ�&ƙ� U��r����W��捠3��	�COĺ��&�1f�S�*S�R7x��[��܌:��T;&֫��8CU &��w��Y�vzdP �*�����N�|��K�w���+n���=�����8�"k�W���d(X�f<E\6�#)�|r,�IX�VL�7��
`c/�p~���Y�#aĳ�3�3�8��,�cŞM�$R�|sd���I��ڵ$Kd�FI@U�T��j��4����!�aB��w��6���H[c��͉��a��qK����Ϡ�z�I��L�|�V:��Ӣ�-����E�N�� ��U��g��t�n�_#�<�b)�RHJ,]�Z`�1�=�՜lJ6;����5سV]b�Sˁ2y��\�s�$W1r�٤j���B�~'�H�m�|Q�����F�:��y	1���R�I��YK���w���tr(T���;�ɄUC;ݾV��L��>����}$�%n$#�N�[ʎ�f{O�tY֍'��H7�2۪�uq{�� ��d�������+�X()���e��?;u:(1�F����G���O�C`�;��#J$M�D	I]�*��*4$26�	ɡo��Y��$�c"���,��2�����`��<��E�o�m0�ļyZ�!���hˉ�C�8��Mbbb/_XEi2��?������˘9~�#@xr�''��B����r�b�͔1KKB�ﹶ�MtX8a)�b�}>-�b����=�,1�"� ���|n�&�K��65S]Y��}��G��=M�J��w�/�wѭ��$rM��IIݣ-Y׳(�5aJνVŎ8�Y~�8��V��e�	}�\�*�|q�7!�����۵lQ�%��V��;J4��N=�J��郎��LQ�xߕ��l����&�Ɖty��{weU��(�<�_��ʭ]Zb�?�j�:��k����&Vt�7��e2��>l�S,(1c㓮�;{b�*�k68U�X�,�o�-{��˸�����9ɳ���ȃ�c�Kh�P�E��f�O�z/���rB_��k�_@噯cj����m���~���%���7�Ҿp�5�|�<���om�౅#��
�mo�'x��j�|s��V0#�I��˥Q�����x�U�'	h$�x�5I^�Ť��{�>6�o��an.�z����	"#��a�I����<I�!�$�Y���_H�61�c����#λ)������~�ڟ� qSbïaܗ���^��'�¡���-�R*�����a��u�����砕ؤy�䖼LxRұs:�A��������'�k�O��P�(ω	BY�����	28Z�9�5f�:=����H�?��Y[�ħ��^��A'�� ���8f剂��۩�5�}�=�M�O��K��g+7���3vY�kL�}�m(���y6��J�q����t������z�P��<-����"�I�9�2��;�J�o�1�8�M=E�RЛ^C�֐�W��o��4��n�f(9źh����J���A|IdS0a��Fڎ.�ޚ�:�>���N[iط�:r]��Ӓ�FC%���	y�Ҟ��N�3�kܢwb�6w�t2�03�d�$`̋��2l϶�oR��'a��O�L#��)[7�����
�E�['�x\p�Jv%\*�I9��*�0�C�``s~�����l[�L��Fd�I	H�U�T�J��M�6%E����ܐ,t	R.h!���uV�@"k�>�ña���/+�kK�'��\ۢ��(?�$�@����:0��ej1jO�rbd"�����2��4�Z��8��h���:�����|��Q��wL~.2��k׮!� E�����P�X�
�"3p_7;�MX�� �
!��t��}�9FB1�Cw�ӊ)d+"�a%n3	2�r��JE��ܛ¢ O| ��O��amW�q89����r=�f{�X��f�����
��J�E�b�`�]�x���
�Vyd��u(�\(k��
^��}�{�@���9�?��汽�����nm.]BI�#Q,�!������;ߔ���-��$,��=,�.�?�!��}�F2�G��-��̢R�B�<!���iBI	BU���"U,����*��>	��$t�{�]��lZ'��N
�v@b�ȡ�$�[S(�{���1�-}ޣ��F���=r�>��ɚ���Ob����x]��a��5�·�����En���[d�v���*G���B!NKB8)���[�, ܫ<�����9�N���l�������I��2NP�T�9<1�c�6$H���1���&p��E����A!�F9[���zN>�3;{hK@��K��j�µ�*�EY,+ok(>�I̹?3=-&8%6�.��P1�� ��9�ًģs��<)�SR�{�V�@r�	>q
�|A;),vpZ����s�X5ۑ�z<q"3�4U���e.�e�X�i؎C��{�r�2���G����k��@}�z�r����UbJJ02��+k���A���G�{.acP�`�-0H��Ά�Ѧ�N�P�h�*��X����hTw�*�^���W��!��|�ĺ�Ĺ��H�Xn��R(��pз�Vo��e	CrXk�"֓҄Ť�Zĩ�U�u���aM=U���˱�)E�v0�#����D*�JU�E>`Y���7x�N�$���M�1�����A^q2j��n�,3Ĥ�I|ه�����#m����/�./����P��r�=H�䦗�TI�IVє�%i�&�k�{k՟���ڬv������6E�`%ɼT�hW��8Ո�T<�E�?���̴R���w-�%�j�u*�����:�|�_y�0��P�]q�r����.� �$I���nKN��*#��Rc���ԓe������Z�Bn���Y#��<�>�Oʪ\i�����{J/��58��m5%��MHF)���{P�r�����Zb@Rb�đ>��7�3Jܚ)t$;4�I�Z3���ܑ�9~Zn&��I+N��5:tN�Qk��]W��?os�`�X��

�����>C�M�J�1)�@HZ���ņf����K:���S>_2c �Zf�e-�p���`(K?HϠ�ex���j9	xYi*�H���`�J�R��fm*����-t)����(�p�,W�@�O����W�@}Ga� k<Ћ�yL&T�l8]��ȓ������TyZ񀥤M��ˡ��~�=�A��pus�RQ�k���sP���
2�7)�	�֟{�
��{��X{ozZ���IΡɵ5���$:��Z�����ȴ�x�3�%ػ��Q�I���s��'�f�RP�Edi�[r�ZK�x�$1���JH"u�*��|��j�U�yR��#ӊ��˺=ƿ���%!1fN>K�m�dgᩓ�⼬ѯ?�,��ڜ�Ĥ,6�Ĵ\�]&nl�s�W�y��L���}еm/�J[���I���[�ۑ���kN12�I+��)?Ў�9�G�<oh��2p*3e���ZtI�⎘����0��sg����[򂩖��jv���pv�r�ugX-VJH�L�l�<������_JB���'
�
��G����v��n߸�BFn��g�G�k��$�"t�m�r�>(I͏䃘��Ӫ�199�/|�K8#�v[��ͽ����ryM��>j�啕Ch�b��+�S*K�Ҙ����S�{K������>x���;�����/�R>6���ؾ����]\[�.k�8��J��%{�����]����T��xT�7�����Ɂ�i���Ŭ~�!� E� �����/��/��,[TA������䝪���ZY��ŋ�Q�@�Cd�;LnS��ռ��Õ9�:H��4Rr��榶~YW�'<�~4t6����CL�WmS6�9����?�XY�"F֐S����gԳ�}z�E�'����!�ؗ斬�4��4p0&I��Ӣ�Q�p�V�I��th�yp��B�쫒�=�bQ���s�e�-��L�y%�&�,�� �����U(��'�)�l1L#t؈gn��{)TF��r�Me�B��l�������xq�w��T���U�\�D�'������4�?	f��&�o���0)�x�Z�Ow�sy>��%6�Oz
xN8m<��1��TV���0����V���,şw�u�U5�WܢeO�ph@����x�\�V-���,2f ���W&om����j����/��E�x��/�9�B����f&�BW�wW�+J�=1�YY����dw�!N.`��0��^K%��-�u����ܪm�h�����f%�΃Y�87���1Цj��i%2��%��"����U����ۧ�Y{�@>8y��19�m��3)2	Q�c���B	l�9[,XZ���]k�mrD`��$_�����쓫j��9 o��_6���j�jh��n��ͼ�-oj�k��[�~����Wxࢾ��wб�I�x���G����i��%�T��/Uc
y��=��n~��c�ߎ;z3ǎ��`��*zr}yR��3m�}��GX.O���Z]t�8j�}��)���y�g?�߳5�������d�K�H�d�B	���������j������ߨ�1W��`��̐;�O��_����T��T���ؑ�t᢬�$�wݦ��]qH��H����=ݟZ��.!�*�Ç��ȯ���?��V:���T����ߑ��0���r�<f�j�����"���+r^���0#��~E4Z<�����[+>W�@�U�a�cܒU��kP ��p
��#�g��a�of�vcx���h���aW��7p�ż�tr�ޔN:Ow��jk��#�=���ۻ�>ǁB��ʷ1bx:���dKlӆ��W7C\G�I(���װ4Y�������Ϫ
ʛ���g����kT"ID?��?���I����x��{1��ø��h�?�?����<6%YN���s�n\E�p�a}����������W.����2��|�����x��Áqv����V$!g2�)��֓����9|�ZG�����ɇJޝ,Ѯ6�ÑCPm	����_I+5��o��^}�Uؘ*�=�D��i�r�?9e(�L	JRro*%#�� ����a����^��~ۦ^٩���O��GoO���/��5	J;��g nh��+�ކ��"a2�^��r�<�(L0	 ���}�%#���>d���@�'{:b�(H���dAJ��OLg>���]d@$Xt���8�W�<��"6z=�5W����Do����������Mu�7q�&��"�>��N������{�l+J�妬H�o��W��/�g�	�d7pD�#��1Tf��t�ֆ$, �A��CO�<={b�%���R	�0F��Hì|��j9���J�;�%��C50ƽg5U{AO��Ո[L:��tI�VQ�pA][��	U�~h�`�k��#��;?x��tT�l4}΅��'��� O���a������+X<<��d���H��(N�b�R@��D�B���s�Z%5K�楾�#��&(s%���vX5�"�(�Ġ7wL���ml��4e���Zg�3@���Ĩ�4XbM~��6m6�΁b'}X��IԾXFI�Q[�H���R��N��d�pk�έ,w����ѵ�!�x)~iY='�VUf��x��G5������ݭ�㷵k4Z���W�I#����Y"9V��sq�Oq�p���3
Vǂ�x@�P�	�K �p�>�\�J�0��w�%���	��L�T�ͪ���L�B���'Oj��n�/׀NI���ib�D��#��@�OB�<�7��s!�v.��=�,�Y��@��%����!~p�*6�vp�m�UJN۸rN��ILLM������M�(��ĵe�,�o҉P��)�T�I	����Nz�[(!j�Z�@���m*6��RV��rv��$H��t
�KT�y������ַ�V촺��iĪ_���:.4v���4)k9�@�3�t��I�	=�řAd��:�`.�#�4{{�*~�����]D�� ����F�?J:(��
A�gV����0�X6�ѧ�F<�PŜ���GIH�b0�`P�;�~l��ۿ4�tk_i��L��H^�y��N~���&��	�Lϫ�[�����������v��1����̉�I�Vwe��e��r���U�|�_�E�}����;��Mbaz����ȱp�2�e�x���0������p���F)�ʱ%�'����.��u�wA�c(~���H'������א �Ei���Vd}59U#��!Y{"rX���@r��0��$E����'~�o����)er�vR��o=��?�=�J�
	��N�ĉc�NH�{�[��i[T���g�噯��:tQ��|�W�EwF��������Sݷ��)^,��Oڪˉ�R�;��]��X��*����{Yѕ�B��J?aG��.1AQsS��J�N���!23S�J�H�᧊b�X�t3.(����c#�tz�Fʔ>��[HRFs�/�1�V�qh��]a���f�C㯛ycaL:R#f��ș߷�����D�\�b��	c�)�����3I�`1�v){ݤW�qH-�s�&�W�紾��o�ѢprMŁ##�U��{���ڵC���V
�
K�Cu7�R�>K�-�J�?V�'����VGJ;����}�у8�n�`wU����l�l^��|�CˀH��Tqm�����3E�,52N%���M3E�0B�H�A7�X-����HR�r����c�^��p}��9�'p�����;$�;�8/�M��<z�ۘ\\�ji���nM�_O�d�r��x��rC:O[e� %�gf~{�d���ke{JyСq'��8�+�H��u1�18k򞜫L$�cezr"6$ �H���ϲy_�H�RF�0���R���O��G����M7Uh���TYc�ajr���>�R����kg�|e������䐬1��F�p��A�ڍ�[&�����NT��}G�m2{q:�TņC��?qj9�Lc�UP	�o��.����n:p�WG_����c��*n:����N������@�����]ďq@�5R�p�$�:>n�����di9����M��ԑY��}�9��I�ܭ-�hju[�b%�S��,KB�˺c����"I��9��C��k�ӏ���z��F��"9�NKƒ�%�ht��rA�C(���ַ�$1��-��{�����U{��(�#)jr8��ؐ_�����������v�:j5�W�Ӷ[J[�N֋�1cA���i�J�p����ü)�N+/�ؚ������zq��@�V�DR�N|��&s}��*doX}���Ƹ;v-����uw�d�}f�%L����3���ܟ7J�����ݔ�D.�TV�Ye�NHR��~2#6���B������n�,��$��f�b�x��X�v���ׯ����8vhI�n�z�U<$�½?���8���LWʘ(��o�5�\C�}���?X[�_��
�]��G8�o˾���ǉS'P>}T�]����Ĝ�k�5Y/5�{S�
6��Ď\���]��W����!�MJ��;ݞV�h7�-L�g���b���/ �j�V�k<�_�ԯ���NM��8=̉��|����O��Ә���=�K��5�k�9��o��|����M�Ӡ���#N{C��9	+�0j��e��E�A� K�Nz_����I��D�t��5R��"�Ĩs����A��%�I��I����CT��[[�`�l�UɾVd���>�I[V2՝��0s��)�� ���5���}5��&`�m{��v��'s���P��Z5��˘�/���ˀ�15&q\ya��y�cA�M�B����8�	쒾����ʊϛ�IԚ�6.7*��$E�H�It.�W�zr�b��t��a{S6a�V��8��a6A,W�x2C�'���(������$�M�!���9���R�iQI���<r�t�I,�\TCK��+@��1�t^6F��qwYd� j�K�k����mǠ�"ugdU�ص�>f�ı�#U� ��|Q��5�H5wv������(��D���5y����S�Q|��4�e�V ���8Mـ��R�3��m3�:�T��T#�)]*>2��@f�V��x.1ʃ���+�^am�*VrX���"�LQS�L���b񎇐�� �n��׉Е�ϔ�-���r)t����<�R�Pȳ�.KF,�8Ѽ8��^M�G�;!��Ҝ�R�΃�0bA���+��#r�����,�%���dm6�p�s�!`c�}1��┬��:&��c�B!z1����ޮV�X���L<�:�sAʨ:B�.� � M�TS�F�a���S|��η�ǝwݎ�$�L��▥ŕ:M�Q���������)(Jr�ڢ���\,�	�t'��LE�~�?*�hU֢���e�L��*��V4Z!-ʸ�;Q^����N��]a�<q�����f��|�,�J���L`�#k����V���p���y	*w�3J��{Bc�O�DR�-���zrϴ%���PM�(��蚗�%�Vk*!t����쁎��j��]Y����~j�Zj I��«�*/+�Ӑ�IC�HK�f�)l�U<
b�	'8t$�bJ�aK��7L�(���
���XT�'Ք��N��b"#kؗ}C�G-�������]��������j�*�{�jϞ��^�������El91�wT^ح���1}�}^�pԊf��h:pB`�3���ƴuS��Ja�SӠ��K��[Bkt�S��d��a9%Jh�c,�`�w�)��WP�`�U!Yq-�H����7��|0�6�I�[t���O����롪$��'R$&5�R�|AU���F6]����P�M�K���|!��>�(~���q��;�,��������y����O����8��~����?�s����)LIP�?zL=5�R9�ӥ[q�w��̕�Q[�Ą�5V�w���\�~�+>�?��2'<r��P�����+}�ŗ�y�:2�2�8w	IF�R�%��������� db;�=����~�8��6�����Ӳ?K��?�,��/>��N�UV���������W���+���_��/>�s�P{��>-I�TW^O���T]���~r�4ffQ��Tq]��~z{7tCk$���a���fb

[p�v��mb��R��WE��VY��C{ז}��i}���$���访����ֆ
4hd���iqȴ����$ ������3ǐ���#�Z��P��9!7]�ϲ�S���鉋o�؅�͖�'�+>f��������U�{�PI�X�U����KPj�8��v୯�W�W#ܛ
9��� C�s�(Z�^��[�3��y��hmcj�9���&��.�>�e��!�e�p|;�P)Q�K�Lc��{9�+A�����(ɍ�D1��T��N_�fҴ�	b�,-���}1�	�
ެ�W�h�v�W����fǲ���w�<�4�bd��I�ތ`)�I��î�'�{:����D�A��=ꂽ=5𪰡-��	X�FK�C��;�zQE���������T�qnY���ҕY1,	d��v�4i�3�{ɶgA��#�Q�����^�K����$��5n�m�3�ku��,�^X^Q����%GnZ�9�%؀i��x?�M�H�9�Hi.�0��h�����f�����-DG� � ꩩ	�vwwG��x2�?��-�c��#�&W����
�@���L�aN�����|�ylnnbWJ�*bUt�����cC�OiE��s��Ӫw:PN�z��Q"M����px��<y�����w��sT��*��yN~O�p��K�"���ԡ,9���y�l�+�0��������NԱE�
�>�D�b�ۗ.!��#	AǍY��G���h�����{�<�y47V�:ז���Tͦ���2�T)V�&�����r�I�\�KU��^9�yy��Vs�sZ�y��W�h4�O��x;��� ��PR�m���+�(��tqW.��l-�Kv�����9��|�րv����@u�8�|�� _������UtU�0�R��L.k�m�)M� Vd�=�
b�Q��F�*�8�)��=����i�H�g�Z��@�����Q3�t�7�n[7�SC�h"5n�{�����>1���7��6p��zP&-�䏿��ƿ���>!��qp6���؉���}*�ctD���Z�vB����������$��3I�*���2P֌�����$����ҫ�lJzo���$��p��e�\��D��U��n�3S��O��R�
E�Y�@�� �{G�G���U��7���FG��W���#KG% gO�Y�/ח��z����_��k8q�4���M|-��9��Ĕݲб8I� m�'���$Q�ӄ��*W�@7���}�|�6 �{(���'?��˗�;��;X[�V�%�Z;�	#�J����ѧ�A誸�}9VU��\�wW��\:�d������{�[C/U=S��M�bK�Ƀ�f7�<hh>)pe:���}Ǘ�I�L��:�%��>�{^"��r��J.j.e�jeJ�qX�;�"�E�L|*�������Aa��YUv��Q^�T�$o�<���G
:���UH&bUR�u�����Yca�u��#i�j;MٝC#'�,�a?�S�6k�9;YN���x�~�֋�׹�_��T^73?4J/�ak%�p)��'���-�:;ˈ�����Hf8���8� UA3=-�l�C��z&e�4�iu�Lo�-]/�W�ί�����*�S%�%)=-�~J2���a"�!N�Pҍ3M����!*L�<S�	N��s��,,��P�c��'�>'���ؙ��I�+�It�c��B�V�gPYX)9�,U*M�6���ƛ��Н)�>���\I������vW�Jd%�zn��,��]�L1��kETwwЬ���)��m��#.0lT%���yQ�-#�>p���N�j���ܟ��4̄xͽG�H-�_��I��{5�9�L�_ni�K��
���z��=/ϳ �����/�x6����K2��*����}�[��gT�`�I.�8�,�"�7h��J�P�c�����ϵ�bόy���L���h����n*%K�ٰ��gZ�
���s�3���1Y2qQ��۸"N%�c.�8��n)1��R�+�\�����0�����Hp�V�<���b�;���Þ�#'f1��U�ak~A���u��X+�B�K�5	}ֽ�~P��=�ElJ����6�To`�ݘ�m���[O�/?���Y��ح֕�X(�T� ��ѸQdf�BB����&��Fؓ�O�_��+jC�o�T�
ǡlN�Y�#��&	�@�vc�����}�9����!B�=[��6�=�cErO�s��%YY}�`�]���
�0�1h�+^�o�L|�+nW���ח��)Kn�[R2(�d�7N�±
����>��������~����`0�����w]� ���}ڼ7{ŕ��<���í>���/���N���,\;��7�uY��R�loJҳ�-�$f&gTiy �)���� �aU	��Ց@F�b776�j�qmuE��Bo��M��&��m���Wp��C	��}�<~}����Ĭn��(��Ŭ�$^�Z�N�v�b�hӓp@�@��v�C'1�ZH�q�U����X��>�a�Ŀ�F���L���6lm^��c��y��)9�#(��S�Ξy]��49#����+��ħl˱��[E�W��a�<���j1��Tl��f�ᴆ�����d�t�"y$-~�Ҿ)�,���J�/~i�ከ�v���g�����㘝�FFY$�t�¨vv��n�?�)�Q�.�H�޶�{r��rߺ(�݊FXD��y��|6���0�x=�,��mv�X��#��Bb�PX���K>Pe�x�������u�0�x4���#ylL@�ih�m��y�"7I���(&���݅$Hg�F��>�^[Vu�����r�rc���&�#�5��qi����o�"�Ԩ]?L�Db�nd��WL+�
qiI2�;��x��}���3��>S,\���1P�A?��M|�O�t0��C]�)$J⼩�9=)?��i�%���2�¡a{G�i�2���SM�:(QO]�i2��R{�=�{��%En���I$O��Z�������m6�L�19���7Ѥӽ�V-a-�'Mu�N�:�ݽ�VI���[j�r]	��&���im��=y
�҄y�N(��vm{[�)�m ��(O�KaG6 B�*:�K��0ȑr��9q��kI���d#������k]o4y�t�'���{�t�	őd, ��/�5�]��.�L��c����G"[�|�>S�l0������ˉ���8"�U�C����3���Z�F�u��IhUEm�k+J���~a5t{{{�����<�.!m#aX-��S�޲�����Ӓ����vlLOO#Y��S�)	>R<?�w�L�.^ŕ��*�3�P�Ϡ�aK����iM	d�<�_�G��VJb�8r���_����=�>�����@��'��W�������Ln6jHI ��O�}�q���/��%khsK�BG����*UR��jG���X���1�r�Vd��ZLa�����,gKd�ؠJ߰���J�3��a��̫���2�������l!�d��"I�y�ffU-A�q��Ejͦy�LZ�U]�ו+�P�VQ,O8��������bʆ����ˆ3�S����p���$���*<Gt�v�q�;��&�9�Sy�8�!oh"1�A�5pCWY�A�-U�0'�6�:��Ǎռ8�c>97���m�;�����)dI2ˤZ����tP�Uqx~Q�h�P?�����
�+>��T^1��G���������2�>P�\��"k�n��h���ᣨ�	��(4����n9�g��5�ju]/����S-)�� /�Z�	ŕ�I(@�&?)	M�xB=�L:��.����)I�TOYί!���J���?��b�s�/,��Z=�����_�.�vAaTP<�)��j��i�^O9�Z�ט��T��@(fڋ+�w�aG�1h�[\rx� �ׁ'b��*�7�g�)b�Ơq��$FlYy_$���λp��-8thQ�gޫ00n���U�$�d@{��7P��X���<����$�ۘ�'P��M�yBl�A&�����_�ݱZ�N���Mcx�0��VO[�G������� �cG�;��U��.��&Dn�*���"��I��l��q�y��tF)n�E�>+E�9]�a�
o�,���mI��e�x8*��4�8�l,�1���L��ו��}A������mȔ�NH�8>؈Yl`l��V��5x�x�"l����gN�؂=;F��A1��k*h:��ډ��d[ggK7�"�)/�����4d���4�̗�ז	��Z�fۮWƘIYeJ�4��Q2x3�AaV�M���"�>Uf� >:�d�ӑ�b��Gi��tg�,���"�͗0#����t����m0�,�tc�{��5��uYE<��Gq��Q�X���$ӌ|Ɣd���_���-LH�F=ǖqm��5�}W�ev�A��2�����#�_Z���R���L���#?_>a�8n�2�j6�b�Zr����� ���1E�d�M���z�q���8�.�H���6_ۮ1K./k�g�r
T���Os¿!�E	9�m�O�!k�\Zd��A���O'�e�����}��ؚb����m��&)Iy�}y5��K�S�xr�&�r�}Y���ؖ�֭cR��R��=���_:�;'f��$`!2h;��R��`��O~w݉~�+�����#O�;�/�+��臞�Z��W����C����ؾ����L�>���dY�!���gp��Y����Ĺő���%I�Jп&��Z����1�a0M�%�u�@�D�w/bR���cK��`����ӧ�P�Qq���q��?�����Hllb*WV�q
�s���aK��ć>�~�GM��tS�<�O�5�y�g�e<��#��=�����^|��` @�K~;�AA�)���e2�]�1�P�ӌF��D�&f#7���	��t}:�Z|�8�<X)�[��Q�-6���A�/���%_7������F-�;V����#q�8��i%g��r��L������j��$�$G��?�8�{���p{{{���Wu
B>}�V%�������?�kg/����іc�����g���#���EI�I�����iM�B����+*%X��Bu}u�K2ԭo�~ ?������&�6����x��n�_�By>���e<t�x�����g�ZY2)b�z����Y*�1?�{m���?����+���5����v���_��ȗ�P���ݕ��/�ww%��krrF�-��=WjI�֮m!'	}=1�=2m$ͯ�d�V���~���hH�-~qA"G7�W%�7ՊywM�.��H\�M��2�6� pH���`��E(���B�)�Sb&7���g^�W����"�{�{5�������<��>&KA*�C��e�ݢ��W���_�W��[8/Im��R��"��-��W�V=�Y�K������Sϖ��^,ՈQuҁ}4LȨ���P�d�&�����RW\)���#��c�x��1�#��Ļ�[G��������s87��/iR=n��&[9�H`�@@|�Vً�r3q�)?����R�h��u�7_C��o�5�к��P��p=v'%�X�4quղ���ֱ|���YɮDu������Q��u��1�P�I��w)>���\ܒ\/.o:���o��^���]	<���<Gp�8��,ŐW%�3$vZh���Z �6�<���l-tX	1v��б$_�I`�YF��"�.��#|k�p�����02C�����+��0P!��\O�+��ضMm�#K��q���e��Հ��DD!xy�,��$hۑ�~��U	�8�� @���w=�l��Ě`R�Y���k��R�[�'/�|n��Nf�Ή�ء�2'+�}J�Ʀ31at�ń�#��IS�?�jW��p��Q���t�-����R:8�c�Lr4i;΢W��j
��8��?�ڬ)�Y^�p�k�VSv����=�ߧ<a���=�kN�t���;1FI��U�X�-�&N��������nRe�3'�^���ް�T�W��J��ԬJ��n�S�$���3�|�\���}��Id�g�E�V����ٜ� z�i�q���������[L�y�y�����#O<�!��<��W�����OP"���Kf��B���S�6H`vj%���~������U�}uu����84�����{~*1�ap�)Ꮮ)#�qQ�ae��>���%��أx�C���CǑ�rZ�����ϣ�`>YP��6���^*W����:O��mnl�%�'�����a�?[�<�	q�5�K��Va���[�kb���cD����딴k���6G�Ջ���U��G��
@�7�����;���e�W���,�����<�@���v�xW�}��f0�����tz�*a�����M&���@����^�c�^���j�?��x���}�x�嗐�%�T����NU޿�[O�ĭ�N����4����Q~ryc?��+��w��꒠�mV�v}�jU|R]�ѼNꮮ�I@ה�k�\�x�JV[ml7��m7�Ӫ�̡GI��ϼ�3�ϓ��!'�%yJH�MO�"ASʨ��ۋ8�����ݞ��.s���L,6��G��C�k#�egL֩�/*A��o%/$c�^['T���$X$���^h
W�T���M�=�">l��ZLH$�
i�U�����j����g��܆���ъ��-)%T�����������Ƴ���uj}���+'Ij(���U�4��{�{.$���l�$�N����½�w<p?����^|�U����u M�Ii��W�'A�ܝe�L��ؑ��uB�6q �ł=�f7��x�+&1���;�n����1���(D�@�ˢ�6(a�/�!}ۀ㙛F��pA��E<kKZ��>|�ډ���5���}��Ű��n(����#x��w�D��~��XX���U&Z����s��������T��ܗ����Y����l ���8��
n��sOaԗ>�f�R������?~P���)]-�3;Jq��8tb�$X��Ȋ ��$��R�\AGt��t%p����#�c���CYq�l7s��@�t�a1Jeu2�?�AH��),�l����t"#?����"S�[T��wۖ�<����M�o9���"�";똞��@zN�����m1|�[[j(����Ȕ��ݑl��#S�(V�x�M���*
��r�'�Sb1t~�� ���6l&ڦVI�<�3u�plc̐�W�\YI��~�|�Y�~�J���ʋ\nʐ�*gF�r�R�LĭU� h�6j� 0��ֈ�C���T,F'a��j�h`%�I���G�-8A�?�
X�9��7#I2���T���8���1C��O���T>ۉex�:���b>3:���FX�)H`>UAC�������K�t^;��?�Y̊#�`�Q�|�3�dq3�)�v���Tđ;���k��?���ۂ\�э&z?<���X�\A��b�ob"����o���2���"/�Ϸ/��F	�N��(j?>�����q�٧�/|��H� �$�/L0��)�����-a��J�Ѭ� ���㏪��|Vr��{���C���_k�"����n�s_H3 �|z͆m�o���#ȋ����%�;z�^�q��� +�1W�V���$�>�2���7�ޗ�?�c�T*�b�|����[m����N9��_rL�2�>Ӧ0 �^��/�ni����a/����sUA#R7��p�vk�v��gD�ꇣ���N��0�bl��� U�[PW�빀��J���gq_�uX`��U�c�W,Y��>�)^���o=u^z�,�_�P��8{�ǽ���Y���!����������g.���S�9tH����������.����$zi�_9�W�ޮ�5���]��{vxv
'n�����-��=w���W�u���Y�������;qxzFV|�V��O�[�VSI�Y��[x쓟ă�}[��U�}�MN���)����M�"�v*Oa��� 1��� ��x��N�iE�#�RV��vT9'Hi,����
����i���*aV�9����$��?�c��G��~��BB�B9�V4���Q{�>�{����,.1: �t1Z5�U@~�/���fo�����Y��ӷ��?��} �Ҕ�S�	9?b���ң=eb`��-f�B�-)o��ajV��id��Е��ݐ�>`'I�a����U^@��#:\�a��#��qp�k3�˄
t�r@��U`�^+�nM� �6ܟ�M/��۵�U࿣	���i�yv �p�mw�~��8�
�P>%�B���m��W�P��cS�	
t�% {ݕ����H��|���3?�	<���b�؆l��� �2,]15T���l��	r�L����
_}�����>���%Ы^Q�Q��Ģ<� �E{�ʓ���H��u�"����gq�y2y���א�����aI��:
�&y�b�$S�ę�9��h3�ϖ�~<ٙ���v��.I&衵#ζ�S�!���]y��h�z}��3�n�c��&� N۠r<���`�U97F�5�|��Jr�Y�I�<lԱ�m������,rS��sY���)���,�S�s:�O���B�s��ֱ��y�.\@���$�)�)g=S_ 塄_JX��G�p��ؓ��C�C�䇪ª�'��g�J�1/�!t���D�B�����deE�P3#�d�J�:�R�%TS8�pV���ā���1�9�'�<x4:i*e�O�Fa�Ҳ����ˠc�#ߵ��p�R�v�<「���a@x�bv���^��T�i"[����ʿ��Z�ju��k�J�$Ԓa�s�N�<�t!g
�!�O��+ȍ&�/�ڋo x���똓L?��:K~=�jՠj�L��-���ɓ��W���*fic$��'8-�Ӗ��ڛ�]�o�~�n|�W��s�v\���đ$Q�ђ{���hU�-��Ӫ?�~������7����I�������!ݥ�g^�(M�a8
�x�l�n�q����������W����?��E_��+'%������Ul=R�w�`^���+�8}�{����o`�����<u�boS֘�{aKb'��$����7Ί��ر[p��^<����x�=���sn~Q'��5q��a��l #�
֐���~�{���d���`��Gb~QV,�#� ��r�Pm��ʑJ �a�����7���߯&�6��
%P�ġ1O)���I��	�cƂ��gUB�C8��Bbw��A3�nRNك�#�� C�:7�c�Y:�8�F�K���\��r�������㟿pG�Éc�tP���Hr���<�R}�7�}쉧U� ���~������b�~��m 0�e�D�D����H��1t&��؄��i�=��A�����S-=^�\Q������$�iI��r޻I	�-�Z��ΰ�I	�����}N�eӂk�R�0�v	�YҡNy�b(�ZhX0���Md߰	�j'N[�����3b�Yh5vŶeT��%v`z����L�ٟ��G�#fdٞ�K��&�$�����mo����ܧ����ȍ�����똹
��XL�(��?�B��A�h�����WQ���=��>�~�lmw�J�Nɿ��7ړ������3��v5�
ǔ���e|��_�+��W�,q��N>������bw��܏=�m쮜C4}RI��n,p�[�I�Bb�x ��.�u�i��$�}>\����o����[��f���	�`D:<a��zdI��IZ�NL%YD�ꇳ�;`9�3�*G��g�����'�Ow�xJ���N�� ��f�zg^@�̗ĺ,ۙ�1�x��������V1�;b@;8rℂŧ&&p��%1�M�z w�a���ƴ<�C��<��������Μӡ,?������'1��Sn�څ`G���NA�ս�Mw*}�rΑ<�#�q�� ��;�[�q!1��t�D�*a��,�l���N��r��N�q�ohōD�=JI%�g���
��U�hZ+��iG�[e$�h�����3�D%��[8��X~Oj�����C'
.�yI��� Z�{X�ZGP�Bbr�O�O���	���:) &й����U$V����&���V�����̧HM���"�C�(~F`��jMy���ʺ�C�2��G�l��E�Ua�u��J��
�}Z6�S�SA�s�62��:8Q��̌Y;
���^�Q�D#ba����˪���Z� �����N�K��kg��J&���������zK�1���ƈ�$6(/�a���	3�b��g$����"G�C�	��3��^�S�Ld0�{YI�JZ1H�$r�+M�#���^^[�p{U	��kb��9���(5�(��m5��S�S"�E/+SV���&s)U��޶a[��'&��p9��PZ���u|�3���ݏ�ᣧѼ��&1����VW���\cŉ9���Xc��gX�i:�UsaK�W�C��}m�}��������$��w�&k"�0��\�z��wQ�:���؀���9�B��~9�W����1��H/,���(UF(N=�眱�x`�<ǎ8r�d=���(��Y$���?�s���Cg}G+�$��ک��2� �χ4U�TN�腴���j
�"�7�5S�����9�������gڻ�������ľ����u��=9'`0 � A �&!�E�liUvɶ䕷d����벫ֵ%�j��Z��[�T
��JL  !��`09�L���rN��|�w_O��Y�itx���;�;�|�;����`"�R)���1՛]�S���d�A�)��:e�X��P���'�[��B��}��l�����p#m��#�#q�ݶ h�^N������S�����X�4��X,��%s�lM�brU\�n騡J�'����b)T�5�/,�Y�I2�CT�������o9Kż��f�׿3%�>�`����u�+�VI���y,�Ơ��u��M��L|@}[����1lEU3�^h`M��;�e�.�t�.їAx�_������}��(�:*�2 ��}sm	78�+IX[�~�������Y��o�|a$��|_�+ ��l쒕�eI���0��t���d�e��J�C���@��UG��SuLR��a��\��rS����4[���+ ����$ٖݐk<$v�����p��އ�uII|�j�1�����'�v���KΙ�55q���⻻-�P�I�GRY�]�}�DR^	��K��9��p��ro��L�!�ұ�A4�!�df@Θ���|/�ۇ��y���kXY_S����3�__y���~�*���ϱ%>�r�pז�=����(��䜀�Z��u�E��u��i"!�4L�b��V7�;��?Z�֔�jZْ�כ�L����XŐw㾟o��ք�uX�����h�]oĹ�M�J�Lͧ�XI�7���`���/�"�g8�T�d��Y��%���|_�8+�[y��Gp��aq�g^�`�JUF�c08�����l�i����1!�D|��iD#	���;,-. ���r����Ga��$$�Z��L�� �i;�
�d���zSK��lV�p��ݨ�։�fN��qڳ�X���ç$�}yU����5?fc3��
����-�ְ�g��ZvP��1��1� ���fA�b������X[2�2��p:S,�"�&Mn�!�v��'?kY����i�	�8��	C.�T��	EP��>����YD���8M�<����#��o���de����XyM�IL"f[F�*@��o�[�I��ന\����kikVm9ޤx�����Vf�\�N���E3Xr��P�Ħ��F�
�@�P���	�S)�M���w��Oq��]tͺ���޳���թ\���>�m���9V`��V��=�<Kںev�mؑ��Zt�Ha%������y�׬�P�ϴr�����*��6����~��Y=[hnM�Ʉsy�Je�$x��:�����G���տd��?9?X[�
�9���L�x�8>36�Ν����ѓG%њFW@֗����[?y	�Y�������Qx�5#�#A�LpD�����޺�F���۷P-;bǓ�<^��^��羅국Zb�.]��Z�䚊].m���=_��fŊ]I�$I��(rU_!�#��4��z-JM�y[�O@�7p4$�2i�������k!��o`99s�M8>�K��D�ܺ��l��I�OO����%,��i+P�sA�ɤ�.�2��_��N���-�/������@��c�p��r�gs�s�����C�������x��7$�qE���BE@#'�k�hoahx _��s��3���5���G��d���{r���J�Σ���oScн�9%�/�m)(lsky�^gdC��c����s�uR��K>���jK&8@E����*KP|��s�crzZ+�s��x�ͷ��o�0'Jy_]�Ѻ$�T �~�[�3Mp��?��������t�w?������\g���sV69�ŭ+�k����h���8��ȱSxb��j9�'$�X[����P�������8r�q:rN�w���(�.Ir���w���$�M�:$�G
�F&�[-����X�\��b��
�DB ��� �9xF�oC`{��*��j7M<y�Y\���Q)�1�V��s�������w]�_G�WKA�O��6�_]��5��3���f%_R!|B)K��`i��B�@�P�t��nʀ�}��u9�H%**�=�*�%@�'��DZaV/�S���͢���;8��~<|�����j��[�g��������l+k�X���ܪ`i��B��Z�\�>�`z�����}:\�7���I��\5��\������}č�r�g�v�kcL��
��Q�:-W�\XAg2��T?��ů����\_o�܃��w��� �{:���7odWo�Yi��[e���zA��9.����C�6mo��/i��S6��.Nk@�]L���"��o)��s�� eqZ��FӒe��(F�غzlck]����IƓ�c��`���x��cK����Na�qX���z?��6��٫9(n�GL@&+]mm:� �m�tC@�AgfC����-��Z��^��V�i�
;�չK�|7~t["��$"��yثU�tںg�:o-��p�2yruW��kw�SoL���"��:7&�6tB$+`dO��!hy�0cۺ�iPW]������6ztMk� �z`Pz�5Q���ʡ����`+�ľ��4�nu`�T���Y%���:аuW1��8���%!�Sta��˵�s��>j��%�d����/P�s/�Uu�N�����w�j���jkUԿ3����/� �(�5����~�Zm�jo�_�G`g�R���j_� �jQW��fW���n7��W���e˿g�-�N^\�������J[��-k�ěۦ���*6�1�|^�?�e�����_��tYM����o{�rV��B��h)=)	S�r�-F�4�]���?�q~�?x��5\}�]<���O���[3K�k�ڋ�$0��*/�eT�^��G���V��N�B�'���]V]�Q�X��s2��%,��ÊӀ��i���7���b��]:eˉܹ�������
����|�/�!�X�(��$����r�7P��[u�ȉ�$�ߕ�Q!�����=���	l�"=6���-�Q�fU�*ŭ �5��###z��c����������4�HI��%��� ��?��I'��wwi�k���وt�j�5:y��>y����%�G��;o�뷰�Ζ�7|;b7lv��W�����7�)������ߪ�GT~g��E܁*6r�\Č���X��O��G?���������%���Q�dm�ib�GƯ�گ!=�/&'����}l|�o�5Ŗ�
8Y��\0�s_�<~��~W��O������ӟ��|0JE�fg-�kbb������Q��+���[wn�u��ہ�(Gi59�����׿�]L8���Գ{��w䢵�ŏ���ⷂ��Y7ɖFN�5�����\ ��/֧n�jߞ�'����7տ6ėǊU�R��_��:�+?�	n
P�<z�y�K8�@����4*[ȿ�.~��?(���8�u��'"�HJR���>Tw�6B��n{��<7=�%v�Y��}���t7-�O�G��*TmS�;�qL)����~;͡]�٧ڤfͧ��!�;}�t�TkUc;�2@\�@[�H��FW��l��PbH�p����MW����iP�׮�ѣA�hĢ�������XlѰ#@��%~jߒK�O��I�c��= 5lC0֗�z߇f�(�$)�>�;����C*�/���0�۷�`cc[�1L�*�����?�(����D�o�8�8K�/��-�=�W.^F�HZ� �5IDK��i�.r���R\ڞe@�����u= ] �􆌜OI��r��OA���v{s�~W_�Jnȓ6�F�%�΄bb�y��$S�L?vwM����B\g��zCJ[�]׈y�����[/|U��]����GR��x&�X*.NS�Z�"�D"�����ࡃ�&����$���1mW����`|������'?��<o��[H�O#,X�ci9���u�^�ɧU:w�;@���f�z�_��}{�.����%�Y��w%҈�S��K���>��'"U��o2K��>����$tm��qh��j[1���Z� m���K�Tі���vuM�~��w�i�/�+�Ҽ��n\�6;Q��0&���aP����]��l��M$5���A�G���a{��7�r�ZUb����k
��]V�x���+��x�xT]?��S��U�D�� uH����py��������zP,�_�J�Ѹ6N�= +Q��n��ce��S+�ъ����c;���:�6/�Ə��܀��	H�UY�a��������{0�D�j-�!����Go�P�:��	H�jY�%l!���և<v)_ӊ"u�2���ȴ����K[����%��:��# ���g�RÕ�?��G��q���:����By}�޼���d�M�7܇PbH7�<t�8Rr337�DD[�-::4Q��W���{������6]�L|:Lah ����=�@�Z���}�IN:Ӈ��3x��w�?�LcR@Y�r�,�f]Q��>�ܼv��lЙ�EM�YD^{P ���"���a��r&�  �`r(=�o� ����1	b���@jh 	Ib��"�ſMN�ǖ��O^%+�`=���&+r���14:�G}�sh�+p�ը9� /��O�6� �ڒ�M�߇/�y��5��x��jrަ��%�Q%W���azr�o�Ӎ�1���M�6Ӊ��d"B���'O�՟��v��IrH5�� OI �'g6��9+���k���yi��f�l���pe���ј\_�[�YY���QI0+�Ù,/l��	(�������:����e$�(���sW/2�~D�F�+��:�F[�+�N���X��q}�����Do�ǽ�X_z���o�k}�?|_�w�?����OP���o|{�8������xT|a8F1[�����Q�����b�ŏ`
�X���6��M�ݤd�ĒX}{�䬐� �U4ל=nq,ߙ��)V8�'��-U���W��v�4�s����/�N�������5y��}ch�5*�cU�����{��*
ZH26�}�6����,3ND9�-���� WW5]}��2��uv]���Vakcc��1�2�^Ӄà;�������6��\�P?1:4���q�B{�$.��������p;]Z�L���䓟�ܝE���{����jȭJ���ħ9s^|��2�v`��i�6<3G�{�Z���Į�j��zq��?�?�Mw��IU��;������C8נ��4pbO���Fj���9z��bK�t�-�΄[�{˞x0K��
��� 8����)�;wV�ވ�*Ͻ�f��b�8�Ƅ��ņ8�J����
��2:����C����
�ZF"bL2�S'O���֦ ���h�#0�/� Uԃ�(t��U��Q5@՜;*YA0��V����o4�P����qq:�>�V�T��6�Zf5���;F��FG�H�*m+ٮ��+�h�b)����~�zv�ykhbɔ�i�����S
�MqB.}��џ��'����������>��ъ�k�����٦7p����1�wW]o�Qf3qq�T0^R~�~tj�2�!��,�ߖ��t��Hd�aJ�a3
�� ���>)2�밐�)�����k�6�E0�ă;mJ��>^{.�fp(K�ڢ�I����%�N�3o{|�݂�F�|�4�z-O����~�^ypc�^�Z��U�v�ܕ��:L���n(_�P�)`cB�$T�))�두9<��d��V{kym㶶Z�ؔ��׻��=��R�o�ʱ���9(�}���.��g���N���*3�0潗��uv֑{fy����>G����E��?�-9���!&�Y�������{���	P�����c��i�8�}���@|f'��
P�QT�g��q�6�5�M
պ��\I�@lR<y��P ����=��i�A-�ɤ�_i��� �������o�'�������G4>�9���j�%�>%C��Қ��3���f���Ψ���b�S�e
T{��1G��J�Z_C�3lWWr���[.mn6��?8�j��5|mVx�hm�v;�ww�7�A�zg�=�H�(@�!�.&ד���rK�".]���Ju����9�,�ǙP�47%	M���s��r��J��ǥ��������8<��؟��:Q�w�U(b[���3U��yvM��Č��)��%�{�MW�Q���k�����\�  Џ`a1�1�u
�G���V�%�_�wf�y�H�3�M*��P��T�i�/��{K}�J�
�D�ܱG�=������M���n������t$AٟV.F��tqsv[e�;_X}ͥ������|�W_ÙB��5��p��/~�5<����c�����Ud��_~UPV
��M�ծN�n�΋���uY���	+٭a�J�Q��N](�����mj���I#�O��`K������v��.�l�,�`]|H���H�o�P����̎a��>�l�=�����^��z�L�T���^���0kp���CU���A�O����r��F��J�(�V������VD��=����7gU�8l!�J��yP�w�T��J�R��Wr�^$�^ɫ/KBy����(���$���Op����T��&G��0&'}bKܼyQl5��ؚ��(���^lV�:S�%��;��fM�n��Q̴�� j�'(�r<I�RY��=㰐^,{�?�B���ȱD끟��>�v^�X��/HkPuM� ���2�J�$A2�n��ؾ���A���T�}^�w��yO�U��y�p�$ÒD���������}��3*���J��`
)����f���̭����0<�@W�ݮ�K�X\Y���rSV�W%��@�68tN�˫f}��l�} ���jn���������� ��߼��I�����R�����m�p�n�F��9z�U�<�=��� q
�ں�H���R�Li��+[w�ru��Rb��@L���!�;W��A_0.+@�t`�����%a3�v�#�3p�,R��[��޼�>�Tf89h��:^H�%�b��m�l��,!�>�rU.��&����@$_+	H紭m8���N/[�J&c�µ<����j�|CoB��D�X4������E���H%�w\��=�+`m�_�A�%p�Y�ڭ�V�u"2N��ן�M+s��N{��j�fz����	E/;f,gR����K�������-u�neՐ|�I	���Z��l��њ�6ɘn�Pet�L�RH�7-��î���jL0���I2��������:7s�˖�f���'9�SÆ��Xc�(�e	�������m6[�J���m&����Y���Op��'x��Ø������a�_������":����� �S^�����H5ĉV��Q�5�����?��uܼuUw��ayM���ZK4���8��Y�e$o��LOĕ ppd'2r}���*�f�P�;��/#{� ����	�����jB��h���D�`��J7`*������kx|�l�S̬hqP!��-�`�%�R�V���y�,�JR��՗^C\�$)#�������CW|^D�j6��<���
n$n�5*	к~�*
[��$⚼j��AZ��mIb>|�=�g�t0f^@��/����^|>���}Al�mc�<N*�O>��~���VWVW���� rzz���n<X`\�;+@���K�b)A���O�:O�3�Ƌ1!$����67��{�ܯ�j׹�6��א��G�/��bH$���%8�ܘ�=٬*�9�qɄ ���U�/&�^Z_�B|`��M� 6�0%g�G�c��$���9*�j��$��G:a,I���QV���>���7.}"�Il+�]��~�šx���~�%�]��+(�}�܇��wv��x�q:p��:���i�O*O��>���r��$��I�4�h�W%���_l�����5^�lP�ɭ5r�ʉ��`fy2HH�&�X�!iB�VM+�~������l:]��}�M�H=.:9yT��:^S�'>	 ۞?
%��s�
�$�LFyAz�+�\r5yV�T�� �2dk�����\�Ʀ��m�����!1&��J�$NR�Y�x%���ĩ��Ձ���Dt���Q����zCr��F��1���A웚�u��¶Ң�od��"V�R��{F'Ƶ\<�/
��Y͗qSpɝ{��^���t)A[M�6{x�}]�|a�7��cxw�A���?Ց����O�:x���^��]o[B���9��k��Iho0pʛ.�Q����LN�GM=
|�)@J���z��?���2h��[�S\�h/�����_y����Ba�7��#������{�����>����ۘ�?"��}QO�ߓ��6�*�Z����/է����)�4���1U�.�hWaw*p�^����q�t6a���M�'�����8�.�C�Qc�
��Z��撛ޱ��Xr��2�d+��̆h�b�V'�l�dR���8i�����<uD�zf��jr%�C4��VV�D���)l����#ؕ̊�5�F��B�����F����}��vIV[Ϧ]K(�C荠@����z[]T�5����A!�:!���&<����`K�S��ħO�`Oؕk�/	D��Q	,U����
'�S�������-��Ɩ�K�Ͱ���4��]]h�^��f���o%\��q"��\ͦ�<z"��IZH��Bz�^�>%)��T>[}<Y��~v��UW���<p�yk�9f�_� ��^pB6�|;0-����-�c���-������r0l��mZ5$���M3$D��O�C��-]�\����~Ult���$�~lx��Hp��8���$�a˷����ae�'��B|��>|�%|"�[/|{��6ދ��m�����^��7�2�ܧ/�	��ü��'�u9�Q�z�Zթ�U:[gMn�(�İ
^
i�b;F���<�hO�ݖk��;%���!d,�Ut�~� �����'X��J��= g���Ȋ�m�]o@�m����:��j�ϵ[t��i�����F۵5y]]t�q熩�$�(� ��(m��mb\|�A�^�Ҿ$��$H�ղ�@^m|ma�k��e��=�y��Τl���E;Q	Z�,F�w��D�����I���#)g�JQ�^�	GVQ�߹�Bn	��hH��-I���cX๶��[~ʹy�ݼ�h���yL�����լ�*��3[�V�2�"	O9?�+Ibn7��Qs�% $N���Jr.ɶR����=������9u4�nG'~}�\� P�INV7�U�w,,�b4�BUlg�T9'�o������9�Ğ|�e ]ċ�A�O�Ǐo�zu�P
�\3'N�!��Ru�������\�� �Gϟ��0�ƨ/dƐ��������mNy
�H�L�O�Ym6*]�����j	�FY��+���"��䶜M�]��ĘV�yTC�ı�8~�&�lu3��8M��!���`5�%����qr9��a-�I�StxX �U3E���,.�kL��0��=�[1��3#�F�:�5T���k��}����f(���׉l��݂|��ʞ��k���+�?�.
>��ɖv�H��w�������J�K05:���F�Q�?tG����a�L��t��Zm#@G�K�O���� B�n��a��=�nP����Q��v7�����9D�*�`�Ӊ]�yj,f�J8�T�\��,C)�Iޙ"K�t�:F�s�3K<`y�����)����6w���C�2$Un<�K�]�Pl.��"e	2$���iH�@�g[��i���ao?����U߫/%C���z�Y9\rQ��00�W�U�����CG`|����A>2��n\�@e���f��%�M��d���Iv�2?T$��ڪa�G������kpj9	�UXa�w��n�A_#Z�������MՕ̯#ADG��^5�Z��QO���d��[��"q��|^�k�Y�C��@�;	޼ms,ϫ� �r�%P�6�?�.[=V[�+r�3�Bqm-rD[9|��4��}HWӒ��Hf"Y�g���0w�u8��q��k�Ը\���
0�yz��/_Z��RN�����/�=�R��3����rm�G���������� ���&%h�d��c{�Ɇ�j+��uS��8ɠ��߸z���4~C~����3)�Xu�`�'�*A�Vki9*�4QڡW���K�F��z=�j����QoM�|܀�k׬�4�Q�clt'N��#�<�ܞ�͜:ұ�I&��d����\ ��(�n]��E>(�&PS���v&n�PЫh���*�b��O[�Vu�o�q]o�Ȁ Ny��pW�����f�0%b��4K�Vvy�[�ٵ�J�����J+RX�e
��MnU��K�p;�Aye59��䑌<W,)�����y_-yu-��9�X�fQ�|E5G��`i}���ʥy��'t���"���7Z�{GW��]�����n�39�a(���q97+@��5��r5T7�*ӓLuM��c�ھGתw85JL�	�:͞��1e����*@�9M�������_�IlvN�;Ҟ2}}DqL|�I9�}�Jr7�q���Ũ6�r�-���Ziz4>6q8���zL�_�$(�)�kg8���y�KEXl��J�7UL�cA�rM�,�^p b0.IQ��lC�gYߐ��(wj7k�1y���RX���1���8⋢"��N�����U=�od��^��4�m9�E$�m�?m�dP�P�a#_����
�]��CT�|�v̧���n�/���8�
�h
7�[j�9ό��fC�l�][�9n��L2� �`q1�7�A����B�xB�7��.�9џ���#��>\�y[����sg�����+�ra^���ʗ1���X���BX�����$�Dt� �u�`Xc��N.�|)��r]�%}�U,�0S�$���ZMd28���x��g��� �?�'﯆x"$ �*�S�a��
�;;+IC�d(����U�Œ�����j���
.�w	׮��	�x2���/2&���� ��$��RC^�a��[��C\GFM@;n"p��$�����"�v�FG�bׯ�p���Q֭��!�w9@'��ǡ{����=�!�C��XY��5�>�#c���C�P�^���V�e\�q_��&���">���$H\Q�F����ڦ�+��ն~jt��SJ%��O��ؤ��Mn��
*iBTSp�E7v��-V���R\�c앚�������c���@�<���ᶠ��?��;��ƈ�z������+6|<��˒5����U����P^l*�[x�I%��cڽ��\�!���S(̆�޼�7?��n���>U���t&B:.�C"�*�w�O��uFK�X�j��bI���i1�2
��d}%�;�
Ȋے6�? @�8��\�r0�ȩ�b�	�f�`\2IW^��ziA y񁔂�f����r�&$w��T%[NíY�]q�]���6-Ͷ#N01�U?jb>5\3Z	s�W��$m �m%���-��-��7���ڨ�#OqZ/����V8�B��ˆ�8:W��b�� �;���A����JV�����@"* �떨1���f��-��J������:��)lw��9���t����3����̹̓-:��Nt���N�����6&a�c��h/Uy�2��13�ݱr]8�z�f�;;f�wmĴ��VR;��P?33� ��2��#��6itl�:�3Ch����Tt
��g��I'3f@�{\R�`�I�{ڇB����_@���R��:�������w]��?����{X��+6���C"ݧҭ�%��O�눍5�8;`G�+mkE�k��%Ǭ[�.}~Ow���/W,�0)M@�I�k�Qx##<��o����_����j[hH�;�,>\u�+���-��]4��Rh���FT�hL2I��krl;�^�]���5q��ɽ���ãl�ԱJE@Ji�n�`��PնU�nj���a��_��W��>7\#!B	����E��.�r�����<��׾��襹%��6��U�u�.�J{�l�1��׈Ż:�ªρC�ȳ`9^m�A�0���ð\�T8_5�>Ӓ�_�ųZ*�$�=�驄 �2&��_v���y�-�������q��B�9}���,�m��rx��dM�\W��X_J�������Z�u���T�|�II~M�o}���QwQ|ƩG��n����By~���3$����Ma
���䳞8}�N�ć�
 �����q�����Dizˁ��ێ�9#8�p,��o�5c��*M F:�C��ơ�'u"��(b���(�A�	�9b�<� _�`@ rjl�@�6����$}y�:����P�h���B�oVu�k8`���VLb�=��_?0�	y��~v�b�������`����-�����[1(���h��,^��1�՚�q=S�o���a�/�*��Ƶu���	`���}a�}��f���8M�)�UFR\���XyjJ��Z6��?!��ؼ�G<�G�Q���fV	��_չ�����kN��C˂C�k���Cc�?90l���MU�U���_HP�v��0/-�O����Nm'#  />�"��2�P�Z�W�`�T���<&�"|�ȭ~,�����>]CF����B�G=8-q{/��4,���~Q&���ę�=q#�~����������P��$%������$�Q���<��[Z���?��1�\�c��]ۃ�qR�������.�	`���Rt�4��J�b�EզXH
���ت�<T�rƅ�\���
���!uTꌼ���@�8�.�b�
����7�������OUK�LI
��h�cƩ��$�s��m�T@��G����YE�~_��R��M��p�3��� 6 O�ώ7��#����7nc����i���@:���A<r�ġ13����^*�(��2<���TJ%�2�R}��t%{�3=�U	�7���'�o+�-�^U͓ey�a�a><A�*�]�j,��	�䘑��h��'��m*4PE�q��Ӆ鞀�DV�m_��ۅlq\��h��Kb�b�����]�~O��(8�k�f+?C����,[YR̺|ޚ� [�laʡH�UcP',�)���g>1�f	�ogT��2��P� �a/ �,������" 谓mS����f+V�L��&91���$謫��d@�f@3EXl��>�nmP��a�	KZ1veKC�T2��~3��m	V��� "΃-	#j�ѩ*�3k�u���6av=���U�|����>}�J���\綹��K�G�Ǵź�����!�
�H�q���M��V�͙�����`@&w��OU�0{������� �9#�NL8`@r��;2'9iJ�郫k�:��t���=
��6�y�ɠ	`(�9$���].���5&*�$���c.?�-�f��jHy��8�`*��T���� FjIE%Ɋ�ř5�Z���l���3�ul��e!I%���-T������q��OE$��")�G�aP������5�;ڗ���%qrM U8�BJ[7jaF��f&��� )Ыʭ1K��<�2tc�LR̐�s�ｅ��y�>�B0���+���ژ��<����ny�`����bh�_������/�&efmV�&g9�N}������8��sx�3O���⍟��Z.��Ѐ\Gs�T,Z��O���>�+x�'u��O�}yF5�(��@� t)-�Gx�$���o᳟�+����[-h���7S)q{g�9�0����Љ��:�-��/v���Z�F�K�{vT��W�7���QI,Cz�}�������f��"	4��ġ�x��/���O������� O}��LVC���������ŷ��=�:���%���u�\��$�]��N^�a���d������<Ixnv���(�;���`p��y �ؾ�HF��^_B�^��r�o���3�a��ظC�cI��&�ރ[�����>7ԏ��׏�)�=6Cpa��p$����
V�vf]��\3�y�:Y��\կŎė�E��)��q��YlI�ܔ��u�a�(I4����
%M����V.*�gY$bb@�b�Ƕ������$@unc���>�qk�s�:�$�6"�ܖ$)�5��:�s�����q�^B-S���KCj�����*ȿ��-�L�n
e�t[a}�<K��8�'�+�zߞ�Hd�ԧ��k�g��,�������zN+��n���_���C�<8$���OC<�}VeT8��İR`���X{hJB��XV�lF� ��@�aH�&2�/z�Y���J��9 c����U���Ju���jH\���������fd
8`����jV�vu�9��,o�c/x���9����v~�d�����9��S�����B��e�޸������0���v_^��7��Eч��C*U����J������ (ksmSPA+Sm9����rcStH�+W��y����A"LWU���w�5�� ��~��kM�op*���Ut��֭ܝK�U ��zK�}Z)e��-��>���v�)�
z�}�|�O[���ƧPK���G�Gc<�/[���Yy�t�bjc$<�U]UF|p�\����3�u�ڇu���Ig~�Ž��V��oHFZ��L;y7���4�y ���	\��]F��o�5��v'�u�*AC�ܴ,m���6�
"A��ʱe���j7�}�iHʁցo�������z��z�M��6u
���B�)?w���)2�	��z�̶��	�R
�I����\�t+���cK����ڷ/;���Q~�[�@ka��7�~?��+x�7�΅��jA+#k�5��0��?�s��P��%�~��;���rFmlme�):��s@�+��\E9}�Mo;T���u9���T��˳�d��gB�w?��b#_Y���u���$B��$F -֘V�gH�g�q5�m�5vԳ��E�f�0����^ba^݅��]W����c�ɩlV�$�q�A�^�|�
rIh�h= 0���u�&��C~݌���B+G��\;��Eٳ瞍�-;=��Ӑ�����l���d�m/PkE�`��X2��>)DL�<����Ç:�������@X����HӢSF��1��m����m��(����Ï��_��b�7>���}�f��}���#�/d�Σxꙧ����z������qu^B@@�C����#O�=�}�:��>�,�;��԰ �>�.�ј l��\QU*kX;q�a|�����QT*5���r(GS�~)c�mnn�/=�ӇtG��̂�,	t-G+?Mr-�0�5�&J��SEa�r��4)��@ ���䇇��w$�MO�\�Qy���\�0*̴�_���l��v��A/ۑL �e� ����V������F�q��%��g���S/ �=����{cFW�}�~3r]߾����Cx�[��� ����������ben]|Py1�-&��Ő����]����vv�z��QO0�p:9�5�7O!�ә�p\���r[%v�$�%��[���Ӡ���Ǭ��Ė,�8򸃩�>/`RZt;K"�S��r����HlL��ϜA��~������+
�$a�좮�k3�3��Ɵ�7�`���#��*]��r�{��^l�*�4Pٯ�<�,ק��$ѓ�6��H�r$Yo��49ޖ��!@߱gdC�}�o,ʽ���n����XZX���=M�cb#��Ĺ3'U �
��9��Ė�q��!�%���l�h4U$W?��2[�<!iQ:���h݋�2���4����kw��^8Z� ���R�·�9|`�?�ӔN��x� �,9�HF���ĉm���A��Oy���HX��,?=��^�����nZ��2��yQ;bL�?r
��=&���DrVC�WWT,snaA�����b0�f�ԙ��~��)��w��M<t��dM
e��T1�D���W/am�	,�Ȟ\
s�pr �j4��h�����	֐XY�#�*�� �e�Cp�π8������1�`-��8��F:�ᐃe��5_
r,%�sr�Rp6U���T�����?�m�����<��t�+�fd�N?��d�~����)%[d���>��#o��u_V�BF��Td���Y�_:Ž���=���#�[�*�-5���*���Rm��HӉ��s��4$��r��9z��t
�&�]����]���Db��ȤS8y�,Έ�Q�������_'<������,���6�W�������Vv[+o���sYow��3�=��=c��W�$喙
����<���~�/\��cShs���t!�?��|�I>zRe�����:fI��5�5�ƽ{�,C ��\ms#��AV��G�;��H�t�
4�]��L
8�U�ϐ��.�L��iwteq����Z~�Us���$=1�ۚK��MfK�����	K\��{I�b��bF6\�/x�������"P��
K��|0�`��D�\U��v9g�\-Çө=ϑ���X%gU�;8�Rj��j�'�RE���;�#�~��{NY��N�C����n�L�둸�ޔ\o@�g�;*4$`p`#��\�%g:��cumK�,c��� �D2�D������X�TF|��^qK�:޼zSA��/ ����/��ܙM��f5���k{���ͻ3�n�q4�F�C2r %h��9��/�������[w���øS��b���v�
�}�=��·���.`niS�$����J��� Y�ח�W�Q��Ng����t�ؓ�i�v���4����?���M�ɟ�9��Wt��[o���5�+��V�� ��2�����߅{�g�17?�:{l�v�v�y���dШ���}9���M�u$���zvU���}��l3#�"�U`���������-9�/���}���%���1*O=����W���4V������៙�D�a�K�7U�E��	d5�;��^��z�<cO��`;]�6/�K�,c�	�����������168�J��j��t2�l\��)O����\O��7ph'@�Z��+w�'�\���U�����1�d?��	n�VWz���ut�&{�����9�{<�]�}&u*�ҠPa�r_���Jg@2�4�b����LH��+d�	�Ŗ��onqUw�,�cyi7g��NM�c���8�wǏA:�D:��/�kmق��~�~Y�ws��,,.�~�������X�1{Rq;���'��gKy����D-@�[�LF���6*����|͢�O�:�k��>��m�&��}�� �Z�aFvG%�Z�k�:�%���ǖ��{励M�*���to���U�x5��A7�<�z�0�\�򈃒e���a���-zu4�%�6�0{���+�#����)A�SXcjʓE"6�9ˮJ��MOcrdQ���D
}�&�FU���<ۥ1ˡ�w��>pi�a�m���{����z�
�N��j�v$!����՜	U~38� %�/K�d��G�42�V�x����C�$h�V �A\q*߯�IR�j�ψ�R3�DnN��U�Z�:�!P����Ga�d���#�H�t�
Ҋr_�>dĸ�c�k���B' �����6�i�!��V-6���x�O�����f~�[ �j%փV����o�� a�����D�!+�&_s�I�M�����dJ)Vs�>����Җ����d�Y9��ɩ����ߌ ��Á����#G5�#O�_���+�$�.��M;��1k�X��i���ӭ�@l� I�ؒ�� 	��7���׶1��D._����J`��~����x��\B�ͰV=6�ۺFnH�s���SO=�?��˯auic��H%�8~�z�<,�}	��p��5����-�E.�uh�q��9��z���coAŢ�����&�۔0��r�+-3��o��s��(�}�zK��r���z)aA.h[��|f=��P��mf�T�yNK��M}''e����$*l�5 3�9v1qܟܸ�t:�a-CN�d}����P��@l=WM&\�>�Nb�w���46�y�G�/�2�P�ȯ�Ge{���2tO�����y%BADXQ �nJ�Z�wd�~>����T4ٞ�$�s�ܐ$�U���:V�r:�x��)XE�E���x��"2¥��oUJ���o𷯿��i�rb�(��d�Z�Z9cU�]'���g�w._�C��GI������d־=�>�-�|d�^���.������ܔ3��c�>
yըmn0&_O��#��af�>~�����6-D��$ sH�}�	���SXe�&�uI������^y����j��H�d���9��|P*+�Prw澀�9��1%�;*����Ӏ��'uR���ۏ��\��[7�������#�t����>�x�x�$�]�s��^�;9���Q�5)�'"�;_��Bu?X��g�D��}l�o����З�ىI,��߿��O~��CG�"�_G��I�1��*�s�  6p�B�q�GΑ�6#`ʪgQ�IE2�YL���qU��_vt���ӵ��5Ce���y�{���(�p��w��x��jN$P�5J��V�VЯk49�ɤ�@����u<����L�Q�U��*����%My.�I9a�ş%%�E�|P&&BB�[7�����L�^4ɳ����X��`ȸL�0<� EƉI�
n4������)6�0{���8;D~yw����;�!6�`�u�'�M�ȁ)�<uÃ��D�~��@�."��e�n�B���-T'�o�c^~~��
��6�� ���$�'�Q����ˤ��èF���i��-W���F1A�G/1Ń-�;w���W���C���W�I�>��50��[[K��MEab	ˀ7*�k��޺+�R�/���LO9&d�XZ��
p��6J��r=@��"P�l�l��SkͱQ�JVz������f~��65�Z
Zx u"�ri[�y�$ӬWZ�#��;')ZJ��j���zpP���Q�Vt�-�����+_���D$c�"��~�frF��^镊�eO�F)\w�:ʇ�]���ީ�p��=C'�TqL��-GџA���r�93�E���dy�6�PՒA[2� �N��&s�;���!�bN�,[����$�~��q�IZݘ�P�ny�%����G��� ���L��r{���vwy	�t|���=<������=��EENf��m��-T�
Vb5��xv��djp����i�����4�3�*}�A����@?0��S��./}|��뚥�����|#�ꤠ�J�趌�&���h�ޢ�ɖ��UK�6��Ɂ�'��.�h�p���r���с��ܫ��|���%c-n-�k;9	c]���o����enݸ�Vôۇ3�s�"�^;��WV�X�`���6m�@�T�2Z��hcsk]+|Zq���Jd��2q�tF�w<C�Z���ցf�mP����T\̰�m-�q�%zT�7���D�{��=@�v!�UHlCsb�l]	$�XC�$06����g��YZM�����H�oHh���VQQ<�����c��6z�TBI�� ��ll#.A��}���*�T O(\�a8�eI:l���1P��7I�e�{����
��6l���|�<�������+7pj� �%y=r�<>�����_���d!�FT^Y��ġ�-4����t��ڽ{�&�p!w��8��	t#Б�gqUl���?�(�=**���7�}�|p�a��<�0��P70����	�����x綾Q��I�k�<�߇/<�y�§OG���r�>m|�!�^�� ���q��S{�+_�&��� ���0&	V7�í�ނU� 	��G$��g�¡� 14"6�b�_��WQ����Қ&zL䊕*��ůU���]\@(��C��ۇ��y��E݅MN�c�,S����0�=�(N�Lj���x��bb�嚊;�[x�8���6~��g`K���I� �3#��`<���2�3w$iJ�D*% �������$kC��w��O��\�紹|R��@h��\�j%1�D(��]븞��X�n����߹w~��6JY��5�O�~�[���?^�D�V��\��S�]��S6-sn��Xb��m:^<0b�ݎ)B�������j���
�jr�8�H�>)��2T�؍09+�Mۯ��V�׿��o���ce̋!�T�,�*�/4�Or�U��d�-V:����sp��W0s���R�j�<������Ә͈�b~a[�+��D19��
ۿF�um;���6R��K�֖q��Jٲ<7Ux�|&'�
�Hș��/+��;��|A��e���1�~����z[F\Ox��;��,7(09���݊����ˢ�r]j��H�*�!�k�A=�r9E�J�V��U���$mok��[��S5lf�.I@���L �|x�̒m�ip1m0so_x�1�	�ci~���!�몪R�&#C��>��g
� ]Z����5�-]�ľ�{0�g��o5���-g%�.1��-V���-Xw\*��%wɖLfH��b�,/��<��`�k��R�i��O]�lS5�Z�a+�O�:$�x�X8��]QΧ�fϝ�kY+���?��;�zI��v:G�u
���m&;�
���$�c�?��8ʄ��r�%���I�%�77@M���1�i)�SP�#�vuʚ<0�g3��\�O����N��#��yI�ֹS�*��Y�.�B�\��f�Q,�kT��Z��(����ʴ<��1 R >����q厮
�l�(ΑU�J����^��eV�|]��F>ü�B���U��;-8q)�f}qF�n���ͨ�0��=bK�# li~E[��� ���+h[��ƊzL�r~��U�J�x��7U(�9e]bh�8r[������tG�B.���N[Z��	yܱTZ��nE���'H��MũTšFt�%@����6�r�q��c*l��y{�^e��u�.�)�����Ex�<���_���<��t�^{��Br_�^����
5��;!��̑�EV�I9b!Oc,1�֝E4�#(�`4�@ksŋ�s��^m<x����J\U�ȋ��l`K�ܳ�<�NL�9�-*�$����xf|�Y�ǊfC��&�q�����G�k��_��k�(Oh��>��3��e�������� �7�����/aC��}����ػw7��.�3(��.��#�zH�/�����]���br�4BɄJO�{�rj�	H ���}��ϢU-KrŉG�!-��/�Ϳ���<� *A���|�������#K��ĞI�y�#���'�4s]x��R�5>4�������l˵��W����1���?��/�H.�$"f��|�$���������wu헞}�b��_��Y[ �kS��F��gnU*H/����O`*3��/��������SV����"}b����G���V��y�L�E���x{y�+�|I�"C�X�k�e�g���i�@X2�V1��$��Q�Á8*u����*'��4�JI���z��R�k��܏6B��M쏚ě]�*�N��=�������q�z�ɨ^ ����i����a/�E���{������L-�l���su-\���VW܄�nN�R���VEใ��s���/���t:�9g'�����f_�$椊p
�t;�:X���Z5miڻ$׼���s�;��(9�k=-��B�g�����8D�b1���������ۈ���9�M|��c��_y����*T
U4r;-?�*�u�������O,�1�k�W��{qnYW��bM8^�}H�A(!Ʉ��=�+�����!@]�)��m��4b��1[�O>e�f���A�G�7������aB�%�����T�|濃�*t�n֐�[������;3������W�5\+C%y�AU�awnڧ��z�+.�of�HZvA����7���ã'`suC�����
����Z���v"8z�8�1�^�Hz��Z�@H���7o�3ƓO=.N~X�.����&7$��l#��=������J�>��}❋�^�*o�B��� @1�Q��VG���l�5o\B+�]-�9����l̰��`��;�i��
��dP��	��P�ω�.3���n�)v���v�������F���oo_Am=�����i����I/�q��iNgi��w׋wOF�������)sk�����v��GٽZ�g�$B�����#ɗ`\d�SC��	$� ��h":�W��m�i�Ĺz�zzZIa���]Z����8�ے�R���-�A,�T���PY��	2��+��{�at��n�9���-�+�L�G�ͬ�j��m	N��JE��l6Z���Du���)���nı�
u�sW)W@�s���Z:�Z�������کJ�����A�٤���xHl��y*�LM����1���Q&@�q`�%Cv	y/}�cod�y��}�޷��^���3 �o�MP�D�f�r$ER��Ql�\��T*�*W�\�rIN��*[VB-�(."E��ľ�f��ޗ����n�w��^�� �j`z{�����9�9�;�#3Kh��`X`���w#:���4,g����E��b���4m�@P�0��5G^,)�S�Mar�1	f����{.�6���o:}��0���n���+7qu�ЌJ=<1y�D�UY�Fi�n�|zՆ:�p@GѦ*�b�3��:��81�1%Պ�}���hD���ځ�6��8ؖ�l:)`�� @;��=�9~'��zE%b��
�X�J��y��#pK����o����U��v�(�����B��*�HQO^���<z�n�.K@��مy�4Y~c�M����y�㇎��2mL(�Ae<���
Y�5�r�)�O�bЪ���?�G�����E<�M쒧��S.=���K�� {�r+�+���&Ӹ��fy�Q�؅Woc6���yL�Ǳ�|C%�L	
�#��4Th8#���'������O���ɡU�iF��Y��3�q�����o���-�����O��c�ǚ؃f���&&���}�fR��&0)k�LF��'�'VNhO�[�T,�[��Q
O?8:B��W
��ؕs7.�,+7n��t6��$����uL��O[+h�RP����Z��-"wt����ĩ�s�0.��.H ���	*�L��d��MT]S���x2Ҙ��1<1�MK<c�p���?K�I,�/`��!���Y�.�W+�����Ǝo�e�l�G�//0�0~r`�~�0ƒhC�o>��)�ڗ@ �="�����f�?��_űC�_�!���Fq��!�!~��E����+	�cq����Di\]^��ϼ�g��D����8P�`��S'�9t�6�B�,�e�=Y��N���uŮ�d�P��"]J�f�y�dK�H��s�d�G9��7.6�Pҝ��M*�$�z�,J�Pds�$��8�0�KU�*�GuDM�st�".yNc����u;rqq�RyDct$}Sf�Xv��xB��#����Vt����i��.�^P}��~p�M,LOabn�rG������v�]9�I1D�+++(V�b�U����?sR����4^z�6w���)<,r��$������m�L��	t�7N��F�﵌ѳ��x���U�hӱSF�y�tI��l&��#�1���o��AX�I�*��1S~T�&���gB��nK�̮�N�zI��@0��4�������@޻�5d����y�nW�/���ƞ��lݍ�x�Y��:��/�K7�%��"q+��� �0L@����7ڨ�9�~�����kMɵo�Ӄ.b�rZf��ǚ�P|<]��D�7��EB2�6�{|���A�cѨ�'���DR��cT<�V��Ul�`U��^M���k�|�n� �r���J�`�p)4
]_J��8C@5TS_����([=���k�M+=�r���ӀGRL'�e��jl��Ϩ+`�M=}��G��&�0�����-�e�E,�B�3ݜ�1S�#��{:	aR��L*�h{�����S�=���u�5q; l��ߒ���NEl,����#*��9=ul��\��@m��C,k�\�@6�ܕ�ؗʁg�9�	9�@�G2��#_%�to�b!pn���a��~�@n(�FY����M��t:�KD�U9S�'�nY9c���̷�ou�dgv�k� jR�Lu�9;�3��!�%pJ�ubi�^۩`JV�4�0��
�����}a�>���F :2�".60d_j���M��Y������i�i6m�gq���C�Y�]��	�����#���%�-��&Ȏ�8Xz�-��U$|���9"+%דƟ���S����6J�Hl|�W>���2Y�ɛ�N���������|Fױ�i+���k7��0� �Q��f� b�tm�#B��:��s���֔���%K��k71x�2���j�@Փ��;�x�E��&Ⱥ%�.!뙲b��_}?�֏`��Ȫ+L�� ���,|F��Sp7w���թD�B#��/�!��cQ�N���N����n}D�iX��K�
@������3c8=3�e6�ZZ�f�&3nv(������(�G�c�
�_�2�^��j���̀���k�1ޕ��֫�a��ߚ;�l#	E�c6I�匵PW����h�<���9��#v�6�U�H"'�JP�UM��3�8�8�O��#*M�%�}��
�^~K7�T���<&
��+���*nksY�c�t����E��a ��l�4+�󘙝A�������.rԖ�����ܐ�86;)k���{Z	�t~�7��mL4P�(HXAc��m#A��P�NĈv�)��H=ⰺ��Z��y��o�q|^(#�F�����my:Ŋe�H(&�͗����s����s�9�T�����S��	��=PB��+~|X��'>�AzB�n�1�<3�3hG�����JJ���ކ�v����J�1G�2� 5	:��dq9�H5`��2s3-��0�LqA�6	��4 �׬��ߕ� AF�2���.aG���ѬV\Z��z$@�(q�D��:rK�F�p(;f]}@6��]*̟B����ۻxᅗp�֎bJ6�^q�7��_*�B6���gIL�5���	%zY�~C[�}�1�q�Ids��_�޺y�� ����ݛU���"�����@�U���\C��R�b�l�,���A��:�Yh�8`9�^? ����k6����;�u�.�8"�Nz:�?hj�eÊ��l,ɉ�=�+��]-�j�RD(��/���%\�A���v���N����zwM�&7Wn`�Pu���ee(�o�?|���Za�R4#��X�^����������������u���G�p�aW��ɜ �il����\'� $ƙc{��4*u�ϻ(�zr]�6td�jRj|?�Nh�OFg_���zڬW���A���`�����%���(�C��u"�����Ã?ę�Ѝ���W.�<�<�m	1�!K�6�����1�$�g\�g!�D&�d�⼖JGtd�:r��"�^���U�9h�={qy����ɛ�%v��d*� ;l��Ap�V ��Ɇ�r8l���+s?F#r���~qW�Y��PK-���j�.���`(X��+Й�;#�yK���,gN�N7.��C�?��� OBb���e4*�Q�q��4�̰�[:��t~'�\��Nif��ML����T
���mvH�W7�sB4�R��������"J�i=x�d�M�0��a�U����>��mU0+kE����i\Z]E��5�
���!'�7o��[�jAM T�#��QC�͛�e�q��!'6��`��u|k�Z��cf� ���܈M� ���cՓ�y�Ͽ����rU�|qZ��~]�c]7ef�Jl���:���O,��:��J�uW���0y�U	V�Z7�xCE�-��(g�E�Y J�p�����@�j�u��I�G�xT��vfR[S쬎=�T74Z��,fNy"������!TJ%��=���k-�''���&�F_�G-�k��F�g0���^ ���o�m�0���Ր�6�癕�Mv?nO�?��N'4t�!���@��f#MBHle4�@\�JD@AO�֓�Օ��DPPǤ�'q;�8�p��y�n�)�vj|��GM usyYy��Yo��lmok�-�tN��'�+ˏܳ�fI9?)�ǜV�HUau�ΰ�����3JGj򠧴$��������o}S���9�		\�'������͟�����<�|��BR��z�te��y1O�4�'�Ǆy��/]���,�y�lݸT��:bm�B��C�%8*u<�#a�c~���B*�Dٷd\�MlH�2��S�'�͊��8�+��k�*��?4z�Ъ�U禎g2+�ϸޟ���\ξ8��rL-�Ñct,z!J�������-�Y_�D[��dA"é�����/���}I��o��s�'gQ�T�-&�'(���[�!ۡx\���6�59���r������>��O�ĭ�\��91>	�I��ɻ��:��NRTU%P?(��X���`,Q��E�����qMw��m0/x L}35�t|�1]z�|*�r�᭱���k�Uk���rd��ь�@�K7�#���Dv��"���X:%W�N�!N�(sO1�a�w�O��l1Fr�&���mq b������ڹ��U������:F����xW��o�t�2cM�8�Жq�=�����<�0S�acS	==�\��ɬ\��l�b�	�:��%��QfM�M�9�QW���ٺ����+]OeG8��mM��iu^t�Ȼ
 m��-�S�|���{���s�|l��#g��o��_��q)z�Q�Y��Ѳv�61&q�O	�X������
�S8���M'���S���6JQC��Ձ�-Y�� ��Dx�ZE9g�F_3�0R�6��z��ȅf+W/ ,��j��YF�ByX@XX+!�����1-�щ��xu�R��ef�	hF���x�����_�����2)��(�#�)�*�!��a�-�ړ�5q�]�d�p=z:���n@v-��@�-�l���7&�:��f%H�o$k�(^�1��(K�?p��kU�M[qb���.��P�M٣�8�|��	Ce���)#�t�3������&�2�U�\�c�kF��6g�Q-bF�H� 5nt";�y�-�#&w�+ד���Zg?���'WRS�~��9�uN���!Ϻ'��;Ze��V��3��
�ژ�XC�!?�`#)j79��͆
>�� �0�ග冀���*��(�j��s`A%'�k/*{N ����77���2�����T��8�,��1Vb\���x����f"G���]��pB&��w��C����˵|j��!�R�Fw�p�òb�Y�ƎFr,��f�	R�>�t2lw߽j�>H�x���G��A�����c%�H��L�!���C�Ā�BK�~�  ��IDAT����gg<��H��d�ZlLK�^M�]kk᱇���:�}��Q�С<���5�:�^�V��̲W{�[����u�R*�'��]I_P�l��(9��DB�I��,�[TBGҔ=p��E�\îE�pO}?K��AC)GjSGc�çzz�I @��fx�#=a53��D�/��9��0HV.;��]��z��+��m	D�,N���4�c�8�����	��S5;��k���U<�9\�p�ʎ�]U�oO�9z/&�<;��ݦ��N�q�A	ZmzH����11a{�xC{JՆ�c��ag��fp�t��6wLo����#�'�mJ��a:�3�b�V���v4=����*B��L6���o/MѓzAw��L�#�F��)���{�q�j�L�낞��/���?� >p�)|�������]ړ�C�+���JnK��WA<�FR]*T���|��?�+��P3C$���]B�Ik
\S�,Mʆ'g��� ����?�Q�����U�sLד�1d���l��+|d��)[|5^�x�K{HL���GԹ������be}�nV�i��Q�1�kv8%8�/,^܌�?.Q�o�R������mnsܶ�{�&�~jzx�`o?p�қCu�ۓ&��3[#�g�~�`=������c:~���w� �=�(��3󔵃rp�B<)k7��C'�D�ҹ�Y�76C�9	cqnL�W"�ZW�tݎ��*r�XJ��8v�]���F�-��?�.]#�˃K.M�;�]��VϿMa@�+8C����k�ջ��0��������2r"�3�ћm�ѓ�:��ٹ>��c�)�����e�#+".�������1[ń��ǉaj�ɞ�&�;�U_�ɺ�өU;h��+fs�!V7��[����9���\��8Mf���E�C�q`���r��1��Ӭ��ɩ����{L�M9�����������f���1���^���1Kt��<�x�d�����0�.a��VC�@�b�	��W�:]q�R�4����t��m&��ܸv^�+�+G/�̳D���N ���s�O�%�Ї�]̊���IbK�N0���(�A^���t4��g慳�(Dާ��P�֮֜ �y�E1�ɚ�¬�NV֣>�È�	bqN�`Ɉ�L��a��y"��G�Q���@�0�KͲ��R[���y�lr��T�Ea��`E �Դ��)	X�b�^��r�����z-̏F$+U�+7������2�Up�Y*���#���#�z!m�!(��mxHt��)�7��</>�J���*x��*�������>93�'�����<�L�Sx[ �R��q{�+<P�?Py��o�	C�������E�w,fn��v��L�;�����������TU�N]�wWס��I=ؚ��*�J�K�����y�vk�����~R�����t���6rة�����`�RI\}Ӹ�U�������;귩�F��GՀM΁�H�)�H-S�1H�Ö�.��u+rfon�^��ue?m�!����9bw��O���7z����o*�2�3��вc�Z��)��(v,����Ǳ${������U�=�

�F��jh�,پ�ܫt��[��ʅ���T���VUyY�C`�Ώ >�����M�ҟ�(��2U�
�-���Q�(ʵʱsy��m����P����3yF��@���?�s���c��[���g��d�8���g�+
^�M��%��H�����/Nd`Z2<0c>��R.�yS�>�@Hs�%���
�-�C^Dw�Y�*�z��(�cs���{1~���z�:&
����Y��`a~r�\�Zd��ko�ܷ�*���S"@st�ў8�VS�D**"<4(Qǔ�l�Qt�,3�ȥX�œ�SJY�r�����@^$J?��@�{C;u��.���_y�n��_�{�ZrX�q�)%����5��~�K!s]^��ˎ��zc*]�X��!s�d�A�ߐh��Mi�R����H�.΅� J�@������,Z�_�{Y��G`@�*n;p�:I�[r/9���Y��wm3�:����\����P>)F�L��lU	b8��P�	�I�i�4�J(��<��)_���	#�>�b��I�Ӯfc9��֊*��ꛮ%J�0�ה�fv�q���6���0C>��6�*�����1}A	�Ҏ1k��+�8z�H�ܿv�jS���A�3�a�Y:��(b\RR7�&2	�w9v�t�<7�M�t���¶�Am�	�\����W����R>.tv#דb��'��1!�&AZ�%Π��h�HL�1�a9�K	�m�w���)���,��p|�P��NI��o(��Q��lX����9|
����(������[?ƥ�.d������˾����ɾ!�#��䞶 W QG�s��M-_u�],�a�a2�B^.�پ��=*0��b7����(-�e �~<3!iv!��q	T��ŚI���!�[V�1��wz��M��Z� �W��Jc�Ɵ���=��h�~hWwt-��E�붧061�p6�Cج���+o�vC��I�ݪ �J����@Kph�Iu��&��]�R�KM+��W6� {vK�bQD�	�Y�������� If�x������"uŻ0+:�Ϲ�%F)i���������/,���r��i˹)$��
Y:mk�'�b��PL�_��&�+��0U���5�mƴz2�ڜ��2��*z�YB7��&uٿ�Q�;9�u9t��	�b'�l��Rs��)ʍ�}����s��� �VJ�3J��ut��G.'�7t�a�w�o*ߓ�bҡZ���KI�5)W��lfa�א`K@|t_z�~eb,' Y C�O�5�ȩψ��9�}l��
r�	�)���&L
�:��y��J�EPc&29�^_��1G):�lX�������R��I�l�p��+�kJ�I"���d����!�\Xa��^0�i$�� �5�}7��"���nҷp_�x�o�e�'�|������e�����{>���q�\}+�W�ruo��@"n��}�gL�%6�عK	3*�D�,$�"<q���i%����������w�l�:f�e4:M�(#��D���b&�gU@6E��l��93c��4�a���s��7�g�P:�ҶqR0�7i��A�L�t˰N�$;S�}�ZUu���X�u��+10¥�m��Z^�E�T\qbyL{�d{K�«�r�67��ګo��G���N�8*��#M��2:+�S¥+��,tw{]B[�7x�4���8�c��dW^WQ�r�-;-��"z�A�~��7�5$yý�n�
<zqFOk`�|}3b��m��d]���QNr@
�(��1�G�?�NmO6�:��mL&řH����	���Dtj]���]�s�\��8��l��Y��JZ�:q�*��2���?�Ͳ���go��P�n���uM�4?�ڙ�����0ch��Qv��yF�}�w���겱jr8�jKGzM�]��vپ�%N�R��iw��٫P�kd��b�vdz�xMӄ$,����N@�,�]*��D�'���(�3y}S�փ�z�����z�-��ۖ�%{��h�4���)�<�V��p�����02X���.N�=�L>a�}X2���#J.0kE}#����#�L;���5�1_*� �_�gSB�ofC#mcܽ �3�&�7c�R�wi�L}`��f�M8Ƥ����:O��G�.30q9�a�,�Ӱ���ͪ��#v�~����_�;�*
�4��&p��(c8���A��L�}>$��h�m1�Wo�'�M� 9�ëWu�G:�C+����k�˙JjY���$�bC�N��"��nm��vq<3�ܬ��F�vW�^�O9����r9��⸩����\�.|f�(<G WJA]	�Cy�k+�Vo�1_�����	T�'P��-v.�I`��cU��
�^�2s��Qc��,QR���ö������t�x�t��
��*]É}��20�@�������.�g#��XlV�I�U.)6=�^5��=�uc����cy,%��iȤ�!ϧ���
�C�x�=d�}`��9\@K� a�Q�Y���KdԎ�@��0l�x��2������ܼ�z�G�T<����V�ޣ���T�����uh%"rݚΏ�f�*�Q}U�
MӺ�)J�S�vF�M���b�_�UC�]����lx��;r�6��o�[(�@x���73YI�uL����%9v�G�fT֦.��ɱ��Cz��劜Mym��e�Fi��~�L�<+r��<&#*��r�9ǚ��{S��2�D�DL��aV:�_Sg��f	�'��tt�/�*?m9~��]��/�`��r���i`��o�o�E:��yv��j��j�:7)�\�Tl���;�nq��[���ڦ���r�F�C��v���c��;����d��ݾ���"�Ջ�?t���N��>p�?�}A}�)G��L?x�{A���`� ��� �L|0j�ʌ6^��7��
��ծ%����#�C�}+�_s�P��8"��M��V��}��X.��������0�R��>4. ����%��E�\}�e\��&&��p�nL�����,nm�S��g[;�⬛9�8��8���Aw�܎m��G�k����&4�gH�&-jƄ�t���=�#��&��_A/�#	�,Q�B����]�Ĝ�0ϑ?�8����D�b�Lwk���Pp}�"�D4ZR�J߀*2�2�T;&#�̃����M�W�+����|�0����}��{q��=�{r��} ���c��p�T�����'fj�!6e}���ު�r�	G���l
�����]DA�u��颺��Ӭy$�\HF�*�-���b
(��Q�[T�����%Sy���gD�=�\�η
��������!��� ��g@��>u��}���}�8�b+!�c�WW�s�!ɿɊ��ɵrrI�-�|N���ی�ά��)��'4P�ߘ�[އ��h�ɒ3�`l�p]�h�b�bcm���lj
F=�H���vՠ�l��ڱ���f� ׃g�sK3�}u}5N�Fth{Y�<Z��Y�ǫ%,6�x�Σ�������. ӊ0��AkX��u��Z���{�gu,��J���_�~��ƗK7������Y)D:!4sy|is�'�G�����Q��d�#ɪ��Q�n�c�<��1ls���A���֍������b�X�Js*B"�YK��F�����HN� 	y��%'u��7"��;���I<	����8�=��BY6�^yщ���>s�I����Q5��(�Y�P2�NJ�2�i��2~*ؒ��l����a|T�W]u�&&&�Px����Ť��F�	/nk�%��D
=qz����+��4κM̲�ufQ�^�M	�u�c�JP����^w	���K�Pv(��|M:S�U �A�Q�aw]�q4�`8���µ�]7U��꿩DŶ)�"�۔5��8�
����Tg�D������)O�% (ו�- ��Q�TzL�oJ %�y�g*�*Ҧfl��	6L���� B�WeoW��JnY��RӨ	*r�dS�׎�Y��^L�<:aٻ���yظ�������n�/<�k#12VO+7%�,�;bT����u�I�W��[��*`DA�fŮʽ���UKeSAu�����9�=���@���(�l���_���K�qYC^�џ�a��÷>c�&���U��xf�� ��L��u�(��k]���J�#=��u\�?��%cF��08e�����HbL%�R�i��A�򭦙���`�b!x���~��VP~����r�-#AĠ>��^j��ΤJ(!3W�2iy��Q"Ǽ��{w5W	���L�g�V�T�6#��YQ:!��?J�8�,
����SJ��lȫ��L��Z�G'���g�F��dR�!@1����Ϊ�W����]�����\fZs������ p�)����]�):ӧ�Yx��}>���k(	]��g�?l���oR4
|����&g[8G&��)ـ`�.0�ҭ�.�p^�ej�t�l��1\]%�G�p�L��<�	(���d񆻝�Pv�����
�fɒ�1��ʽ�$MC��s�(�Wۚ����d�����r���MSv��<s��Q�e"-��P�q�������]�~�g)ל���c�͉���ͪ���vr����ue����i��e"$���>��,;8YV����Y��F'бU���uhr&�v�u��-*��A#����)f� �a��d����
D+0���!�e�h�K��mL�AD���(I��N�Sg!��K;j
��]`��a@fk��V�m�
y�!���7:�]NMy�VU�_q��r����N;kU9�z"ZF�e��P\��c2���$հ���D� +M���	�3K��Ŗ��c&��Z�^��5���P6��8���%<r�*�>�?~�h�J�c*/�I%�,Ϡ�C^�+N��+k6��V��:,��]����n�����N�����G�){a%��/|�Wq�3��F����rqS�a����q�2*W.�R�a��ݸ�G��8��4y���$�h2�|zr��r1���q�\O�r��,pmR��AwS@�ٻx���jjw�	ً��q����!�n��q�fc����Yv�L�pW�A-��N������	Td��H���[Du}�b�&Xn�GLl����o~��aܔ�a�gq�6��� i!+ !&�AHD J�Y��2�����6Jx`���ذmJ��- �/�T*j��QDX�v�	��8�C�v����}K;7�#�h���Ⲗ�f�V�z��y�8���d&,-;�T噑����t}׌�C�R(�����[��k�`��4��!�!�`V�2${!ᅵk8^H�Y���TN)����I�TF�{�USJ� �qm	�R�
��}�cgc�HH��8J�
ڷ�p���P��(�H�a̐�Ϡ*���n��
������׿��[Ľ���B�����U�ّ���W���f�	��Q��v����3���6S
d{�	���_']�'ϣ�uu뛐G�r�k��]�����ġaDm���j��q�{����}�n�Z�t�=��P�u��4�����!V 82�]Ҥ�8���{����O�}�>�z]�n�%"�f�ɞ��UZ-��j̶f�H�_L��[����g�k��z�`'���s��o�ƻy�涬!��2�{|�@��)߶��N�#r4A�_�W�O̖�������O����:����q`(����zCV��Y	3�N6/��ń̀��O`����}�����	؛<���
|�����;�J���Y@�Ny�Ȉ�q�æ�AV�tJ"�ԌD�(4s�� ;��<B=�ng��l�	�iD��� GN����N+���i1 �d���`F�	�H���RPi��4��&zm���|[lL�
(�3���t�-�*4��s�J%t>-�:(_��D(Gk�km`H)��|�c��"��X��FF���T��	)�9�&�X��3��!˺m���gxȌ�/x����>�1��1,X��4SF�"'(���<>S�b�u���D�ј'����*��+Y\��e��>XX�#��}J>_�o��H�n���h6��Y����Cm�o�0�!ߒ��3G�:KK��C*j�-��r=Ӧ��z��ې�5��o��<A�<��-�4�曡R����UFr/�"��tV�ra93���f���(��&U��jz��:υ2���U�^K��ֺf��`��6��,��pW�i�(���� [�Y�mªtp<�G[������\�^����&�R�"ru�L�r$bX��g,�(i���ݓF�,����N�
��/bxM6.����-㣅Y|82��2>}�0���������F�G^�n��ukb�.�����5|��I���xxb3����m�MG?=�����tu	����e�o1�>7���^|�9�����T��k��nPYӜ8ށ8�fqK����$����L��C�%�}�#�'>��x���p�~�2�=3��k1v͓�Ό��_�t̡'�t�|��ϣ���ؔ�y�#6�թ$	Y�� �Ӕ}���PBI��l�8=<�y[��9�����݇k����� �^V]��kɺ��h�0���T�:e��_�ϓ�ىYy�	�{p��NĨ�����9���4�m��{�Q��`-��M������㳿�_���O=��^��B|��@77) G�⋷��<g�f�
.��%ȋ@��������7��|������kH���T���l��.�k{�]9s|�$�)�F��3p3�GŃ����#+��ţ����6�M$�uvdW���ԛ�M�:`cla��{����
�}�k��>-���Y�a3HZ�I���t��*�����=�g{�CO�ɿ�9\�r�������셴�������q0�Ů���X?���cW�c.?�cG���t��n���W̊r���Q�Yzt�4��M`3�֩"��D�Ј?�(�V�+s����J���� ����BǞ�[W�g:�FK�"��ӡ�b��m��M����P͆���NU(�W`Zf�J�cP�'���{`�=��%W�snU&_��#�`sK����K�u�eiC+|�0%��h��#h�5�f]�� ��6�K@�CU::�ԡ�'n�J���`�(gwU`���Z��u�I���QݳF��שO!	�=�����̄�L��)X��<������Q��e�tH"[;W�Vr'��&^�d,=��_k�:ؖ�׃�Og��^�P҃�&/�nYh��w��%�1d'd�6�����$�.Ar����AH�5�Tz�P]��8Q�S�ˤ󴉮�hX���e���h�l#��|�`ŔT?H���u���pJ��}��.�h���d�	�I^=0����k��W��3��WB�� �ݛM�ن��ǫ�5$@�׌`�b�:h~�&:��O;�C�j�h`2;���Z����XM�%H��+t��mv�}A����9�&�6S��UXw��Q��ցɪ
���zV�������h�K5qt,�M	p�e�爑+p�;%Bi��R��b�,����3�ΰhD�����l��і�Y��nX�ՆS�e�<[�B�h*�CΏіet�jx�j�"�1Y�)�{,wX�Q���,A�X�����3	��-�GgUO��!�o�R��-�6GTp/#Х���R����ff�W�.2-!�	P���jrB��b��ݝ��=�{md�L�LE$��]�}��	deؐ�I[^�&��C�>�F�P� �SQZ�
r����A�1\W��@�$!��F��Kܛ�=���qL������'	��s��,ªE���0"g0r����r����*���a��v	�=�[p�\i�&&!79�����>i�&A��Լ ���;����զ�O�P_pb���p��1�0������Pj��s���s���1�5�|P�'�fW�1eJ���y�N����ؖ��7�����)|��ߐ�����t<�ϝ@z[�
j�&�Pp������
z��;��=� ~|�G��7��U�����K�0�x��Q*7�i������
����àM��Lv`��Y~M�&r�Ҝ�m(����g�06���
&�f16�����
�w�2:�2L�y���ڗ1����/���������*�_���?���*�Nu�iT��5P��|���q��X�p{r���q͉�N��XG.�F�#�.�ӎV����-��J��]@�ԑ�����x.'�Glw:�������t4�C�~����zu�rm�{[���Զ�n�a��%��g�ꑓ��������H�<6m@�Mc�J�6�._���o����z�	:p�o� ���G���3ȑ0��)��³�����u�	��#iŵ� !����)X�u����%�G9�0�+���F	�w%��U���f2�]��*���Jb#βy�!����|���XF$�	$�T�=��;�������

�A�J���4��	���@V�\�dÂ�� �7�L������o�Ѯ��Z���i�i���D�ҹޏ*C���D���I�����)�˟*�TBnR_�J	��NԀM��4����ők�:��s �O����`=G��U��2%�
� s]������:U��Udb�Y���P�5$1�Z��;�D��ñϫ�ǁ���5.�o.T˧}_��<�z�d� ��D*m���^a�
�����Q4�p�W_��e��-�' ��cq�)���C���C$r`%�6�x&<1���&ѿ�F�z:PI?���ҞH��υΝ�+ة����S������CK��U,W�j��3���Z���� ��'A��� ��M���D!��W�n����9�s�,�kX�Q�1��m����pr������޵Th-%��vO�X��1�;��	�^�U��qd�O��-AIZG�E�*"�I 5�TK�8�0�5'�S���!_HH$F�SP[�ׂ�g�r�Th��^TX[�_ݒr�������1�܈>G�)��"���~̳eY�}m}�����i���Ks����Rzu���{=-2�F��>Ѥ�ک������M�< �;�B<��-�0Bl�q@��k�N@-w5;�
x��Ł�\�w%j_o _q1��1e�t|�r5r���::6��8֥�l@B�۰��BF�l���r��Ű�=��4����fBzè
�$"�]\�n��~+)`+�)���������~�����G4�9��rN��;�J�6�+m똴OL�#ӇU��7�<���u|gk��4J@��^K�����2y�ԛX.���;����ip���״�!�SF�uF����4��)��ٮ�o��Wᮗ`��;��<���El,��|o��M4���:$�iL�����#'мp������2�feJ8v�8>�+�Sc�ݧ��ݹ޸C� /�J���N#����w����{�5���w%�j��{��'>�1X�.�}	V�(dq��r�1����V�'�~A���̏q������L��y��g��k�v�-�ܸ����a��^�N���$�������?×���
SY�RL�w7�~O���ڲ6�\���~�z�1]�B.�ѹ9P8���\�*���&�FZx�S��'?����E�Z[Ö �z����<f3Y������B������K�����Q��CY|��~��<�=�
.�]���L����&��&�?�1|���x����������X<���/��^�j��-���=����PDY ��C�������Ϳ�v���8�ɘ�<1N���Gq��;��U��܋�#gQ��ko��Mr�tKl�8Nɾ[���X���.�z�ѳ�Q��O���(�����*i��j��-�8�����L3��ȡ�?��M�����:�V�FbS{~m��'�K���2Q�a�蔳����z��I"j��X°v���r_+ ��*`G���$B0��,d*u�[�F��ay��k�$�JK���+�Fg����z̺+g�3f��_���40%y�!����4���~(��?��,3�\�~݈v�TmO�Z�",@��:euv|(��5�3y�dף;���Z" ��WL+4����t1UR��k��^y�#A�k0���el���T�+dZ�=m�p�i*�Q�t�(�`-�!�u���Ηf� �������یb���o�s�����F���ݽ��e�Idy��-��]�	�[Z���G$niy+*���o�p���|�A;���$�0�$�oHK��'����<�.�Pn
�"9< �;���3���}�w��F8}��[f��b�8ᑫA-�Z����AR�c6�J���eʝr�8�!!��-���æ
��>�Ďn�������4
�q��ٳ+����8Z6���H9��
<������$h����ލ*?��I�LG�Q��
ሖR{����g�I�M��);���!W,����/yV߀�5�$8q-M��v�L��4�Z.df�1�cD���'��0��sMIގ�6���Z]� ��T�uѕ�i�{r�m�J^K@A����4f�Q9��w8���Z!=�C���L�����췋�v@��t)I#g���l>��*1�Q0?��c6YK(�Ja�8w�c�(Ӑ ����vMn��\"���D�͋8s�0~�c�?�KkW��'��TfU�ݒ��������f`���y9,�J	�O�&�w��P��l����-I�X��N��S�bJ�����;okP�L�01�f?� 4��3v�<�������_~]�� TY�=���)tS��s��U�v��������;p8) :�}V3ޅ�c���BGe�����3��<V76�����MXKq���������^���8��?��I��칗Щ��Y""���w�����O^{K��*ZV�>�$8�Nde+u�v��=�8~�i	~���:2����$��_�'O?�c$62��֜����_�����U����'>��{�9y#7]�D�#�ݏ>��o���{�%l���U\�ka3Iʎ��bq�(Ξ������/�Y7<Ӕ�i	�>y�p��͕�p��r)��/R�_�..��@Q��O�w��?Ƶ�c�T�m�>��{_�U��|{7���d������+�ߒ ��{Ξƽ<��'��������q�W*7�����T���o����Г�zH�*�7�1yw�s�Ç�u���\3�$�����e<������+x����rI��j��^EQ�����������������
Z'�M��8����3sFMOF��蝪�"Uf�݅-F���-�ΚN���G��Z���
�F`l�J��fʐ+��N�eO�Fi�F�m[3yAC�H�� ��A�GX�E1.��D�ث��]��.ǎK��Gê��*���Qn�o�b�&lj�F�;�Y� }�$Ep�'jj��Ć��=�f�6�\(#��Lq�S��?E�N�y%��:&�_�t�ket���l���Q�����?ㄔ�f�M`>up�i��Υte�%D6W�x�8�O`G�r��@V~\"⬀?��A[�h#����]�R�b�F���=�37��K�j2�M�ֺw�#��Ղ}W�ESCY�Of�.UĔ�Wҗf�T��#@���:?Г�Ԥ��-1
�^����{���'�\�d�zY�4P���7�Y	��v�އ��kז����cXo��#���.B��{N�ƥC�6�##0�CK�PJ"Or�t����R��㋓r�<\>���4��1$�yT*M�x�;�3��)v=��D�6ػ	 �qn֐�q����!����7�P��7�I�OQ�%Ps��F�ɍ#r�N̟�7�~�ֲ��<oNV�<����`��5��ֱSl"�Lf���Rq�CW�����w�F}�a\�T���}s��J6g���O�Ҧ�(݁E>yy:J΀<���m�N�9ЙMZ�uMnd ,�Q2ZBSjJi@g�J��q���� O�Lǫ���>��nW�l;�#(��\R��.�%�F�\���S�J�R�-[�����F��R��Z�E��!+ߟ�J#%�nC���;Q�G�Ҙx�4r��xM��K��{�cb/8���YY;fK�l]�t��u�\����-=?J���p.�o���_�����[��woY���ǒ����&�~�!|��i\���ڕg�U�CF�7ONf߬1���޽�U��?�;L$���38S��E�i����D^^G��|��~aa��E\,o�����uy�zSrސ����P��&�r/�x+�w��m"<=�d.�{e����Ьy��7���Z��K*$�%@������	^\\�?�1���Im�4�bi��=~���*a	ly֛*��W�`s��ɹYy�bg��#s�e	�Kl�F���������Q.Ց�@i�C�y��I47�~�)����13ΑWl,��Q''�5�k+����_�<<4vUNoC���ud�\�x	k��ŗ����?�/�q7
�o�X����N�?~��/b,,����N]��n�n��+/^�z����ث#������ړs���;��o/�>��,aZ�W�.�M4)q�������2֟>��Ǐ�7�އ�j1�SD9��V_����?��v��{)�NeS��k#�,�E�j	O��70�����b�R�zQ�9��f�կ}��/mmcyy	!9���޹���K�M����8�p�%���㙑=6І��jO���_\��[r/fsS���[��V���K�W���Ꮝ�����@�n�y�K�%��7�t,��=���=G�DF*̈���Q�o������Zn�g*EZT��B���C��`������Ԑ �$��ꠖ���@:ܮ�L#vT���#��2��(��=B9Q�MuT��C���) )zܑ�4l�
�c)[�|H��U	lЦ�U�Ȟ��h�0�3A�� �$<uɈ���[g=Ԑ���H�5��y�}���f=�Y&����v���"�bw�)؉c<�(�%�xF�{*�Aׯ�}���T,�/8��N����o�0�R�3q��섊Q-A@���.#Ҩc�����h���F�l����ɦ��tg�L���z�p��D��`��<�2� ��  )x��LY�%?>D6u�ZM���V71�$���>L�Z��0Ȟ�[�ܦ`���3��p[��=J��5�e���;0s���ۡ4�!�G�2��N����yUk��dA�Zg.(_X�t`����s)�)4\7��=7л��x��3���]��2'�K	���%�|$�9��P�Ĩ���r�0�y���l�n_>���<-D$�\��,�v�ʡ�Mb��	��b��:��r۰����uNr8Xw&_&�9pk���[Zi�;���%ld�a$S!�S��~d6&E�'חO��G��)̓�aDj�13R��������UNj,�uVf�
5,ɒ��g?���D��� �l���DȌ; )5�V�eO�r_�q�3�����Ϛl�Z�����1*՘���%Ƴ���f�[�<'YTZ}=�l���R0���!�i	��o���M��Q��Z�^��y�5bӉ6�;b��tk���5y�9{Y��gi<|��_���ju혥���A�8B\�K<+:Z��--�W�����7�-��XB����[�T$��컭��#���s�'�%�Ӯ"f�4x��j�z%�(�xnwM@e�����9y�禦�])������f0ّ���b��X}c�ԷU[la|\u'[�=u@�B��6v�.^������''Ԧ��J��?���X�Í�%L����S�"K�k����تJ �NcK�{c>tJ��З�*��SO	0��
� }�p4w��#]�Y3������T;r�x�c���cg|��M�X�TdM���E�(�� ){�e8j2���\~�L�S������an^6�?��?�F��/-�") 6/�������c���|�����x8�;�~ ��*�Wo�&��3?}������)4��%Ҷ4`a�z��%T��(
��`���'Uv��gΡ"��{Y*n*w9�cg��JQ8!��`]�^����W�<NT���{�e�)A���+��c�4�vʈ	������bI�\�37��j�8z�.]gJ�����e�������r�j�Fa�ŎQ��*c�����-,�}Q���#A���$}���E�k_C�t9�	9����f���x��~��_�>{
Q�ݪ!��Nv�x�:�,t�=GU⬥��p����bpƇ���F~*{u�o��!�m����L���&�j͢<ˆ\���Q�QJ9e�b�Mʒ��(5f`d�(��ˁ�w�_�$6g���	JM�(ܖ�=i9�}�*w%(�j���7�7����H�<�i��o8�[��������mWU,�@�*N~'����Ke�y���N)�1S�ȣ׿�jo���T��q���vC(�B�`�^�y�n�Q��2�=�ksb�)|�����X)����t��*F]ޜ*�qZJ�(@��Hy���}D~�1��<��Pk�2�����c@���C�Vh�k��<ߤM� g�Dk6~�=��� �c{�'P���F$䑈��Y������lT��ށ^���{Kӕ&�>�|�]�]��<h�O�L[��!�йA�x<�V'�#�cq�kuX���5�����D d;�T� @���j�鳫�B��h��u�#�z�-W��yM�2��Μ�Ɯl��'�D&�d6��ZM����s��be�X���������7I������&�P�AM�a8����l�r�����X�%�z$�JEA�\�r�����H��y"1PtzS��1�m���/�U$����h����̙�	Y�\*���"�u1�ǳ��ٹ�����@;�B���;	�0��L�ǡ�Vٍ�-�+8&��<��it]�h��3�5�����D�e8,����K���,t�	�>�N�Q�g�:a��]_�Ϳi���9�W֮�)}�hX�-�rDY!g��)�XjN��{*�{K���˴�A������}>�����G�{|�� �fθ�x@>?56�{'�n�z��]�z��I�,>���������k�-]�Y]�g0����mn�L��E�w��q	��9�m�~��IL�R����!��m�r���V�1.����gd(|dz��4R�>I��^�Zn�+L��I�P�Ъtp���Fs��?���NȺe�Dl�
�r:ܜ6ĉg����S�!�p-ROI4��\���\�C�} �xBe�t?0pI�1��t��Ⱦعz�-����w��vK��#��O�1j(�
GQ�ְ��-@�զ�����/-�������ږ��:�	 �Q��gó����ER�\��#™�ϧ����Zi�J]���6��K�-�"�͢^*�^NNd4#ߪ��
������]�$��B[n�e���cq2���y�י�G2�D8)`1�F"��l���-ܼr�xS�s�d���7�;8q�a��Wg��ރ�%�f]�uD�r��Z�o�{HHPǌE��-gE쪜�� 37�3s����Օg:��JIP��JK�,�Jt�	5a'eOE�X��#�܍�?�q-��eͳN\�k(�Un�p�;���'�ڬ����P@�2j�-�?*�j����$�)���n�K(Uv�FK $����y����Veݎ�MaN��Φ�+�+#w�6��$Z�V���}6�f)�fC�H�a�t`$��4?7}�aI3���&�@�1g�u�,��ZH.�$�je���}D�'��g@F��PR PB�Y�!��,�a����+g�[�/�Y�(��`�C(������r�Q��p�%������ٛIv^Wb�ܷ��ګ���t�  p7�8G�则���H{�K����pؿ���;&<aό4�F4%�Hq�H� [7��F�ku�KV���L�s������.��ݵd������{�=�˟U�S�ZǳsP7=(=�4��pc�Wω�"K�2M?�K��$��(.�{[��|ޅ�d��P�*j��l�@i��p��~�3��h�E�� �����i�KHdR�ii��#��/!���Ƌ�\Cߍ��ټGu�p�e��2��6_���¢H�t$w+�6�Zs�����Y|�ߠ!�'J�iޝ�s�;(5l���&C+�i~f���Z��1gOe)ə�H�*E\��)nYg�M�T�q`�%G|��䪈�O$�5K�<CC����d��t�6�9��#���R�{$��c_��}e� qaG���1#$:u#M�$
ߕ��% 3�><X4�Ԁ�tsh �E$&��	2���J�������xj�#�R���dz�b�횔!�T�����W��Z��p���M|�x�2yj������"#��/ g�g�F����M�,ns����u	�M6���H���_o���ִ�,Cb9�l:E�e�+���)���
6�2�:�ں�j԰q�7�V��o���ʵ)�m��a1C��A�{T�B7V�\�-C�'��ȥ*���#n���N7ҕ��p�<�D��]��z��n��0�V��U�����FĕU�����lE���l�mԚ��5:O'i^	�i �k`qk���/��|G��Y��ͨ?�uc�<uqWh��pb��@-����&��w��'2��B�T�m����'��K������@�`R���ӌ�_���I^W��e���qZ7u`{K�B�L��u�S�7�x�qj{m�Vů=��Ku�1l@O1��&m��[k(Z&���{�������|�j�槔w����NrP�޺�r��//��r,��ֶu]gy���X癜h4Q'�����}:���"���p�����+㐣�G�f�����?�������^�����g�2��3�f���~�4^6�fP���[��_���a�`na~�eG�V��"�;��/~C>?�w�QiZ�yp����-��������{)1�j#;[Ā{W�>��������)5 5hc��*���V{����O��x����Q��8(q�?�������I*ɋ
"`��,��ut�<��E?��_`��-��vhg
++X9v� o����������6�������Y<��3X�s��E����;�|%xo���d�3gN���� ���Z��Γ���5�jyV����q��C���qj��lf	��	�<����C|�7~���m��;`�ɀ�΍�a���?��{�!���Atd��O���_�Hfb�T�$�Q���~����������g�awo��$���Z	s�)|����
3Ks�N Z3`�^�;��s���w�����0�ux�]�1zM�3ft�~���(Pu�<Ep��a0z���=?TH=�M� �Uއ��}�ؐc��4���#�y̴S#�͝��)І��߿!ڎ�:<`鸍s��QFaç.X�~�jMD�u���,�_�S3���/ХGz.��t""h���W��Y'�~���~Ϫ�v���ԇ��Y���4�w}�|��~;[��LH���S���҆��[�3I�I�Qt ���8���Z�V���1���Oeh/�^X]����C>!~��/y#(:Ê���f;����f���1�qj3�[��NUC�&n�A��$Ge:�$A�YC!R�^��ԝi❁%��F\����T�x-"�:��qLf�9�9+[���s'{LY ���E�����LZ��5'�t5V&�������4�tm�X���bM:�&#��$l��xf�ǟo0`�Ӊ��1�Ė���m�j���W�f��a����"�q��)9�#^K�4�"�iT�����h6�4�!mͷA���	���K��X��	�v����'�B�E�4ΩXƒ�AGWN��& O�g��C��I��X�zϞ�Vi�|�"��q�H��갊 �q��l?�Ɯ=e[��V�C�2�V>�\F&d!��M@��ȿo0�v��IuAz) ^��y5ݶl��AL'� N��&�&	F�Ey����`&R�y�xu4��U�6�b`ڃj��\�&��&��7R�P��Ou����q����*	i|���R2WVZ66�I3Z����C���PÇ9-��4�1Vjw�Q�(p��e��]j�����LnDل�F4���\�tr���8ɕ�uގl���IF��Tb93�FJ�͉Kg��K�	=a$O�(T����.���֑[��^��_�~�*v	䞟>���"o���bCSgj���wU��i��l| �s�W���]�	8c���.T��r�*vWW�����Oaz����$P�����
c��������]|n��_z��׿�{\�l^?����N�{i��[�2._{�4�TPc��O[�ʩ#��;?�7��Er��{��p~�5E)��(e�[���13=gN�����'ܴ>뭃-s�#�8��g��ѧQ��t]W�x�"���j5\�x� �C��U61��N:
���&���o�K����*~��Y����E3��݋��uj�E�J� �isH[HO�0}h���e�l�K��B3vs��Ә�]�f�|5I��wxO�|
�����ˠ#5̣�5��멫�ڬ���o���oo�N;�Jd����*��`W3Ny�wK{��l�T�X������@]���qi�� �,�T$e�C�46P6j};���L������&����ޑ���g��������]�C�s_*�&�S	�:{{�����L'ѧ]nD�E��%�=���Jo��.^�³X(�YF,03�����g���x��u��=~�цZ�&j�!��.��������'��ghԚ0�+����_���ui'�����;���#�e��mq����\P`�$ef�{%p�X}W	Y�,���MFL �k�#��m�^�����?I1�*G&�ټ��m� ʟO��n�NF�5���bȅA�H���,z�	�G�8�]���F�����G��E�RFb�J�ְ�;e�]��@�,�ʛ�g6�#���Y�*l(ᣤ��M�*O#����h��U��s��8��з�m�v�@�d~
�u�jU��R��;�q����Jw�4}��/Z��f��Q��Tv���<�͖�KܯP�+0n��k@�s��c�6������|+�ױw�:����� ���s��������U�n]CnzO=�e4y�������-��I�2RN0rV�vD�!�c�����6P�����j>L��#@��X�,�&��7K�l3��+Θ")�C�DO8>���R�ܥt�xhG�������7V}$�	�_SV!��2.�K��q#Z�ú}��%�kzx��5M�p�@��1f�4�D�:X}8��
�� �Z�,�R�� %�F�'j�@C�&~ƥ:�����С�4&�ց��4-X6�e^���2���K�6E����Ìv<ܺr��`��e�	���<pF����y�qL-,���z��4����|G7��[��V�}n�8�Ç�x�C��~ч.�3�;2�"�8�|�f�l@$C ��͕*�D3t ]�N�e =�fWs�~�m�;]�o��YWYQ7���>����+񬁿��4c�<nL�u�{���O�O��T���A?a<*/p]�~׷x0p�����)�K�EY{R�D��Yrk����5'hL�6ME�!���u���E⽁�w�{*c���$?n�|F��F��"���K�-�P*8�[��ص�lz�c*5��HxvoJ�)VQ T�8�r�<����F���~��q|vEu|��!�3��$�I+��7�����D�1[�~�p>����>29��6(mT�7����6�-��V��,��nt5�sř%�v֑i�F�:������/�}�|&�x����a�!��h�{�|�6���%����`g$��h�p��M\\[E��$�g��_đ#�q���z��7��4ku�g=q�Q�fp����+��������hK%>ݰ���4�����޻}�
>�ܳ�*Lbz�h���
�\�ɟ~?����މX�, G��j���A=�W���Wo��S�"*�|; ���͵{���^��\�ӳ6?V�ʤ~�ѭo����*�g�sR���[��+?�A`�l�·���|�FMV���wʛ�g�s{�9oܽ���K��H�y��jOk�c@[�������$A�1�VW�{{��&����!�^��><�_�#��Gָ&[X�)�\/1 �Xg���P2:Q��s��(ï���Y��:uZ"�<�=��G�����$�`kw�2l�};�n"C������;�ڿ�7�|��z��\H����an�
SӦ����w�*�2���:�%Ϝ�XA�29�L��"�徘��՛6CSFVo���w/���d����qm$И7i�J�L�%ʐi�|�i�:�.�59��t���Q h���}���a�ldhg�X�j�B�OS�ĭ��~�Lz���L�l�x����'���u��^\��4=����Qж��v�v��/�����D����<qI��3p�Ɂ7��Y�:L&x���ݒ~�s��q�q���G�v��@@���䟢�(#���>�$��%��ӑ�r5�h $�]g��!ȓx�F�i�7�yN�����D������Z.�I�y��?l�D���kBӸo�����L��V]��T�+C�w��ڮc��=Lݮ#ï�6jD�-�^|7�`r�
7/»v��S����0T#=�2�*�lC �<0)�N���m�&���h��ӿآ�m�����o�ΘE|����(j��	�l|���=��6,��D��}q����A�QG[ޖP�Џ���0m�j�o���%��0�	'S��HS�����$t�RG�,��I�Di����*��Պ�_�O�t2t4�F3A�hu�N�ƢVE��l� �k�,W3��D'pCT�t~&�gX7͛#�w|�ձ�7���>�lf��-��n���'q��gP���N�6�$�9&�����-����������>��o�1��s{�#��������=^���I��1��%}tJ��� `���k�Ď�|������-��82�����Fc�(ό�:[�p��3_��S�Q�Ɯ����t�
���B��P~�7 6�n�3�A`��xʕo}M��(�f?�فm�-Gg;TGt�79뾦7m�f4����wS�������F�	#�M��-���I��/�A^K$⌚"�^�5i�z�-:Ǫ�\��EK���ь�� E���T�{O�a~>�Gx����P�1�\�k֭�4a��	�Zm��hMAp�Yt��I�D~��[��푮Q�e����������+(n'���ϱ����>X�G�9|,�a�y/�,#s���W��ME�єu���pd�pd�=��:�,0���ޕ���7����E��#H&V4�=,^����ӏ�'����XXx�������i��E��������h�7n�c}�jb�Nj@/Jdm'�o%P}�o�@{�y�"6U�mҹ�<��.����=�����ѣ�&�l�TJ-�7Ρ�l��poV��e|����;{I������������C%t
��)�DTN�k]��J�&�Gj��'�CtT�rj^��ϡ���P���#�
�����L�R�7��m�Ku�)42x�5	�x�����t�}(5�N�lG�
h�U��6��Kͻ���}�w�b:ZD+���	k�/ѧh}'���f��>��m5PШM�VӤ���x[c4sd��;��إ}�����	Ln3ϊF�%��NL�����7~��B���k�N�3~� ���x��s�c��h��Ȧ�ػx���`kmS����94K5��׾�3^�4c�V� ��?���G��v��A��A.Ag��uܾq�Ϫ����.x�E�~hj�jF3�TE�눺r��	j�.HѶ);�V�Eܳ��bwM�xO%с��6����H�)���S#�J�)�1����4�*a���w�qq��z��i`XN�p������o���mҖ3H���z`�p����-��y��G�PP����b���pjP����!���i����dէ�w_�_�)?����y�Y��[uw�]{��@W�hN�?/��.�(��{��G�QCnF��`$��-F�oR\C+��?E�3�������aة��R��� O7�Te}#����ax ���qw��Gq��_���n{g��L~
F���>Ʀ��4���E�	��H�j��6n�q-�2_C��Ym]Rɔe���7�<�J���"��g�l u�F�D�?��F��H�R���;������9^���	�ꊔO�Y,9E�$�k�H�|I��\�G'p3󂈥��È�W�ä%t_jD�p ��ʴ�|ԥ�d�:	3�it��A�n�Ə筜ӡí<w]F�E(�qx�(���Ф�H�42Jk�mc��W'd"�C���E�Z]Ed{^��j�x_�{��� ��U#r�tj��M|���9؆��<�����ÝJ��YH�˨��g0t�%0�Ӱ{�H'
h�e��1L���Y��+ȧg��#s�1ϵ�����C���!�܌�2qN9�P�XB��D�R�hI��8�W�V?7Ҭ_Fh�f�ȹ�ê�K��Xy�{Q�RC�Ӟ�幏R<2U�M@V�%�j]oy�6�e?Dl������Cߍ!�6�.E)�@��$�caL��~��=RwZ0�>4��W��7
g�=��1�X�:��q���-��t�5o��=�7��?����eǻ<�
�"Ꮀ.c�~�ư:���'�&N��u_��ndL�����JE�xj�4����E�����~����E�`i���K��8�ni�&>yd�G����� �Q׺��2MR����xC7�S�!'80��ξ�*���l���t�qL0H|��Gq�3F�X��6[0Q(��*���E��	�J�pk��'�"RǬ�u�<�qH�F�Bs�3����� ��Bt���iUsP�[]q�m���^z��{�@tݲM�~��6��[��j%L�1��l��*�1�@ah��1Gf�S�g���nOX �IM�y�v\�f�Az�{`�g�6Z^����-�/n��źz����g���x�|df
��Fgr̪F.?Lྰ����LN�2r��e�7P��C��À�i���W���|���EL�RF���2X*�&�:�`2�(�6׷QAG ]�I���CS�t�l�e�4ƍQcL<_�N�<�?s�*��}��JO�⥩i�w�6&y*4'�E�����n�lC*>��i���s���0�@�{�Z�HΞe�U0�u��)4�4��_�ER�Wo�i��5<��c�ڱы��|�U��F߄�}�`t�7T��*[	\�JO�d+����36y�?3���K��fg�Y�Dh�c�ُ�(&�D0�V�?���{�-MR���r,p3t�������KJL�K_
���ɱaݸo	�r��r����=7X5��5���mI.i�]��f�p��|���*z=GkIEcf���Jؖ���UTңoY��#�|�JU�l5���fG���N��� V��z-w}#���6�Ab�H�%&�P�Ev�������-��9���M��j��]k��)"ۯ�1r�*���8�v���Ϯ���Ӹ�~Ә�dv6�C��E^m�r8�i*�aq�f�kB�1�r*u�ۖp+7G-9�9��D� (a�r�Á�u&1�s!�랕�� f���Ж���AV˻�u���t"Œ�`�`�W8%~/\7�׍*2�7D�	�j�)�<�K�������)#�IT�5��<_+� ���-�׷����%�e\��"�a�M�ǧ��بE��BJ�3^l>W@1���CF���9Fr�*:u��L��Z*��F��E,u�ܢѻ���QY�#�TuUsc%��&e�"�DL(�9�>,�<#�ȷ�P#ij��e�J�G��C6n���e��4��L�����|�33E�]>�.���)�P������=?�#(B��o):H+Q�\]��r���1h�~�N0�(_�9;e��q�>�r3��!��}e䘒���#iF�j�D�ٵ}��X$,]y=�8���Lԣ�hL�/�2޵B=*j�PĭL^��=g@Њ8��(X��:��s$����,^�(/qV���c��F�E��j��.x��+·L
ҕm�e�t�ڢC��T��%M/sW|\�����|���e�=>�Lɠ�!�xF*9t��P*I4�[Ð�c	��Ġ���Ր��������>'������{��D�� %�V�"�<��):��|iz���{�/�]ڲ֠ɳ���������6�8��1xr��7&��VM	zӘ�t{ؽqW���K�-#�ֹ*����ɹ)kx�*tP6 �SI���|�����ҡp�w���~
���8{�,ο�>�mK��i��֖z^���F��H��1�@@Aг��g���Oc~qW�v1��&�H3�n�vh$c4�[���-��jXf�m/�}S<���:�}=�U� jd�.m�g�8�vݸ��ЯNGMz�U��hƷ�3�:�Źg	d�=.�cIzZ1�DQ��fP���0X�/�����6�F4�t"�:���r�\C�*3�f�Q�<���Y��<ML\�m�[B��-3�T&��r����Y�C	d3�HH�!OR9�ɴMW�w�VK�d`�L����|�K��A�_TПH����v�2n��]�)���G��813�~�F����Dָ�C��F��=�1.�xߵ߃�N��@�0�~�!�P)�a�k���n��OÍ�0z1��Z��Ѷm��P_�=1(�,�,����C��Ą�)���d����\�q����T�cpR���$�0t���h���LDq�v�+���h*�)��������VS�ݗ�8��N^2�����G��o�yh�]�����U��O��T� �濏�q��e��4�
�:�Ǎ��I=+�<.�+�6��\h�Z3sY�Zn����.2���3�"��� �}��==�4XQ�3y��%�n��t�D��xfwG�+q \�����ģ�}� _;�vG`з��Yy��?��-ݵڄ�PԈ�Tdԓr=����T��^��n��>�O���i�����*<tt��E��Sw��R�7Gcij���K�0R)��0���S�B}�D�9O�s�SNhѲ�\iƩVc���M�ʥ��YM����:�2�E�Q�2G{h��,"��^ԗ�\t`�cu��q&�Z����!o�A	���X�X��k7M�MeMP�b�'m=���e�\�����Ǩ�hw-tz��U��	hh��܈��qW�h�(7�x3"�\�[׮�εk(LMa2�����m䳳�ISY�T���[����?�\�n܆hGm�C�\q�{�V����H���لak"����V|E�ﰵ*X�v��l���Av�&����ƪ���1�sE����saf2��jY��_�gtZBC�ec"+��/�d��9���=�g��B]�y���ʆI�M���!ek�-�<i4X4�5�$'#��.��X�s��އ�V�~m'Hv䚨.ܿU���?3s�aq%��չ�?�&,�x3��Nn��c����^�����J��,=�FN���*����kK���w��)u���#7��B�ƛ�'�u�+S�нf9##FG,:
G��2�H��`�@߳�d��X�>��u���Hq"��-/�Bl��fɉi���Ϸ��t(��V��r'�)|i�(��4�0x�<M�J�,m�v��1䧧�����?�GN���y��kNQ��Jp�;��bBǚNR+�\��?��_� s,�zY��s\$��,I��*�MM��l�\+[S���q�(v�"�m�P�����6R�<�H�f����ԙ38�ԓX^>�R���簵����h� ������2��u��A>�̙^`�\D);����)������rQ�*��g��wC!�P�UB��y֢Q�~4?������#I�������7�Y4�	N��r�(N�z��eܺ}�lPqfބ��F����-`��U�;�t���j�,�)c~:�$����+r����Le���;[ƥ:�*bv*��+KXk�%Ȯ���}t�C��fJ?,�����%��	��S�	|��p)pc{��~`��J����|��ճR�����:ڃ���<��4��J��
��:����u:�_��mI;�5M#�΍�?�(&Մ!��\�#P���+"O�3�9~{�=��.j%��h��Q��+�����n�@,l<P�)j�����g��u���nБ�Q#���4b�ͷL�T*<�k���_V��g@2��}T���$�|�/N�?t�#��	��tD�U��[N<b�'�+���1�������B^��=�@�͉�k���V����>L�M���������;���|�bs�.�4Q�d�֖��jm�d�ռ�,�}����]U���u /�9�2z~��C�_�l�o�Z�̌�8ñ��/��� o�
m��u�t�rʮ)�A�U�Fɫ��.��e=�Ա��)�=�It6����9Dr<��>����q�d��I����4Q�FCS�#�#�h.�Qv]F"u�x��F�����g��3.IZ�XL���Z��Icn�F��q2�7 �|��͵m���*]LM/�M�K�n��d��G|�:N["z\&TD΁7z�&.'����$�2r�ﺃ���3>zl��@ �b(NV4b�<a�l�bj������*�zM:�v�9?S�Ѹ�|f���^��FI�2��Z�|���ˌ���Ap�8�2K��e�����>���U6�`�@��s�ꄢ:�F,b�-���Õ!T�s ��x��/&b-� ���VZ���-���'�Ȝ�r�}{|�5L�Oڌ٨��4�~�YԹ�,`��GC�ܳ��>��ݸaWRU�ʀB�q"�
��i�,Q�t��.�������Pl#�J^$:�L��чo�'���Q7�V{@�o��TӇ��q����H�Ǎ��퓈�]���CK���Hڒ����ܯ���'����IE�H�����'�A4�TorV<[[��ϒ�J�Ƨ��3u��]��A<�F#��HټE�+���t��eܠ�b��9NOG�R/x`��x��րjO�/�l�r�2�y���V��(�/�WFj��w��6~Nk�6�s��U|aj���'速�-��O�5t��Q��@R�Ȳ9��9��t��KԲK]Dk|���[8W��D'\(�19=��wL��đ�hη��j��M�7��4m�N���7VqW�kI��߅Lւ\��i�~�d���l}5�i<:1��z_|��X�_ƍ����Y��W�ߧ�IMX�?���,���#B�������<��0����`����#p�|��@�۟^I޴$���e|�K���i\�v߽�F{{�;r<aǥ�[����CmP�����~u�8>=�}�:��m��޺�u�v�R�3-cff
�'��^�ٱ��x� �>|���_�\���ş�5�jy�����=IX%o`پx<�6�W�s`�:H��x���ON~��̠�-���-��*�'���](���,ډ�GCΙ�/Y�S�I|l��B2�o�w�/W��:��F;��Q��ٗl��?i 괽�<޺{��_:|
���3Hs^*o���K�P[%�-�M��̥�f�3ƽ��ihҔM\a�����&P��M ! �Wa0��"��q�M\*�T@0�ADI�������Y�r:Ee�-Ol�?s#h��@�g��s[�f�+
Z�a����Ȫ�vy.��k:�bsˋhml;���Ys�в�J�hx�]����v��xKe����4@p���!I£�L�9Wh�g��Ƅ�U2�w|D�gx�a��^�5Z(��ďǖȺ��-�sȳ�)+(k�.�f��+���N�*���A���Vi�!�%�,c�𼐕�d^d�<E���-vS,�z���QuƷ�����3���L��D,� �!l�U�[z?|0�yz��,�D��;�~?���:<~[7޳v�>AFmw��Zk�F���%�h�E$r�ܔm$��	���>�/�a�v%���0�R��#���8�q"��%��ș"^��)=��K�FíA�S���j!�K76��n�s�ԓ��K�n�E'����&m�NH���Y��\J�X'Q(�R�6N̋Y���SQ���D�
���Z�_Dܰ摵}k����1���M#�N�WD�v$p��rp}ל�qkʤI�O��"t&��kh��s�t�6y#袰2��<i_�ޅw�6���a:h����0�2��o�|�e�}?���ڵ]����[C������E{C�GÒX����3��Y%�P�<���gPx�Y�������V��1@,)�陬E@��x'q�v�N,����0���0"�4��6Ǳk�{�h���� �nV��lY�.�LԤG�nz���0�.[���ךrb����'0q{F�69ʀ�W@�>C�M����_�j6��w�ߢ��Y'-�fcާ],�#Б�e��t?�.��:r����j�Q,c<>�!XW�����$��$����dh�6,�e|6���ɹ�dpԸ�[��"�D�{�����-��,�����wi\���*QD�p}���r�Vr��c��m�31R�q�ګ{ۘa��ٹCX�W�e�jOJ{)\!����fq���[;` U�9���֩B[��kee��GЮ�M�!Y�ZVK�>>G$�׿�G��_������wp��-����d�&�>�x��,�k[����}%n�Bq��'p��y\�q�ʹKG���H�֝��5{�5�)�������Ɂ�1�ˡo�(��O=������S�ɠ��g?�o��`��5<�p�?�GFi�&cm����l{�w��:�}7���ٵ]�

�j�`�9�½-��˙�5)��W \%+�#�wqA�p�f,�	�=ڮCU�B�>#�Z���Z�f�4y��u�ުuWJU���?2���� �{�ܪʎ�;��]g��Fr�5�$����gȘi�F-ۃVg
�x,����<z�%�ݾ
�*�E���S���vO#�#���)����s3h��7���T��3@�����N㹧���W?���7l��>�	��u���/�R�BGM�q�,k��=��D�|�q�iD��؈/���k��y���>](�0�
���TP9L�͖D�ufdz���d%r_븉F�#��6M���4��	����5Ag�����kLp O����Z����q�}�]��S��	58��OQwxDZ�Qe��N�O���l��h�z��s7�l!�dVB����ժ(v��|%��5�g�o�6\��)�:�@�d��T�ߔR�&V<�t)qb63� ]��裳�i'zU,�a~~�{�nF�?��;}��������+�r��9�� >1p͆q���2��6��a����n���u��1P�-1�i{���ɨ���1��B�7��P�3�>�&��7h�.Q=��ʝ���i�|%��z	����;���-�h�J�~{���.��6�:��	�G��Jo���9���}��w# �����Fp�����{풍E�8��u�[{x�h��?:��=}�����]A�����g2>�z&�O�8�y���O��K+����8uQ��/qW9�XF�94x��4~�iA�������<�Xؗ6��c����+�n�����z�a/h���2�u�I�%�x�o��٬f�7=��h��B�,>M*�D�Q|f;��n�(r,1����.әL0��G�N����s�~�;8Y�gd��N[���f�~q���-c)��HF۵�����C�Ī��	��#M:�S"�$+����2�6f0��f�\q��o�G�7.�KC�G�ϱլ��b�X`��Lv�F��K\��-�V��	��4����e��L�=��h��0�ce�x�F!�6F,f���v�Q(j`R����6|�hOzuC�����J�ȩA@��8zg�4�U��WYL�!��qU�?"�˩��8p*�����0�2rR1�Rf1�:�x�����L���`Y�����N'p��]+�+$�1�tj���u�+�U�@+u?��5�U{�:Ö�s��y�A�e����D�VR�K�>��	>��fFV&^>�u�c�0d��k�6�]9��̾Jq�t�B�!��A�Z���mL���]:�W���jP��e`o���7k�qjj�f&�4��Ր�$��L6�С�F8���3Q3�˛������'�}��9Y�qw����{o���+8~�$�A
���ݠ��7/ᓩ|%��7�������ҩK����Ϝy��ӡ���5<�����m���E����+��j!39M�X`y�����?��t��ۿ�S�N����6�u�|7z���U�@�\9����f���+5�HXV�uӪ��y���-Бq��E��.�q~m4�*��#�i����iF�ѫc��Z�ٕ��D������]��b<{Vo#�} ^nOg�����!�2^x�v6��px��6���[x����k-�}W������V�����X׺�;:\��{!��G�E�����B�7z�N�R�����j��Qejq"�lx�sٔ�~+܍mο��}���x���(YS����+x��e�8�8rS�V��ܪ����H�H/D��{x��m�����+|&S�Ԥ���G6�F��na�A�b�����8��:��ȥ2&ꯤ@��,��7�#���l�5�lv
��|3]5\)�6rd���:�#	um��'&����^<�<A�`�d	ӗ�\�`_�5p�(Y� @�g�S8w
E�}F�`�$�B��m���V���u�:k�^�/5r��Mqa�ó����elܽg�VڗYY�5�si�46��G�f�Nc�,�M;�9u�FURV�W$�s�.ܫY�7�f`�T)0?��.ab�{n�AcņL�˘^��­��q:����h�p+��A�����6�s�r��6Z6ũ����^=SC�Xb."[I�9`>a�)hW�d"�v3�EEO������#��㴺�96�|�C+h��!6GS�%:/2*+N��<���*ܸ���67�AN$[@�{�b~SK�,���Fu��q�@���f�&U7g�:�ĥ�Y����@b�kXA��u��"�y�����E����AG𱏜����7��k�p�}D�����/`2�����e��r��sF �T�H� uh ��B�{E��e��7�t��K\8�E�{�Q{�Q�K
�}��u嚑'�%�h5���4�EC>��%�箬�f׍a�ɖ�q�����	<G#"�G���j�h��lB��E��~�����is������c��mL�=z��h����p�����s{vj w ���#�X�Í�cNZ��T�53z�0��ݯ~K%5=�4�@"��v�-�}�.\:�z�lr�z{�8�hI#�TR��{�A���h��oU���v������"`��y`�6mŀ,���J�q5��+ъ�9t`W�6>�ϯR�8c/��r�J�V��݀�V�ې�m,B��՞+�B.��DFe�DP��� +�Z;=\dJz�V����m��u��Y񠤭&�[��Z�.���'q���*�C�����ǿ?^��,����A�U.!,�����W��i���R����% <�����ʚ�ṹ�x��y�@&A��b@��)�-#TB�x<��.�����qC�xF�Xld���=�i���m��Q�ӹ�vI�)�x�7[k�qm��8�sLRڿH�[�=*�b���u��V�=�V��\<o����0@�բ�>v�8���P/Uq��؟���x�՟���������lO�Ag�$���+�F�����'����Z��˖�Q3L����3���t�J�R7�XC���Y��r��A���έ���q��i{=��K�8�yyy�
z���6�+HЦ��n���g\_i�A�5I���?�1u��V�i��1e�+�E{n�z<n�<�OB遺C\ڄ��3����K�>�TK�Ө2POb&3 ���c
��lE��i�������7�s�.lmિe���֡�j�����&LnJ�J��I]�1ޓ��h�"{5,�	v>h���'��g�8���F-��k����L��w�<�Q��,��6:���%􁚪�	�	~��V���_��~.�7�X:�4	����>���g5��ח�>S@�N[�i
���o�\��l�������ެ�hG(��g��j,�Uv�@�ߟ����J}:E}g��1k��yÚ�3�mR����j�j��k�|㦋1�Z��(�p���3�WCb?���6w-,N�ϧP������p��*�6��C�1;���̼����Mx��ה�D6m�sr@�^�j��J�h�I�_��-M0��\��s��T�"�N�Q��E��Kp:��M(j�����oW�����!����4	��֐p?��Y�N��
�jx�)ڀ/g �'(�#�IP{���N	{wʘ��+�#��fP�@���s�W�%����w���������/yNMy����G���ztK��AU�/�FTq��C�ï����n��]�2��`��N����j�N��d
��ک6�i�Ա��Mu	�##B�����s��eR��_���8I�؀�������G�d4>�Z��>}�<2G���4��)F�g���cX�a6=��?y�Z����C�x������l>hߨ�vč#�M��S�D$�Aρ��[M$��%�������5#4j�AC��j}���s�=�a�H�C'^���znJ�Ȏ��b)r���[��AgPƨ��_	L�H*�]]�$Y���AK�+���_������z��7e5�/$ШY���$ت�ZE46�ٺ�{&Y�ڋ�v��mD���ʂ�c7칒������Okq��)�������{-��fKRhh3�Z�!�VG�X>:C��3��$�σx�@��A��g�A����A��X��1c=ǉ0I:=����-���U\T���ʪ�r���>Ml4�f_5&M:I�I<��o�PǷ�w-�������iq�<"#K	_@�5��.�q ǌ���'�Z���~w�u�k���P�f8S7nJ���Tڇ9[�]紛�2��Qv�U�1�8��1[4���2��h�:�2tV~����Jx�_1F`j�hx�G2�tqSʨ6��9�K(ӹ^-oc[��3��N:�H�nʚ1�Jׇ��H������:hg�Hu;x|�ziګ�U|�}ԣ3��u6����O�]ڗq+NK|u`ߋ��a�l�i]��+���UQ֨l"�[��_\�j���G�ane�:���I��&mA��(�Ev���,fq8[ē�G�S^�mJ��N>�m_;��&{��zxyW�\Cf"�T,�r�i�y�c-��y�>�Źy,-.�S��N?�8��� �._�s�>���|����(Й��NP��i[�t�F�yH�[�w��$c���5���������,��C(_�����Ӧd��^7��n��Q9T|W �&=O*=jr���2J�>R	�m:��[F��C���w߳��ޯ���޻|�o�����)=v�[��^_�d.c���J�ٰI7�͏��|��GYp��Z1�s3݋zx���\��A��)���f�J��d�F��I���y"�G�몮�hv�k!�E����E���(b��:7Q�M뛠�}܋���w�_�MNZ����~[sr{6͚y����L<i�+���d�:I�M�0Jψ��*�5�H���N:��I�Dfp�Uh��R��H����V�LF�^�&%Av����' R@�������p�X8�v�Y��Ȧ����d�{�q�u¼Qצe�A�?�zP��":?���<&/[�����{���y=�j%���i�9ڳ�iMS?�b򳴭)�k��@M7�[��{7Λ�����ۘ��r�eGO=�|>�{�\��$��V�?H ���g�Hx�&	S��s9�f�ƒ��
�z�,/���6�����x�ӓ�]�x����fv:(�눴��P"&�͌.H��[���a�T���I������|�`��\)��?�&f6n�S����>��6:o���s3�`�ڻ���h��QtS�g�h�Ҩ��J[<2 ��y)+�Ʉ'y@
�3&G��+��r�`n�`��K���T�Hrmn܃�mT�+������y�*���I<��G�]�ݫ`q�q<y��x�7x����?a��g?}���\�r�;9u�2O���(��ٻ�����"*u�F2Q�+�7�#�.[e:�� IXi�g��TYˣ��0"�������h���~�&�0��u��etW�̅�T��F�=����}��5���tnd���]����X(m`��}"�h�9.�s���m��_�������Aw��C��8�bA�]y�Iu��qf��{��חӞ�䭫��=�L%��AP��Dtg"aY���{S4��n�8-��	���9ퟜ�EA�lڲ���=��	���<�1S����%��S�{�������H�R� ��1]<����Nq~��!c!��83!����Q�X��7p�Y�@٪���������F�:o�K�(#���`���Db�a�S�n58Pig�v�zn�f[Ż��OP{�K�?��Np������z��������"j�jfn	�� _���u�y	����xx���	u�6���fV��M��׺;t^):c�9:h�(zs�0̃,r����&��yS4�5����A&�t������=n^�^�`
:1�:�-#���*�n�QZC���Q��~�o�
^��Q�ܰ��h[����K8��Y���<y�L���w��)$l&j��^,���q���7l�y*7��ڽ5ܸv�J�O?��e�:W��u�֥6��>�ܳ6k������I�H�03�����~�:������mℂ�.�qog�G���/��o~�[|���y�s�ݬ�h2�8A���i:v�}�L�	z6���9���ŨYFk��j�������t.��騝�h��`ߺ!���{�3���K��K7��W~��Η2x����{Vb�~�&��k����R�+Y0Q�q����;��_� ߸s~!KP�F�ǀpr�2�����@�.e��7��2}���=��sշ���
���Jj�`�`��J���L4_]<��ۍ�M��^��o��w.��W^��yR��֣�?��i�~��7Q$P�i-��}->��̯����[���[|>mTh�s�H����2(�CWɀ�I3q��7�\%���|��!���ц�Q�'�$ '��&8&Ҫ���(��@צބ:�ք���o�|�����$m֠묂�,���)N�ںV��XW�ѓ"��T"e�`0��]�g��$x:���G%��B���͵���~�Aφ���Դ��10e`��m��뺎~��_'�+؜beoe���l�Y�(0�t�X�?�kd\��G�ì�,�N�K/|�\���/0T�|�`{�����#�$]��ϖoJ>m�d.����}��O�������"�D�~sŹSXz�0�G"k|�����ƐޮqҞ������:F�[Y�u�s8.s��Q��:e�����}��LzaX*|JB��na��%�(�f�l����&-�{:��D�):�{�
*�.z�=�[+���ǱZ���z�ѣH������ˑ*��f���?���m<�՛wLp�ʝ]|p�.��Tj-Ԫ�e�"����UTwv���<6+������/�pW�o�ݷ��_^Ba���Ʈ�;N��0y������o�dwV�hT���^��jb���_:D�6�.#�^��Q�f��5s.�姀�d����h��tK��QqNusO�K�mb�&}"�'��a����w�-dd$A�4�fa�i�R�uVʵҁ���N����@��(��u��h�2���V��}�02���1��D<��f	�x�r����ږn�qK��hT:�����g#�wM]@�w-�Kޤ�h�Zh���8�%�V�������=���4����H�8��[�@�z"��O��3k2꼱�gB�U��ۥQ��WТ{=���F&IN�Q��~tm'fS!�N���L.��  �����<��(�2��ϝ-?ԝ�x膀ˀ������.m���.dߜ���֕<r���S�>k��9?��Yf�{�M�٩&��O��i�v�a�SqUɷ���� �Eq������V2O%kӑ�B��Op�Ƶ^���q~Դ���[t\+|�3��贊Խ�>�l��yԓi����W�[��g*�n�"�~��m������d�Q��N����ʲ�ǖ���a=�c�RŐ���ﯵ�n�iY��`2s��n�����$ ɳ�Arе5��>�t_���{e�w�:��|&���)�?{��E\�."I�8��X�Sk"Mpr��s�~�����7j�����D�՛װO�vo����to�/_���R�ʒ�	<��_s��0Ą����X߸�z����۳_��bii�dU6	��2�*������_������F,.�g~����a�@\%B�G�e��WZ5T�l���a��c��	���{���==;�����[���N9]0�٘��<�D+�%����uX9�8��r��:�)A��\�$�魽X�3M�"A���g�?I����$�QUI�R;tr%����2�����O������\�4��9���6��M���W�㷮!R�a��It^�g��x:�'��?����Y����!�ծ��U��j����b��[�s9Ti�J��MMhh6������}S�������ޣ�SP)$555c Rq˔�X:~/��E��,oҍ�w�C?��ao�W_��?{����r|�@p�g�A�`#�=ު5��Y���{',��l�u�z�!�Y7~�xh:��EJ�Jv���MzMy�-#&� �3i�Y�2��y�͋����Gjp��v��5�LH���q51g>��O~-���W.c��$F-Oˋhf�v}l3��>�uv�)Ĕ�c �Nd,�Xc��8d�$+��f�[9l���g'755e�G��mq�xm��<Y�cA"��GM/5` �gV�3;<Og�]�)1%v���O����÷��؋���j���*����Ϳ���zo���=|�����ƫ�k�䵜H��|f��{H�l"ҪrD���&�"J�f���d�l����d#����ڇ?�䅍|	�hr�'��F�H9)��Hse��N2
f��+�=��AJ|��E���ւ��#ǹ�S�b�;�2�.��*V׶q��U����{I�v�xE3�B�J��Z/٢>�h�3 �.Y��g�����db�u�;��x�'��r�����N�'��Υp���x���X��4̮u�0��/ �@�A:R)��ՉkP�9�t*b�o�!U�Y#��I*�l(�l�b����{6�9��AK2,#�}'���kE�<'cc�"a��6�E�PƟ��\�jrg�V��4�m��Lj�Y�������R�^0��ⰻz��B�1��:��!GCoӹ/��YL��i0�o6�Ѓ���Dw]�Q%�z[cl�NҨmlma�T�w�.�qhҧ�a�N����굻�S8��f4'¾9�Df���>?��WQ�Զٌ#��*�k�XϤa�y�u�3��{&*���/�f�*?W����5��uc��0e af1��Tt�ш5��eLG�?�Ĵ���@��F�Ӡ��2M Y�M?�=d�S�]�f4wx�5:�^�Y�CDe����
����VĭSVq<�q@G�$Ȼޭ����Q�J�`�%���&8I`�A�G�#I���_���M��_E��oJf��#��tONP��Zo��3ϻ=Fy��Y�Q��ڧs�=���cPn0�H�s�I6D vh�m� 3֚� $�8d[8.K��7�]��李x�b�;r��,����H�b�����%9ﵵ\�xg߾�6�Z�N�:A�v�*m�1(+��`u���8�wʆ���0=3e�#�A����ѥ'����-:���F$Vm�Jw��G�{�fЩtQm�pPo�mTb��<&0�|+�=E a��3n����s	�=�j�AW���$��\�i�+��q�O<�G������#R��Q��0�7�����goa�����f�d2�@-��R��A��gvع9��9NO΃`��@$@r���]�eY�ڒ�Y.�T�~ZN�RY�Jk+�6s�& @d�`�C��L���}sN>��nX.����4�o��}����s�t�}Ȥ�tƳ�V���������:6
u���Y)s'�� T�*��Y�2�$RX[�����B���T�Qx����J��A�֫u��H,��<�}'�B���AL�и��Վ31:5w�7��k8:2��cO���U��[ �����	SĹ�8��\�1]O<�@2������}�s��2 h����rr� ��;�J��\���x��u+ͥ���N=�$^��[(^['�ia8�CC���Qt- ���Z}=���M�3���J�0X2~�>Mq�����7�ֺ��mw��_� �A���:�ԧg�<�e�N>��')��7��y�����sYm�~��	"�?���GP�z���|�*�tTՋs==q�b��o�P�{�gCY�tƪ
�PD�d �S�PV����O�#C0��㏡S��Q��&��z�j�蓎hj��u����KE�ˠ�E��N��Ç�lC>c�<����I,ݭ����kp��6~�?����u�6	r7o㍾��	��b�Y��u���$�'3�.p-h��׮F�ںz�f��F!9T��(�P�Y�3]k$�Ǔ.�_�s��D� #aaMԶ|���!��$��w2L_�cr&UF�K�C�9��M��|��o�d.�m�Pc4�m<u����/ß�����۸v}��cJr�*��h�\�fg0I�u65�E�Re/������O�ja�uLf��{|�F��"&�	|���+�l��Û���s�������c��i�GS�r�~�:�-�S&�p�=\�X}:�r�fD�~��۹��T�t��
|�|\T�HD�}kX�k���[n9��Ǚ�3�޶ߑ������s��ĮwA��߳^"�uQO�4S5���k��w��IR=�j� ��JZL��*�fc������G�D�OͶ~=�������A�����j]j���oĶӝaSC�<�=��fu��
K�������\7���v�X�����u����i�xКtN�Z���jv�����d�����긍��Hg]j9z���Z^��V��5���p��h������������ǫ�N&�g�.>��J���O8�7�6SY��!�Gkp������@�g�a������{|�:�w�R��5�J�%�/V�0j>��]���M\~ۋ*�(p�#M�yD#�K����a��qG��tR�|*�]~<�A�P@��ne�hr�4��˭��v;�b��%i���*>�M���q$�y�L��9�����A�N�����6�5wp�� �����PQ��t��"��z3;P�`zTvF��:��TU�^������D�\�u���+�!	�'����O���t`}�%�|�q��ڎ���/�Kܯ�AA��Q��5��h4��'�a�>:���11>e�0�n��]e����N�7�8�	Y�N>�ϜFg����O<��eE6��@�.c�{o��w��r�,3׬4�4x}��穙)��T��t�2�Q�X4f�Y%���w�+wm@�S�X�H����9��;�\��#m��e����K���հ�UBI�ע�bЬ@�Nv��i>s
����ı#\��1���:��L���.��6����������C�u}��֏���J}��V��C�T�̔7����͟h?��6`iu?x�m\��΀�����^�cR�0� �������Ȋ���yfb�r��x쫟��?b���k�e��Oq�$����h���������}�32~����;����{Q�6��A��7U?ƈ��tas��2���������s��ԭ�۠��J_�2O�������J�_2�}M3�҉�n�G>��^Wh'r��<�s���D8�I% DV����5+��p�8�ĩ������F�z����� ���y�y�CX^�ƽ7^Ecm^��L�{�`�	�@���}�~�n,Q��Y�h�T"w3�,�WЙ���&��%���ác026�Z�ό�F�A��;��hs���%���� �OU���l�ru��m���#����m$3����V��\f
�8��lɇO��O=�?�����-����ВA�����W����8��C�����x��f#�c�,G����!�
��v��~���$\~	������X	,��D��C��8��8��ԳT"�A�gl|��5����~����|�:�{49:��'O �hs����{�𣟽�<#L9Aq��9i�I��o��Ip�$=,)�mZ��P
❷�+����g��go��ߨV��1.���-Ń�طg
�v�+����qIa{���~�S�SI�"V�}ꉧp��Q���|�ſ��\��D=	w��4�[j��y������%7���p�6T*�8�q^���.�&���A���-U�4�������x���!vp�Dߵ��K�J����=��J��4''ׂy�
���W�$�<�@��='.���s�v7ٮ��q�~0��bJ ����h�Lï?��I�ʍ�V��2��O��P�J�"E�z.):��h6����E*���z��"�̯ad(�<k��ע��>�䣎���Dr�����;��=௢�=�C@U�v,3��:ݏ��ݾS���:w�v&:w�E��Z����9�V}����c�0C9��M����6x�C��_���̪��e�š����ku��e`�ɺyl�4Ԥ~<���W��䦚6���5�}�����UHTT�F�)
"�yp?-��6� K���m�z��ө=52�ϺD�u���IT�)�#8x�QE�Q�8[4�c��MM�c���U�AW���<���o!Q�'��w<��������L_��r@@�Hmu��y-����U9zآ�tp�Y�tL^���Ҕ^rRM�v����oבJch|�ʴ����C������3���a|l�ʯ*i�=���B�"��0Ξy�?A�v��eѪ�
�����2`�/ŕtw�ؾ���&�|��E��9�������>+�Eh����E���=�ML����m��S�얙"�x��w�B����H6c�Ze���xU�
�Ο���V�g� Jۛc@����K��XD4�u�E�vV�w�`@mj�W����w�����ΣlB��wn?���1[7�i�TÖxݒ2+�X[\Ca��p��E=��D�{�����;��2& �'&L��p��U��Ji��/��Q�J.E`����?��Qjr����c��%K*�Qe��)ثWQ-l���0��X\���kױ� �o�6>��_�������gx��|�-��7���i�lvŭ2��� �A��;/��w��\5@��g���2k;��W��ZDFL�RA��'rw�3w�|C�{�N{�]۲޷^L|�7걔ġ(��=�ʁΖX�%X�%�s�{Nu�H���r��ʹ����f�t�о�#-_64`�����m7�g� �
��翌�G?�+�~?��o� ���6��!85���j���QV"ES��$^�l�����ԪW��㷿�M�=qwn���ͫx��s�#���Po�,tM[k�>\��
m���T�M?| 7�XO�z[�JR�,��4݋��uo�ј�9��.�M\�y�N���wvz�d_x� m�m��.������N���,���kx����!�OL��!~�.\�y>���"���tx�V�Q"�e㮏:��>
�v�^�ئ��r��� k�FB1�*;�h��Ũpl�Oca8����#��h)�0B��Hԏ������r޹��~�Jr��w�)���X�z�.�|P��)��ξ��}&�⁸���?�/~f�<�ÿ������$n�ӈ���\á}>$���_�B��o���+�ب4��(���&n/�p`l�}�=t�6iD�����o؀�8^�F�ȖZm�^1FG���D?���-H�SEQۡ�侼���|�	�+�����{ ��z��U�v�������!�m`�Ƽ2Ğ5���+eQt�a����B[�m�����&~�w:e�fÚ���E�4&Վ�L���IC��פ7:h�u!�6�6���t������P��=�v���J�Z�y�ݶ�j���r��p**M%�q�g�(�[����Rĝ���&��G,�o��z���T �h΄��1\�`�^ն2�qSl�y�әl`W��~qҗ���Պ��F��V�s�o0v��}���g��(�u?�������ݑs��n?��WN��u�w����1�@`ݲ8�׊��0�8/צ\)���C���5	�1%�@���h���-j��O"�7
#m#�&��0�EWm:�j�����M��HQ/Te�C�Эw����U\�}��~��a��ȯn`���N��W�Cg���>� ��ҥ�Hh*��9����D ���<.uK��l�[T�y'�9�g`O$m�j�����{����dJb�X�گ�h��;o�&~*���}49</��4��dǏX_Z��t��w�+6�)ڎ�2���_�QV鴔��(�m���G�c�R�KS�,�»W�mW*��ʽS�P -�щQ�ml�-!Ui#^�#}�!a��|�����w Ǔx�o`L����$G"�%�oI���X�Wӟb9Q�TT)=5�ӑ�Y�|��y�!�{��˒��Ў�L������g��	���˘�gM��qc���??�@�3�$>W�r��H�(�Q���Z�`���ps��|N�}L��x凯�ʥ;�35>G?�RK���ȷv���'5�Qg0Ѫֱo���3����T��xƲVު�9KT^� :ѭhBX��"�u�Jq*av�l���tg��q�is�<�D�u�B����X�n�K֌lه?������n�?��峏�;�ϴE*���
`W�n^��}{�P�R�	p��;��Fv/��Z*SfV����~�\v�Ri4�5��Nk�N�Ht��Τ�!X�I�����A�K���@�Bm(�P�g� ?�EW��]�����ew�;��<��n��j���rYo̙nV1��w��MB���V�p�'�9��=x�[/��w��ô-9�m����Nȋs+���=�~@���<�����}��F�܃CI���ۃ��!�}��^�����;�k�w&=��Dso_����V1ټ�`	�R�a�0[;��ihe5�nm�����
෿>���0}�&�L�~��K����b�,j��g��D�g���?�V�o8�ű��ϣ��H��ǩ�.��w�h����a�ڻϥ��~�Md��}-����K���EI"9�]M^=���R����n�#SV͚�՟�qD�#��jA���	�;��4~��Z�e�4�kx|��i�}�!Fn��|���K�D�?�L;y�T!��<2=[E����oih*��8�KZ-����^`�_��w����3�o��_ǵ�1K<ā*#������3��w����]��#�S�m3j�jF͖_K��+��EdFG,��կ~���)�����3J�"K �2vv���A�ƀ�J�Ȼx	*t|j]�F�!t��Ue���m@�? |�Y��\�Ӑ���0�T7 � g �7 iv�Q܎D�J\�l����d��{G}q�J������	Ύ��u��s�>��ڵ<�(��j�`_ξ�뚲��]Nv��̓׸�v��}�/�x�(E)o���>;���oÁ>Q/��(��,J`Q�ٳ�����XߨX���qI��z�u�oO3Ȧ�XY�Ğ�"�.��UE��3�;��]^�@����t��&G� =��}݇^�gwj�ծ��z��>����X���_����\�?sw�����>��u(SD�#-%q���QS?_�|:ט40�n�6vl�L��ceI�E==� �|�T�-{���Z��j{}�	�q&�zêy�y��J\�s���{���w0st��U$id�>�0N8��7�2Me���'��C��.}�;�.�\�غU
��]څ='M�d�������c��������I�T�*��DȲt͠��P"��g�����X#X�*�㬹�g�����}wq�+�hk����R��T�@bkk��!J�[���������x}k���m��s?wM%@Y)�5�ߔ�MemLR_�<z�L��3�}4d����":�~R���pòi�m$���]'(�j��G�'ԇ���e�M<��æ�٭9׀T��:�胴O�6"��@4`��]H��
qs4TJz�bB�D�V�n��q��v��婧����&�j�Nf� iys�|CC<� ���m��|Yz�=+���B��m�:�R��2}�tS3�q����xE>�r��j�fͼz|y.���g߫R��6����?�k�븹�D0۷LW��0���P��U��4��!�ȎN�����V��Y ����;�xF��:�M�7F������ӠI ������c����M�[me���r��֚D�Hf�LD�1���ׯ��=�VVR	�>
�b�C�(>��Z�t��.)���rk��Yn
>��R(V��j� �0�{8<�8�M,wc�&�ü�p2�h����GKm6�����g�^�ij�v91�G��%�	�����ޅsH��y-��i�g���������3;�fs��y]��0��:�g;�w���W>�4y���\�r���{�[��0�E���asGRqTP�r�^5�ʇ�':N�r#n �lc����`%0_�aseO��`�L�QCqs-k],����B	�ن��,��"W�ك>̎$i��y�F��X$���,m�6��&�Hcd��wonb�{.?>�}{g0�}U8���1H���!
��FN>H�>�_���G@��Zz�5hp������#h{B���JyD	���g0�oW��^Z\�U�VG%�����ÉS�Qc$��{�pg���Di������κe��8FP�&�:U�[]��*�*��T�:V����Ľ�c��? x����9�3O�l
�n�F7�������
^����(� ˖���QG���UT��0�Kn,6�Rl0�px��8s3����[�b��]k菌��U*��߱z����lr6�� jv��ݼ���7g�h��>�����t�o�-��*nP��p���*���''�PP��ɦ �z.�s\�2�^�4)�`�-������ZR߅>�;�s	z�6 �K���H��.�_&"D� ���z���E*�\Sl�V�3.3B�r�Ѐ'�dcN��S�e��:n-�SK��S��"+u��>6ɍyc����`��rb�7�	�t uTiHGf2��>�5;7��.r/����a��\1��t���C0u_�x�y���a �>,�>���K3`���m��e{�� ���S)���)�����)��w@ug�+!��Z�p��.d%S��U(Xv/�}�R#�D�C�ξeI��>������)L����<��О�e��Y��fC��\���;Kx�SF��'0��Q��G��O���7��ǰ�A#�D �ײ�Nb3賩>�2k�V����.�X�P��a�a��S�)<M'[{�.�vP���MfL��#�p�ok�^ú�oJ{��c<��e�\O��J]�C���jwQ�z�!�z{j}�j�oW�!L����V+�%���hf}�U�=H��)�C��۷��u\Ig�	��v^������;���Q웙�6���K���Zx��*j{iio��:�#��[ �	�{,@�M<|
����!�<���38t�~��k���s�̎a$�Fr4f�X�@3����7
�<��=��H!UX��#�a�%&�u7���]��G�&GL�]@F��=>��J�}�o�m�1�[4V�J)�I�7�����ׯ���U���C3n6i*��鰾����_�
�����,H�����W���x�O���W����YpZm`r�b+�<������$&�D_��Kf�F�Ƹ�}�e��o�:���?��ﰠgL�\#���py{�`��a?}Īn�5����*ֶ�����@l��0���N��}�������:�1>�;�,@�p�Hzmv�,�~�y��C���;(���^�֥ʣ	z��f�88����bzj�x���Q���n�~-��5޽qw�^�+�1෴�l�5)��t��l{���53�[H���bP���,"G��T�@Fݮ�67�{t�F��H�22�<E}�%�ٓGPȤp��(�6¹u����O�?6��V7V6pkg-�/�����Op��\{�0��i�<xǏ�Ǳ�q��޿r�KkX]�4�
�/v�埾jֿ�Ѹ�g�Fϝ�àC"OVoi��o�H|��j��&�חhfl�H�Vm2���Y���d�geц�}��7n��������<�(��DзŠj��OCt�Le]����A����q��&}/���V����}��~���ާB�_�4��g����p�_F��*܌V\4 ޡ	�&��A����6pyc�$�������D���,��0���Jƒ��U;iz<�VX���/j1���B�:��+�TϜ4��� ���n�|j&zo���[�^���}�C�#�f"*a�]*���r��p�"�)�{k<4j��П-Ys���{�����CW���2~a�A��k��ُ���$�;�ߣ�z��E�dR? :����UP���V�NZ�|Yw�oKL�������Kk���K�Κ��~g�zg�����r|�� @�!'��;���QgP��8z��>�h��ȲO"�� ���;�D�b�#8H��K��jUᗌ���z�&vMXI�~_��������&����/$��JrKijgJT����; 9ѤDs�}�D�L��V�1`�W�^4�d"AF�4>���Il��`sc��S���n.�nl�\�\��*7�+UQ"f,��{ ����h N벞�꽻I��9`�����w��~��z���˨Ez���u�	;��A��k�ɸID�#Ҳ�7��/����a0����J�	$�aϗk����ɳ)uf���QxsĪ����@���/�Q�/n�M���QXe����8��������Gt��L�m�:��Ԥe.�M�p�������\(po�$���"�u�C�x0��F����x��I߭�<����
b~�7y�Wk�S)#t��������~B��Ce���o�Nա֦�����������!�c#�l�%UF[���7������w�����{7ǡi��>��M��������$R6M�p�'at���O>�,�>�$����㤆3h�^�r	��!��X.��%��Q}��s�l�l� ���������������|w�"�b������_�&~��~���?G�@A���!�M�:O4����ĳ8��(j�y\��������?�������o`�@%�@P,�U����d;q�x��O���#��~�� Gp���4d����#�YI�����\���#�$���>���6-�;K�D��j�g}��
δ]6��õ�-���C�{X=y)گq>�&���ֶ%,āX*k�4q��"<oc�{��O�/*�:yִ�=]�����;����O�Z��7n����iԢq�PU�M�X@A$RF��7ࠁ�d*k��_'�+)��Svz�>��gf��v���(�\�\b�mܠ1��/���SOc��v��u\S�� :�,��w�����la��ҭ����?���*���;�&Sȷ�TN2������J��؞ID�۠��Di�f�	;���F
�Ju@�6���S�V�^~����4�����Op��71A��G�S2�M����:K�k����/%S�(P�agc��Cܛ���6 &5���oƸuw�@�2�������<Z���o\�}��>Ք4|y`��/�*�|�@�_7���+a��KZR�U�����:}�_*�:�
�#C��xQ՗[����A����kwq���f	���ġ})�P_Z-p��^=^�Z�~Π�� )K��{�t���H��CHr���`}���yQo�z{\��=�	p�ⶉ�o���������c��>@���15��Sg6g��;�����Oh���l9S�pJ��F��܅��oh��>FI4�V5-7L@Ӡ��fU�QS�q�9�g�7�v���.�����b��ŭnm�h�!ɰ�XX�S�}E7���2�>��J7�%l/w�J��e�l��;ik�*�m\�������x��ag�Fy��QlF���u�k)i��ʄt,�ne�,���ĚUJ��g�W�x�t�Z��}F����]n3�M�:ri�N�Zڝ����<W���K^3x�����_S?J�뾑¡�Gpv��#):�����>��0V��=LG��[� ���E���O"hz0����W��J����0O��_���0-�z�k%��D$�Q�\R�� �����a��6≠Cd��!���ԸM#��%�#p�_Hr5�0�t��}�����M^��B�Ԥa��V������ (X��P�W��w����(�l����[��s�� ��ڢ�1C*uF�����3��l��&h�Ni^`���H�o���n�YC��྘LM�k�q��y�u��0����������%�)�f�o]�$�nfԍ�c�Y��B�?�wr[�_Q��y2ҝX+!�]�����:��pe�V��vř����Б��_ǣu/N$�0m���rn����!/&���(հ��eP-^D�ήƽ��-**��&iڽճ���;۸īx�(V\����	M���X�ob��~�?W7��|����^���;��G��]�5����Hv��O�����u������s����MdP�=��Y�=�֖Vq���#�Ocj�N�B����⊁�(�~Y�C5V��a�6�f��D�볾�Ǐ��5���+�����E�Aʌ7������Z��k��,���;�Z_��U뱜��?���X�:�#�X�6-i@(QA���p�ēx�?6����q��q[�@,��utz������tS�|���M�C�=���ۇ[� 5x�Zt�yC��iW?v#��D[YW� �侽8�y
�`����[)t(5��#ñ�����N�H����o��7_����g��O�)cz�<���X���?��?5�G����)'Q;W*��iǢ�;��o�>�Y���F�ӟ~;8����D����b��4�2k�*��a�L
7�_�_�1���N��hg1�	�^��d�AeF򟾈)eԺ"ӠI4�D����Y���x��m����b{���c{���|;�N��-߹kӣ�{&�`���8��ie�vo]���˨`o�#x��g�E[�R�#� H�ک��x�＄���0���:�� .�����K��p�Oa�s��~�S���ۏ �aix�r[�G�n��o���c��XUE��0�g��_S<�ֆ�C��U�H\�#\�s/� ݋�1S.[u'2>��׵���,�J�|]��'�s��R1-�
E�$�x��C8r��	��|��W�& s��{˨�Uvl&NR��z۲�jQ�x��Tu���� Dg@�!3K3���[�����4�)E`ѹ�	��/�˕T�uY�X��W��0�<���h'��~�$f'r8{,C��%����b��d0�e�_���26���\\�_�*��=��sy4�z6�P���Ӷω�����_�;���2?=�`O��Uс��Ȏ���M�����,���N/����N�2���+�r�&�dQ!��Gk6��f[9�Z�a�4E�>7u��L������F�)�� �W!��	�Ș��+Q�TgO��\�&�o!�����y�*�$�3��=�F��͹��={���u�� �ޡ��U$cM������h�0#)��p�:�n`��I�?0�?{��_���щ�e��kK�~g�Q�A�Z��������Av�5P�p@�ǿ�!�Px��`�܃Ҝ��w.�j}���|�����l�����A��5���!�>t��6n,auuӼ�ւ�ի�q��O#��M�mv��AM�?���:��f����_NJ�mї��"tif�\�o9�M5�{�F�%PI'B��nBe�^?�b����>L��u8��j�u;�Ӷ�<Et�gNfBH�'�M��<�%e��v�b�a�o��Zh3����j#ȿ�(5��Z4��v��Y;ym�;�]�3ݽ/迿���]��k�Y�+�uY[N��sx��;�=�8��!��Ǧt�8�-��s����CvzC�p�����H��^ǀ�����(��aF�� ��=b[�S��]{U��^�� ���U��=�w��Ba��Z^�\�{xe64��D���\\E��~���R�q4j !�A�P��&��������&�mrO�g�&q8��jP��z�)e����L�Zl��Pn���)i�[���z��<킪6�48���D���o�6^���1:1fӪ���h�+6u����v	:�䣟2�%�F	������a߁�H�2vq\�q�J\8����آ �Fg�Eh��wL٥��8U������a�f��w��?b��)�6&	2SC�C$�oq�>1w��m�@��/�_�2>��s�!|�+_�s�}�R7^z�#8�Lж&��E%̾�t	\�SB�j�N<�1���,
�×�Zp^o�g0�u,��8�� R{q7n�F���/|�Μ�ӟ���Ϳf��@������~%ՠ��E ��ayk�{1j�M�W_�җ���|��E��^z�j76��J�h��z��Z�n��
�bɄe����;p��,-���Ƹ75K�+>D��o�z;���:���� >����,�"#'�� E,���F�i}nIe�4E�/M@`t|�8X�V7�w��?@�F�H�M��%g]�z�>f�/M
��)�d��.�έy�K�q�׻��p�#)D��7q��;�6,ȉ�}}�S�n�po{�F�鐱T	�<kǇ�X�.�½왝Łg���~�c�]�i٣=�c���`srK��^l��~Օ��j��ʭ���Z&N�;wew�_E8��d� &�A�߭pk{��~�po8k���2�;^N>�_��sHgx}K[��������E����UR������pLK;@���;�E0e�]�����vF�ξ�j���TY�4�b�U�^P/^�8�nZ��[U��z��r���Q���1E,�.��|��qxo� .��`��R.�B���t g�����#p�:.ߦ/�u����Y�Zq��,��Y�vvP��a�g
Z�:��]� ?�3y}ڰ@�A�*Di�Wv\]�[���c,��GB*�Ց	�10��x�����Bt��#���hhs!4��G����������s��MZLi�Ww��(Nݏ}��3�����Dt���e��K��R��N�ڕ|�m��x����x����ai�e�9����g��wP̫_��� �Y�??D'@㏯�­��Hq�m����(�ˌ���$�d��.�1�?�5Y<w�:3"q�9�b�zʭ�-���U�������?���p���vKs�r��{6Mk^v\V:Հ�I���&�&�I�?F��n��#�M�`��	ܻy�7.!Q-bu��?����N�ϥ�����Z]�5��|�+S���CVC�R��_��e-��ڐެJ�Ҽ�A�D��u���0څnǍT2`�z���^���¦97?���ɘ	�KI� �'�H�C�s��`0� .	�l�deb4ҡB#�:K~/��=tp���J��Qoi�\��E�/�U����v�4>0���Ʊ}����C�h:�y^�����֖`=�}��S/j�� �7�0�>��'`oDخ����@WW�Gb��P<Ĉ3�=��'y>3aQI�G��G���JG�&�)�42����q���� T[���qT5�!~�f��H�C`�a���:�|�5+�����k	�z1���<%W�Q�NG�S� A��{��^��u�[�� �x�8�J#�i��3�5=SO����2R�J-�Ie��R;�c�>Ň0�g��b��m�>MË����DӃ��K��g^�m@���a�i�w�?�ľ=F���)"ͅ�ע�(W{���*��>�y�Өr��w�TӜ�����sݷ���ݕ;�+Ej9�!M���F�¤DJ��%�t��8_C�V��}6�P$��}��>�͍��5}��eO==�&�gl #ǵ���ύ{t4�Ef-���"\�-�VJ����Q	֤�,92����z�f���Ӥ`�������(r�7�R�c��׈�Q|�|~=ɢ�1��@��K?}�Y�� �t4�i��j]��˔n���q���U�_��k(`dd�h̆6LiC�H�ܽy�a��+��o淭��@@�j��y���c�,���|����b��E�N�-�9��MڐU��k^��C�����ؘ���d�	ܛ��R��&i�L�]�ф��꛶F�ꜞGZRp���.p��6K���<�|+��s�/!�g��I��y���E�^]\]C��5�V�����w	0Π������ލ��:���w���O"½����ZQn��ޅUt�_�����6|���9>�m��{S��Ssǐ��	�v��t�d�6�����[`� Fc�\��"���r�|��ݸ�����"����-��#YQ�	X�|�����˘�;���?�W޹�k�F�&9�v-�3۴A~�!j��k/(���������f,�3��K�cH��ŒF5�l����-GfO��%��\(o�w��ɥD��sc"��&�;�(��O�W^���m5�C7�S�&磱e��{<G�~�(��Et��>��O�{������Ղ�����9�đ��r{��џo 6�v�M!���A��o����h��ұ����k�/a9�Ëi�pt�#�Hٟ��T��G$�-�^�lRJ�R�~-t�u[�鈂nL��a���������S��������kp��oh=��A��e#�QF��8h�I*��"Å�7>�O=~�6���Vp�r����ƻ����#�ay9����6�3Ofi|zx��a\��+6lD_Z�u�Cʼ��Wn`����Sx�_��k���w�([�j�F#�A��*��멑�c���Z6A����s���K}^�l�݂go����r}D�v7[k �+�J�Jҧ�ހ��？q��PN8������7��4�+��Z�"�2eq��Gv�|m`�󌞛�L=B�l \ŗ�&H�+�{�dְ���-TJ�k?�X���柀�~����\2�p��&�vs�brfR��g0�)&��N��~+�p#D��-k�Z ���N���g�|ߑ�4�䞇�?6����i�����~"�n*�Gg_�5�	���n���3y>Q944��	G�{��3c��J����H|��5�P�QQ�2��Ǟ�e��A���P]�
5`��Ժ�	^�Ǳڷ��z�ڢA:?���	:�bq�Q�(Җ:�Z"^9�_S�zŖ�\����J����%�H�@jW�/�Y�#�ۀS&�h��͖j�s/=z�{Ʊqo�F:���!:d^��V��������D`���#ʌv��}`���{W��)��ϦYŘ�o��Y>ȩ�e �\�V����Z����?C"R�I��pm9�w_�ceԵ�%���; ��,lo�����	(��;֫�'�,_*�Ig�C�>�����
�i��ly(��������t4q˂��mm^�)�.���3c�.��?0��l���EQG�um���@�)�Li���GGk\���	��/O���&�U�{eSS�"1�9�������F�O�7Ȫj[6=fo�.�Z繞C�PQ�PRl�T�D��Az�k��qe{�Le��6/Hrh}:�Y���� ��,�ch8��~���E,D�	�t��-S`0*�3e�xտ��u�۪f��h�XemUwT�W�]{2������X��%Н��z.9���>w�#c��󸾽��i�6=�o�P�^�_K�7����ln�j�����9WկGy�M��v�����y{�[�\*���޷]_�6��'���U��3���q�(X�j� ��f3�T��ɛb���,�R;�O�=��J�\Y�(o{�����8�lǳ$#1�7
H���z�����kK������j�4Z����";����u/3��j�8��k���c{S�C�}�V3A�ǳ�����J%�\b��M��u�k5]�����a<t�����ҫx��y�S7���Ye�c��b��W�{��w��Ҁ�� R\�	~v:����]ڳ�ʾ3���L��"L�ڨ�,�2hp���u)]0i��,��,�+�>oRpH��]Q���'��g�N��ў,�X.m#��75&
�b�>Ѥa�A�*����u8p��X�;�B`�j�y�g�z^�V�Sm��������W��7��#j��rE�6eÌ��t��]��W�o�a��@����0r<�"�m��L�L����r�c֗���P�6���E�]Қ�Ј����������هƔ�U�9m���bv��@C�eй��n?�25�|(�x��9�d���>p�xΏ+��bu�=ܸTB�I.Xp�w�x����aN�3Ϟ��H'�����2征MwT�#�t�X�ll����w~_�ҧ�O�����u��8CÃ�i`�Z�� ��z�Өe�T:���eE�6���2|>Ye#�Tq�F���:�^�r�)��a|���=g:�=�7V8іx}���!���jWK�22�0ji�@����WٌQ�r}	�f��IxZ��y��w/�SD�jG��D�t�z��pUD|�{�E()s�kt�*"^l��SZ�<��V�΄��%�K�%~£� 2#��\�����Bf:O�W����\�?����OO����	?̀q�)"c@�h�`/�F8��Z����E�g$\->���D�A��m���z^o�XE�F���.�^�N�ٲ�۶�z�$7&�b٢������ ��g}=�F�ZtT�uZ��2�}���t�&8�|n'�'n,_Ȁ�A@>���;�������1�b��K��"�� �q��:�=�y�͠�������fѤڊ�ޝ�t'���n�ʽ���6l �cA~,|�M�z�����y_�F&�*�У-8�໿�'�I@~�.��o[������4�]O�������[�$�-�������|-;O=��S�3�h�{>��#p�]\�(�G�{���]���&�	ԫt��Wq�u�a��	$G�P�m�U*B�Z�ꛘ�x^Q�T�ȥ��
z	�o�gH,���{h�i�<4�O�`� I��P!�}��8[ł�D�L+ԍ8A��Ui����$�.�0AJ��[��0p��@��w��.��,���r��t�܏�J�Wna��L��&�x	��Vo���e��aG�Z�&��6z��зeE6ᦣ�#��?Gd��N��e"�0@%2��c�)�����޼h��A0�2��@���.��R�h�M�"Rۦ�%5��s*u����������~g 1(�%({2����vZS\^�^gԂ���]��c��x~��F%Ѷ�����{vz�5n������q0"I���Z(���,��l�|���3�7�'��`��f�3���opk�8���v)��v��H��"LV��\1�	R��k��VE
����4�i�4��mz���bjaC+��=l��Exd9C�3h(ߺ�2N��Hn�A�v�4��ѯçO��O�B�{o �S��s����X)�>���Ɵ(բ*�-䋘-P6���z���av�}�{�:��=��m>�lz.>K�6��S'gq��1�`���_}�E�X�k���`���ڼVM"q�>�Df{��}��=�t4���Cx�#8��n(PPR*� ����	��L��CU��g�-ҧ4���)�d�;ח�I?5�}r���o�vr�le$�u��--�Ҧ����<�'	��7�̳�v���q�q�{p� �X����m^��O�!�2�6A}�D�k�W�hc��% o������D^(ի�/�b�����y�E��c0C�ĪҬet�0�.��d��e`b (.�Tu!���U�M�[t4n�;�gO�SgN㓧��>��Z���R,g�>��n���?�>�Ԫln�ؠF�@է���)�c����47���=�N��x��?��s�8vp
sI�������}Q4��;=��������b�o�'������m O���H��*s(��	Ak��t�[�ѭu;�����iX�N�kM�JQ������q�9v��}�K&o���N��P5�j��n3�.NE�*Ie�	T[~�h��C�*���K��N�O��d��h"��Д�3��V5V�s�:���5�ֈ�/��"���6��4�'�7C.�����L�a�'��h��(���0�^�`�������=��7���!�}]�p~S$!�5x�u8��0w� ��ݧ3��"�S�TF�IJ�+.>��/�5�O˙[�G,�-g��P�@��;��4��q;L�ݾe�9��柆eBl�YM�]gpF%�eODgS�^:��Y����2�T�C��}�c��*�ϗ��D|�a!I� xp�4$&wMǆ�F�mױQ(� ��U�W��v��B�j쌾?�gjE��~�O*�5TZ�~�@*��)�3�,�/]���]x�	|�k_Cs~	[�k�huh�<��z�8���#�N#��^x��އײ
zZ=eý�1wߢ��۪Z�c����3��60Z��\U�#��hk���	&�؆�'i�nU4xo>e��!VF�.q������-�Y�w-��K*m	$T�V��2f�ba|��q%�ٗ�;FWc���RnJ{jx�z�4���d�ܦ++!y++Ѷ�Ru��Ժ��J���`�J(`g�J6�:׸�\�8�4T�������f�	!~D���b�$p)��i?hI,s��O�ut�2d���[�8"�Ze�[ʐ�F���kjoQ ��q�a\޳�t<�geY�mH�UA�b�gY&��ډ�Mv�vKӞn��
=�����v����|phM<])y�}�B8�g7�g�ʗѦM�����lx.�kPv�g8��{��p���T��� �i�@�Y��}28������Ѩb���865%*�0 �V��IPe�{Vղ�^��0_�&p���Oygy�--#HP��3�K?~�;�8H[�,nhy����}�aL?�4"�,n�YFH�E�Q��~#g���G�'���@|~�{�k��gT@}ӎU{��ۼR����3�P��wЊ���=�=u�QCN��|��U�E� �o�����>MP�M�.��&�Qk��V�eʖ�
J�-��C�"��(A���66��~���죏��0�����O��u����Z�>N+�~���[�2@�����X���ƽ�E�,]C���F7�T���5S�9v�@��SH$�	B���M+�hpO���Bi"��݃��,�����Z\ù���y�1l�nc��=��8���dއ�����A����}�0"Z�W���k���h���TJ&�,�X�F�X�r5=��9٣�&H�xG^��)����Q<��|�38y� &��U��FX%1P
4�v/���I|�gnk�9�2H"��w�,S�C#C�$���bD�>"�>��ҁ
��o<84-"��}�:!g�Wo�c4m6�Y����_��?��?�i�Ϳ�u���WX��!�I��U3��(��G�7�������{��Ȕ��ŉ�|}g@CW�,��1�p�����_.�Yy��W_��u���.�k�u��/LC-�����ۑØ>z�j�k4�t���"a��J���ͅ�u\�m2�K %P�z*���qUOU�F�u���L�E���	YV�M�-���bcQ#9n0�5��Hc�5��Z!}��Qʿ� O#��b���{w���!/_�c����Q4�;n�~�nn ��C��<����^˦��m�?�@�|�`��wXX�=8�*�F�̀�m ��jHк� � E�~:�pCΪoƹ#P��A_�X�����&~���ZE:��ښ5i%��DL9E��L��z�

�8��]~��ٸZi�J6�+� ��sATFͮo۹�5�������Z/Q 췬A�N�$J�
�Q[�K<Nn�"�3�Tb�䬫����/c���Ծ�H�p�`�1O�Y�"��!�!�+c����&4��1:v,�(���V���p��^SA�u��7��m�y��s��sZz�k�O��xQ̕��!�^�#�	]� M��ö��A���W���|����[O ����m#�fp�QD�QB��M���~g�O�C�鳖�=�LJ"5[{�����qzn͆��Wk xܖ%n��s�/���P�+V�d�0�5�@	T��&�cV��-�k�QM�zmU�(�������y�)��E���R�L6�A!���nٞ��`�z��tꚨ��&�U�j%��Ccr�වa:�lԃ�r�x�}�~�Zۏzݔ�UU˗�_�	Y�G�jG���z�	;�m�Wf�� )�BC���#�!��ex�R(㪿���h��x;���B_�y|v|��@�L�����d�T,����n��[������������f{�}�y=���ۆ��֤��p�>�y�����{�e��*�8���C���b^l����1ܩ�@���V�����*A_����m4���>q?�U����?�ؿ�������7�L�+�d�0��ψ|�&�Տ�u��7�3QS����d��ɑ1�}��U��s��3�|���x�
����A�P$̳�F:Bp4�mb��|�>��X�Ҵ]k�k�M�7^x�{�I߷���~W�!������#��_��P�(��@����>T&G0lb}g	��t�����5�q���\��m,�%lH��8��\�~���Y��z���^��/�M���r��b��O*x��E�����?��7{�(r+�K:G����_ܓ7�f��������7n���e�&g��y�Z(ի6���;4������!����+a�AOB�ճ��O?�o~�380;	G�Ǝ�����w�#�kM��1�0 뭶��t�~O���=q���i*3�HX�v�r��Y��n�ޚ_���-��c��k�̗�� >7�\��&ff�����o��'�=�,=�+�s�����===9`�3@� 	� ��$S�d*�J�U��֖]�r�ʡlo��gU�]���R��+n��#� ��8���s��9|��y�{�{`���(�LOw��}����s�t���+���U�E�P�k�>7��������J9Oe@��<�v������M9f���$8�ڰ;�;�h?����2J*�  S��gI^w�^�`����C�Fn�|����%��''[����
AF�s�0�ቂ�{'L "ްJ���(��h�k�J�����ǖy}-�G>�b>��R�@}c��}��&�t���&qh.�k���B��4ͦ�@b�o�܊�{��b�N�a����1�U�AY�ʚ���4AF����9)����/�'`.�������x���h��r�z��~��}x5�$��u��r�^���j�!����h�fB�A�E�[G&n��VC�D����"�,��m~�Y���/I�X�>�0R޸���,+�3ڵ��SV@@R����~��P9�g�XC���~�Cl;�OmP)hxh� �O�7s}��!���}�B<�}~�d򈖶Qn�͆S��Μ���%#w�mW��	(T�#�o��U,a��e3'0���y~�@V�!FJ��p8HSĢ>�WJ-��I�,1���nس�&�8�<W��KY���)��C5</#,G��+�k+1����o=mz�*��d�O)�j8,�� -���j�𙦸F�1Bp;�n$��@��4v��48���Dl�L�e-70eݬa���|7�c��ڪ�^�V�n�2�b�� ��cX���^F��{07�[y���ބy_&�N1E��({O��3�X��
��f@��O~0;���so��ZV9lk����SE�^��:�Gr��'�@��,~��gL	�w<�\�B	��Uk��Y(�,�&���2�F�!�X��,���w/�B6�`��j��=Q���[��?�u�[��;F���9�r�^���$W���7M�k.�AF���<�Pu@SӦ��w�<��t��$�7�l RF�MH�A#�M�e9�*H��������脋����K{B�O+a�_��2������'p�[P9]G�gx� y��5loo���9���@m}�x��io�܉��[�q�%��<��&Yx�A������*�0N@�c0R/�,�(��j5�R`Ҩ�ʕ��*2&�=����6�*%�N��MWX��ĩcx���ͳg���m��%y���>A��-C�'5�3gU2�GS�K=�^_u
[�݃�����}waVU	��xkի���P�L�?�F��g}���i�'GB?96�1�n7�P���Z��~��]|kkg0��?c29e�Z�7y�Oi�_@i#��q<�F$V�vq����6�巯�/^\�K＀��
��������u�&/f�׃�L��E���r3�x�ίmZOU!�gP���,`SN�!����z�ɧ�D�<8?�/|���cc�x��m����x"iJ��V:�jAtW�s��^"Ԕ!�҆Sd���X�#<������<� R=ԺM<����]B��3	���4Z������9f�
N�YNf|n���b>�����o	o�sm�Ӥ8����!-g������1�i��A�U�}S��B��\o��k�ؐ�f�f������)^v8F�j�Yٷ�0:�F�����/� �}���YFK�4�ӷ@]N��Z[Dwfۓ�&�?~�%�~il	�H�&RD+�xN�P��x�5����*���{Q|e��ayu����*�#ƊX�W*�`d����*��ԸV��4&Edٲ��Є �k��o���CS`a2��\��24@��ϴڵ򞚸�ɊMՅ����Y��c`��px+i*2�������QAݼ�\��TF)��N������2���D��A/a�mM+����$;�q+Q���um�G�Zj�F�N*��(vf4�I��(�(�90��\����mCi��pJ���m�U��V$(g������M��N�Q�6��&�w?u��t��\��A�EP ����T�.s���жK�1 ���ȷ�x�Hw�yZ�׌{�Z���X��?����%���h�2^�X_�І�$:��H�����6��G�6ŵ�� }'l{AZ�>�"��y�=�O�ݙ%P���E��4�%*�e4�讬ʨ��Q9k�9aQ��sK��kCZ�$��a�@@�Z��a��	��͖��tU2¦V�ID���#����[�>lp�g��q'����;�WFK��^���������v��U5ޗ��f��h�'���s�ƳZ�矩n`��ՑH��TB��^�Vƿq�_t!봗/W�q���T�X�&�.ƣ�BH\���R%G�

b4� �}{�`G���/|���+��� H��~��p�����q��W�{'��Y�e)� ���ئAYI��Fb6��[m ��1p���^ѻT6mRYRh�d�����u��Oͣ�H��~��
^��y��h�ʺ"�M�дz|.
آΥ���v=���vkf��(PP_خ��Y��Mjđ��Į-wL����W��M�b�gѫӷ(9rp��y��ޗ�a�t勫h<Ý��[���sm�[��&|>�v�kװt���<��+R�'X��L���p�o��Ϛ�n��ج�)vxf�X)^Gav���=�F�a T��/_ƵkW�ovS�.//��Dҝ���V��s�=8{�,�>}�v���k��ӳ�F��\�v���%c�P�H�Z�~��g?�)��g�Ľ���j��E!�|��/beW����Nps�V/뫖⓰M4�. ����p�\�*�+<q�I,��0���~+ۛ��r��<rc����O�|_���x�}3��?��o��<���W�nڪw��qp.���Փ8|+�ګ�a}ss'���]���������p�[��ԣhz��V�]��F�>Y2�50 =�z�n���7:�n2��+�̚t)�{o���ؓ�97��"��v~2�������ڻ�7?'�t|w��Ӳ�5z�7?\ߜ�:�r����y�ߟ�ոiz�s'�@���Y��9�5*���f��?�ӯ�O|O|�#Ɲ��_�n��c�"RM�i:Yr�#����3��7,ǎ@�L���MF��$���_nvW`0�r5�+�/��p����W��Os��rhrc�E��(i|~��݁�h��1-��X[�T:)��"Jg�Do�QJ�g��)F��S���ׇ�}z�b�x!��	�j+XZ���̔5��4|B�8Os����"�<�E��m���7�8uM��R��V+Y�(&���}>�C!�t���� yF��D�t�$���Y�*�q]�w���;����3;����E6��	�ě+������DT&h�;I�A�Jh��m  ��IDAT�q����-���ȃ�����D)��lB:�{	��Q��ZE�R5Q���8����\����2��nm��n�W�G@�Y\ĕ��|�6��r��iK�U�~�>���&�.���Ie��'���6�\�gɗ�R�L��]~N�����$ԭZ_�B�����Jњ�Ó����ʪ����H]��ҡ�kx2=�D� @�m��ITu�_���m ���C�A|BS�NQ�΅�0p"Ю���PFִ���s*���(G����8�X�آ��u����V��Eic�#"����H�<+Ю
������!�v����1TY��Up3�T� [	;*�Mr��PA��ŴW(�6�8��H�V�4��R�b	)x���#�&�)�2ziMī�e��Z�o@t0��T�+��6��r=�]�����4��L�#J�>�K��򭃨�v�"hw��ŉ�\K���<K��_��ci�q��B�R���6�%�A0'c��:lԻ��Z�,�#���bq�]��7;5�b�?��Z���+L`V�bݾ�*�#ܠ�˶9��Y)`�#㨤���]?���=�а/^Ԟ�|z�5v�c0$���}����O���������>�g�!��el�~3قIQ�y� K����򒈜����:mBͲ�X[���|KA݇��?bJ7O���9�>���"�L��g1V�ơ�����4X���X[[3����I��peK�������8����C�5]���(����{�34|)?�:�^[Z"��/���I�o~��>����F�����S����n�gw�߫'��z[�,�o��{84�Ň��g�qumϾ�.^������U|��	|���#�[�qu�2�����8��C��#��
\�r��s��Gǭ��i����|.��YSx/m�=ӵp=`:0�Xd�6���ٷq�����A����i5�lӹ}W�u���{�����w����O��y̦Z���5A���%��E�v�kg��&��Ξϸ�5%�N���9�ԏ^7�>?<���*�i˛E� ������������?«���n!=�D�H]����%g�I�g�EL������<���u���l�wU��R�b<$F�(��7�2x���!��tk�Q����T/r���w���d�F���X�mFk�wi�u0�K0DX�1)2FA�m�_zn�$W��nC߳�М=�J��ɕ5�7��1b�k4�KѮ�C�h��%��(�+E=��W�R��4%�e�.l81��Ř�^�7��[-\��I0V��BΌ��d������X꠹ݷQz���C�ب����HkQ΋�r����}��-d�xc���L�����-FWi�����d�k��C�V�<��/#l�!IW��$^4�l�9pL:*�\�?�,�k7�1ʋ���)�Iܨ�@�E=a�zJ������h�c�(��ְoC6t��5������������,|��A�v�g�T
j�P��PixX��`����WW�o-��\��(6u�6q�X"A��~�NQ����@���ʡ	�EپS����=�԰�|������7P��w[%�h�4lۢg���xJ�(qў�q�NaÀdX%�6߳o�'�8�\sx�A���������ȩ�w���uu+�Ƌ��$�]G�FA�ڣ���2Q	�j�I �%`+#0��Ǟ�/m��=�ek.we}mH�&�\::�V�b�=ӳ2vdX]�k�F4K��u��#��7��
���4>09�7���4q0W�t2���Dv����n�6J
h�6܍��l�Z�'�I������e���%�u�i�Um	,/Wh}|�c���ͪi���Ľ-���<�n�ʖZɓ�n�W��������w������~�E�#61�h��uY�+�>�Ͻ~��#� �Ddb�M�����x���tV�so�ƛm������>ܓ�@A}����}U9
S�^h`�;�68p�rC�I-D)�l|td��aO��H�5�<����@_�<�$߳U,�K��*N[.Hjy�r��&���:���@��n���Z�Bl!���.ob����Lաׯ#x�[��A+���[(���5�ѹzA���������8
���L����Y��q�����NQ��da�����s�Ў�͎Y}��eA�h��Fg�����������Z�L�.���2����x��K��L��W�Y
ۂ�y�υ�^m0i���Ɵ��G����'#�J�����;OC����'����k8�E���<>�n�s?�y���{��Z���߇�Z���[�?}'G+��g��� &����b,�F��g��4�k�ﱤ���ޣ�-~S�!��+x��\^�b���Q`�RU%�IX�X�ڰ�곌��kش���:<~�A���3���6m��M���=���,�s���",12�4���4r�ԍ��˛J���Gu=rȼ���$>��4����������׭T$�#�6cQM�e��p�USԘ��auk�����?�}����7��R�i�1�|OX����T�:2^��C�k�^��K�z��9�4��,��]Cp�z#��a�8|èZNؒhu��r�5�Kb�F�@��j�2j���Y^Bqf�����ȉ[�왷Qy{^����iT����f���G�N����0��بQj�L�O]��,�P�WK{�+&:���$.�{�Kۘ;8u9��6�����)4T:U:5�^���U�ݡ"�ʂQ�����c>�*��&�?�����:
|�����&�1)��Ʉ���qk�	��8�TrRߡzH�I�>MO��a��f����D=:��o;�>L�-#�a��5>��s��0�&�ML�F���T�JL���b�v�҅ȟ�gD`�z��Ԍ?p��ڻ�F�Ưge���H=;��|��jy����.^��^i���TgT�)d�v�m���M�P�ËZO�ӂ�qs@*˩OO��>N�-1�GB��Տ�$Po֫bBw��I�y|Xj�o4��71e�M�V�����ʩ4��U]��j\�V���x�k�x�h5@��Y-.��p�Q)���v.�3�Ȏc�״�jб,���{h����){���YoeH�9ު���Y�0��E{le�̵J�{�|��%��I���])�"@'B� fcʆ��*��J�|��p�*�Ƣ	���zSO�:�àΩ�g!`��q����ې���H�AYseҸgN0(�Oz<5��H�8����̣z9���m�1��Lusc�4��l�J���"�=���������3�#�wX{�{��o��W�o���r����`��qum�TĘP�7x��VfU`��U#(�z	4��[��y�X�=m�h���>r3���F�G 3� �\���@p�ML
<�>7�x�����V����dfq���F���S�T$s<������^�E;/S�ZFv��čV64,՚f���A*շL9�z,�2�>�t�^{�~&C>΀�-_MP�q�<��z��IHuj���cϕ5��А|V�N�"�r�M����}\cQ�5?�3��7߾�2���Pn���F	��f�������͍0K�}�VÅ�U4�>�'�P��Tn�,��r�Xs�(3p�Q�Y�Z��a�BEy~�Ƴ�klc�0�O�C����"&��*Hd�X�L��?i�*ңQq}����{ɟ�S�=+/�3���V��mz��;�q�p���	�S�����o�p�˟w��0���:����񭿾����#\����[�6���^��w�q��>�*U��K�vp�K��}!�hu�J���ܨ��s�7�8M( ��3��z!i�i�TCE&^M�$4��7�G@��C��'��}�y;�"
[�����H<Le�t�?.���:OT�X�޳Zm�O���&n9y+��L��,�^hg�v�36�@`�������M��g��p��k%�Kn�IK��;pao����V�Bg5�:���.^����=��ި�������F�|�Rc�Bk���6�Q*VYK|j֊��O*#���J9C��7��4YwЅ�P��N+�P>My�"���h%�����b�����W;M4y]FΫ��\E�ہ��,�0���,�#rpSdy�
�t��A��q���xd��װx���h�^M�KO?�~�d%o_�ܚ��{}����Ȭ/�	��Kq��Q��fQ����0s8�{ 	Th/
�(��X0�;���RG� ���hԤ6���o%Z�U���r��c��$p��u,EG�3���0.�Y�J�R�P/����F��z_�@j5���E�3�W7��=��^�i[)Od�>6�#�Þ=E�V���ф�w�S37��B���&��	��H/@'z�v�oD�5A�0K�*�׶J�*ج�I��i�\D�{2�M���&����>�w@��>r-��X,c|W���S�#�%bHT���*�l���
j�8ޓ$Ж�$Ewd[g��/N�mC�~
���,	��)<�z�h��������Eݿ���`A�Q��-mx:���w�3ʅ��I�;�����ߪ����Xg������t����=���@����*?��(�66��y�N��^�q,��������` ЌgP�~�qHj+#��=ڄ�������O�^�D��U�V�1�R��f��d��߳ll:���h�ۣ�8n��kBAG�����M�F�Jgm� ʽ+��4���ԑ̤مd>a�^�PUE<��&�����\�p�}i�{��m�����O�>̀�n27�<��OZTI	��6��/�^���3+���o��c�1��߯���o�_m\����`�M/����p�<�ַ�%2�^8�P<�gK{P�9j.a?�����h���B�ɣ��n^�қ��ǌ�r�<Js�Ȅ�8�O��=w��P�ݛ��]f�J0�W*ֻ,ʰ���l#��WU�="۰��M+PS�D�@�M:~(��|`@%0���U ���V )ڥ(�΃�3s���I��������j(x�҈����Ӥ��j/��|x#��NHо%�vi���(�Bs�(�c��<�����	��Tp~���T�Z���+b�$i/��g�r���"���1�9��D4b��L�u��YmQ]�qϨB�j3���IJ�N���o��R境_��c����e�$�j���f�2/�[S��b`���� !e�?	W�3a��C��ے�^/�Z5��:�}�&ެ�#_�I����1O�P�+���������Ͽ����o^�w_��j5@��.μZ�=m�;�x�e��"x��6���8u(6��X���!�p���68����+�
��x��%T�����V���c��:�]�N��M7���k�X5���?�(��������HmdEd����ܜY���5���z���׌(t~�����'����+�82;���+_���/��4���&�]���&dE��*"��H��i��x'`fn���}�u�<+ΠN�1NcS�$�S�^��k��M�,�������C��̮o��7\Wϥ���}0�N�yC�rrCV��{#�-"��v��C׷�6����-��m��.B�?�)�iX C]�U4P��I�|��ؿ]a�͈LĲ�lꛛѠ�%�L���D�/Z|�-:���H%	J��Z� ����tĲ'O�`�D�\������uu�ʈL\:le-��"��������a˪�2�ZFE�%�Yjp}4i>�"�=�Q�^$@����+�E�d �ό�/�ձl)��p*�o��6z���lU?�ٸM�̞�S�X9Ic�wk�I�a��`�<�yNX�0��
�:GP�,;�& k��_ AӳzFp�~.nձI�"�K~tEZ���&(���{�U�x��,�d����!�?51.�ѲV��A����aW�����*U��ipɳ	��M.��fLE�0��岁ʔ�C��wA!o<leO	��-�Uw���4;�.M�X,l�k>���U���',��ϐ�T����ג�6����S�R�H��F;���^H�	M�^���t���*[F%�K�"��ym�Ԣ�$��C��J�wR}Ǎ�Ya�fza�qnL��w��H27j����!���p��P*#�8�qS��6����M�2ٚ>U#%��>��SD�*��Ʃ�j%0F���̦K*I�|L�Fr|�ROZ� =[0e�3������iRR�#5z�u:��p?������ٱ<�������K3�K<C�Qot�odxYl�9\��F���
�_������¼)ct��}��ڷ��"6�)|೟�G���s�J}��3/���,^>���1���U��/]s�
G�g�>t/"5o��Q~����ph�#ܗsك����&�KIz��__���5�,ԗ�1�f{~jP/����|o�(�-�!J�����l�~܂��Up&A�%�vT-�m%֖c�A=ы&��	w�'h�C$�7����e� orΤ	c�}k(Pϧ���B�����M�����U�WP�fƍ�T�C��qq�Ʀ��\浔]����U��54J�86�5���߃�MS�|�� ^�q�*���v�o&�����a5�){�I�1�/|�s��/~��M`����Gj'4�'q��ď�0�k���ӿ~<� �L2�A\|�)Z� >�q�ߖ����w��7��:~�j墏K��滧�pb�z������j��_��R<�#���?t+
�Ӵ��p��3;���d��,-���g-["2d�6�UFE3"!����SD]�� no-��n���?�n;j4bzi��C�ݞ�л���T3w��22�C�dR������ĝw���D��z��s�zָࡻN��>���:���i'���*]P�OC�-1��X��o�5=v� �㌒r��Z5�^�ue�а�֕Ok"�eT�sO+���^V\v"���g�ʷ�%XoXX��h��������!jk�ʿ��P�x܄�-P�P�ɤ	9��CU MT0<4�H��E� �g%������6^~�-Ďފ�@��!��ji[�␚bԻ�[�W��}�Z�ch��-x��x�w0>s#μi�f&�;nۇ���om�_X���-���QQ�N)}���z3BB2ѝ�{���tj�T�8��B�
�^��TY�3{J�6�z&$l�� 1�������5)~��#W�HD�H�a�����X�����1$e
F2qj���ke�;��4��sۮ+�5U�4�5������-:R:��� ^ඈ&�cRp�&	H�h;�����´�:Q:�(�w[���)��qF����1�ε_U�S��i"-	)�,4�<Z��J�RY~#^Mݯ�|���7,�6�*�t��D/v�V6J��H��b8��h[��MQf$���f���>�J����-Sl��G�c�����&�b8�jKC��y��&)*��<�hY�k�A Fg6�E�{l�{��~����^�W( E'�L��<f�>r�&�}�m)9hJw<;ij�4�чF�[�zu��#�ށ:�Q�;<����in0�Ws��ް\n=�_�����?��4ALNY����8)�����_���m!?�1:�����non�Y)�о�8O8I6�^�Ѳ�����U��3:���:�2�{�a<8=�S*�ǓF�5�Na��>C�\P�i���o�pa�k������6�= ���;��Ɵ����Kv���E��<�܋�|�6.�`R�F|�[^=��7�5c��ב&����N���y����݈�EE�4jkM\x��<��M^O+��J����d���n�l�㮓<a�Mb��d�%10�����XL�����Л�*�V��;�}{o�;@'PQ�V�^�^�����SL9���Z�Z���yg�{�ef���3*�$�(Rm��U�=p��"jX�|}'y�łP�U�(���P.�^|u�W��#"j1T��o`2�{!�,�>/7p���z���S2��8x"�Ր�xC��X+��f�=S[T�ϰ�l��}������/���������G��<�vG��$ �33����-�l���I\�wU��L��z�|�����oz����GP�L�u��3Wp,��gr��u��,����I�������A��pd�eh����C��[�����k(�k1���Z��g��^��	 ��M8��4�'o��?�$�'�k�K� ^������i��������8t�g�x���^@�gyo��X_\'�'�O=i�m?x�*<eM�r�#�P���;=��I'T�12ZYF�?;�o�^�A �Ⱥ����\*7���^��A�,&��L� ���>F��\*���+��]��ĭ�T����SIk�W)����4E�ng�]��s�������v��L�(y�J��:���&^|��и�Q ���o�N��dv`U�E�D�%��Q���c��Zĕ��p��q<:�Vk� / P�p��4��T�����K�*�b=K�E�@k�9������X�����3k�O�WB�S5����XT,�6b��������	"7���5�i��M��~��B��<�t�F�!#�V��7�|�ST���D�:��ٲL��:�5��^O��٪+m�4�pK��*3�L�Hz�#M�%�MDhx�a7��>-��KK�/6�<}Ł�,�3��j��X���{��D���u�-����3|�@*���u�Z��\{�a�Ϻ�J�y+%���ڰ��DhOh�j�k�YN�U��r��w6�`�ҏ�Q��qv��S�II��j�����E�׶����("N�҄��1M���
����M`.J)�I*k%n=i����nKr=f�9Ǎ�Z%+=�J�d�=����E��n-"H�0Ƈx"��������^�N�e���e����ѥT���\Z��7�S'O��_�"�ZU˄����j%�D�nR�d���4�xU�h�xq�:�*��{yK�zue��<��J��O�$-�r�B$ڍV'n�i�]�@0�2���חO��I>��*۪���u���$?�o��>�s�2���Kh�+X_����׈���! ��L���G[|&�Z��?����y=y��$Qw���8��@ci/���Pzᇘ�fqۉ{P�g�L�W%�j��l���u��ErX�O#�[���rl�LN��ă�C+1=��8�U%c/�"�Q�W�Mv�z�ɓ&x4f�,]�alx%���w�ͳ$�7tR:c�:���K��RF-I���1������K���NII3j�pZ�୆�٫�#��mT��E2A;��?ϡ'�:�k�$3�c3܃S��ב�/�26���y�	�q~�{#������5��l5���Qĥ�u�[m�9�7Ĕ%Ք��x��kYc����t����9�!��'Ҹ��#����
�[5�x��"#d�N������?�$�¡�7���v�{�>n�'y����``��2�}_������u?u�x��?��w���4�+���**�f�&�C�(��AN�._�}��	޳��	k�{�Pۨȃ���3���ί��#H3b�����X#~9E%�H�E��ϡV��<>��#���(#N��D�WFDF]Q�Ϟ��f�<ǳ�\��GNZ%I	�d��h�ǽ���&�5���~n;����[U��k2WfF���+�g'i|M��w��[������omk���1'TC�a�^�$GIbM*��LJ�vmSN�FS��ј~�����V�����|Ȕc}y#Vn5u��u湒BXtƙ7'��I�s��R�Q��LH��t4�>{*�ձ��]�Y��L��kU	�Q��7Ϡ����>�3���8�m\�r���2�j�6*�ݏ���ηZka}{�w
��}W�������!>�qz�{4Z4�w0-X`�eG��Rx�`���T��Z
=p G S�#rQ�RH/1�뛺F��;�ce󾣽	`F=d�tฯ�#E����G%����ݳ�G�`O�?����������q�&��1������� �2���ġ!�\&�P#���	�c�����x������)�r������ʛ�6��2�se��2�꿋3a�tn���#/�;�*��?�i1��)��Y~�ީ g����pB*�em��ek61��5��������2t��� �fBdšd۴]"��Ӗ�i�t~<s�鳊O�F��6��� 7��!%L����k���@�m��X��rs�������O����L�O���=�`0����hjM��xoD�6$�f��4�E�ڞ�L�i3��U��6+x���`��y�$�a�/K���������� Ko�7�,�=�߇��y����\�d����!��.	dh�Z6Z:���T�u=r�~�E������$�7y��\�_�<���*+�&U +�m������g?�����?��S���5�O����Y�61�d�k�T,�s�"����"׽�.�H����X�y&��������'�����,��ocPna�{bI���G����N�5�'� ��.�L㝎wZ'��2κ���V�l�P�p�#�����.��R�J�g���穽5�3�"�Y����:���I��ƆD��p:�S^�����~��y����������;��'�R&o��m����3�6 S����_A�>D�dz�
��9o�V&�Lx&����z�ф�>�X?a�	��(W5R�Y�^�#]�#�=����bvj�Rpl�&�K���b�L���=w���/����Rj�0k�kC?&�6z���W�4���ZŽGh���+q�̲��w�s�`ZD��mŗ�ꙗq�B�b�ד���cp���.5�P�4�ɳY����p�b	���b-O&L���$�*�.^]���6���.f+���(�0J5�,����h� &qǩ[�ؽ���򰦟"#
�]��P�g���>^���n�`��kQ�Y��P�F����%�dϨR$|��5�����O'���)^E��г�9�?�ʚ�$Լ��&�(��hU"�e�yMr��4"�f��{G=.*��~jtc%E��:��$���|�Y��~>���р�˪�,�8���,�z�t��Hef�<���n��h|Y'�J�a"��ԗ(-N�3�bd�����:U��ޑ�R�]l�-��	8�<�}�	�]�f�1&�K*g��LV�gT�M9q���kW����5?`=w*'D<�B�{��]?XDh�N�%��eG%.�뻒���,{8�rO�߿y���8���p�'�Uh�{k��pThO�����7�l���^T����}��	M��g��M���5�H����o(��B�$�_�s�d�v9>��l���bfJ�+��Y��]��S�[�rm�xD���
A�K�*�Y�&m�~� �7�ԟj�$Q�ҴzE���:�L�E��R���݀ � $��1O���{<�	W��� �>g����n�z0X&�h��搛|�A&j��1FM�CJ2j�۩���Tћx��RkV��m	2�:�G��z���Z ��z�i+2R;�)Ӂ3	��z��o�Z	��_�O�<������_�\ōU��[$�[:w����%(�=�Jf�,��?G�M&׸��V˕�DR-M����;?x�G�EM�j�ۢ���x�]�V�2ŝN׈���5�Foc]~��o��1MN�[6�Qo�33p���hX�`��4��+WP�gUy˗.��t���g�wZ�s	�C��(
��UQ�ٍ|�?|�`��l:����V�[ o��{OC7�J�1E`1A`j�܉<���}�@����E6�n*�E�(&�C:�z�q�`ےQ7�'�qҵ���_Z�J1�7e�4�#�>w��ʐ*q����򥳯���
05���;5��-����=co�d�H�;}G��ѳ�mBZ��TL�89�T�m�Pc 2���6	F0q�<F���S_���&m��W�d݂^�}1�ZЌ�эd�P���U�DOυ��FJ���c�A�찦���*!f�o-�]�z�-���j����2��Tr�f�Y��>�;N1��5ifR�`�d�{�LVU�ipqɥ�W0�C���%cRH%�q�m	\Z9��z��|.makk
��,
ӷY*�]'�������|��$;�῕�t��O���D��Y������C͞+��x��%l�f,%t�l��9�E9B�F�8��E���4X~s3S����ǽ���������{��ޓ�������{����MM��u�+�w{���-���hx��X�AQֲը����-�W^e8��KR�j���"��}�V��I�RDO�p� 4,)n�x���m���1�H/TXet\�;�-�p�N��?gL��0�	�fr�z<���VOe���&D��҈4%�޿�y���&�!뽌�Lz4��U����g�2$z����u��m�=��KK4v>�O�av��5ޟ�r�~�;fL��ưX�z`��F��]��	7p�Y�q�q�6_Å�P�Kc*��R����aj!��p���4���&#�+�7���Ufu�t�5�b�X���^�kGvMhȅ5��=�������jX�}WY����n�{\��_�_�CÀj�v�r����ΎJ��;4���%�n����`�������	=��y
�Ys�TZ�zC���S�f5/�b4��V�ƹ�2�q]e;��^w8�2vʢI�H�[���L\���p{�&�R���aX�J����fWY��M�y��o�Ìti:t<�	��2-��Tv&�w��I���-uq�%�='��}�ت[�.4�"rj�@U��?��k�hjX?Rk��&j�E��N�wT,5��~^�S7�|�,��^D�g�m�b���T	.��.��K4.�G� ���&Vg_��Ƈ?�)�?����+�00�" �ĺ@����<i���Zo�rڲ��~�{��<�z����]��kq��29��|��O����~�\_��?|[�2m:�m<�[�w�y;���\���z���J�޶�IбOMO��[o��[��	����A��gp����>�)<��3�DP���LF;�o��}[N70������<&�&��_�?�Z]F0G?���P*����Y碨F��j��M{�NM�(A������>�l��^���
�e�Ta�p"�=�W���M�7d%O��y!W��R�!.�!UW0���{{^�J�6��u��N��
�E���\	�g�{�~��=�����_[��}ܶ�2]����?~n9�ώ��f��ųV�����+amZ�h
�A̲z5�b���r$������{	"�!�m-Q	D:<��_Q�_��Ӧh ˋ�m�#%
��ӻ�G��x ͷ�8���H���d&��?�Q�ﮓ� �u%u�ǡ-ۭ��h� �2��l�a���z�F��z/�l����GưZ��O�S��|�ʳx?�t�z��V��׻��O$�?|m�������0?���gꨗ_���q,�?l�UZ�PO�x�|\��:ʛ��m�#��"!JT�S%�2��DX$d�j�Z�z[n?~�=x?R���4]���e�Fik=��K6�H�R�697T=0��C*���9��i@>��,�<<��+_ķ^xo_YfԒ2����^I
����!�>zm�9�gE��z|τz�i�yp��a��)�h��U[�L��F�+��eք��nI���شW*T�]��liW�o5�(���l4�dI�/���w�+#p�Fb�֢�~�A�!�Y��������,65���@|m=���������ʯblb��+�g��4��W�����1�,}U�Y������F��Tdx�}�.F-�x��+X�2��X�4� �:t;Ǐ�7k`����kP�^��p7���5�����Vj�Lב+��{2k7G�{��ݢ���G4@�\k{~~�kϏ�����}�b�ݟ��Fe��!n w�Hhy�FO��:� ��a����|��y
�}��g�g��	�M{�h������P� M�o�k��t�D��x:j=pڡ=s0 �s�?&J	e� w-K!�سis�?��0C��u3�z,�H.Z�f8fX�2-:�Z0�u�N���``j)5����ٶ�'��߉����c+�Y�,p��T6b��ܠ�����t`�h����GUe�:O������bS�߾S������t6g�)�R��*G�L'[æ�d6�����&׷���|��G<ß����gr,��d��Qd�Tr���Ǘ��8����w�A����qD�{S&�p��x�O�K�&k�=�p�2��t
[�:�Q��6�&F]� ���<���9L�u���o�3�Y����쯔��R�P�7���cb�kǉ�}x�7�P����!��#���������PF����� 35�"��@�@�&~��M���	���rջ,�MU4�)�� U��O۽�����ô��4T�@���J�_S�J}�z�q�nM��������#q�+� �l�p`MY.�v�YY���QǥZL˗~P���P�� o�GMYؾ%VӁUB.PU��U$�ج�*&i,��K%���0�e�$#gmS�k��*�gQ���u�k���pFR�[<���y�?��SO}H�@*�lo҆K�(+�!�pf�y����g4N�j����j2p��
�������OL���8�*������Z���8��	�E�g��嘒o���a��(�����=�e(�(7E���Я������~��d.�����0�	��bn.�\a�{�26W/�{���1h�pw�/W�,��|I.d�^����tSt�Q%t�)��,�<��<�ΛƇ}L�l���!J{�����{�x?/�7|����FӴ�^��G�!�'�;��h5�6%�Ç��$�����M%�I5���pt����+���1c���67���4��;}U=��p��@�)0�PKa��ݳ,��ne���2�W��/*��
��t�xܔ�lWPK&���/�E��B(5�)��(R-�⹲�\�Jd(�tU ��m�$8���V�2��Ȑ(��焗Bh����C��+�|j��)��r�V�x������M3�2|!M����]�d����[Jt�X�޾�y���Wx�3��,����M�&ğ��1`y������
YLF/�3���F�hR��_��&��j���zv�,Y�;�/p��>aH*=��\�J3���h#�= ntF�d�� DS�6�>iM��ɴ�2��M[z���{�BìB�:0C�p�H�K=@�n�a-�'1E 2�o�Ⱦ0n;�ǭ��03=��M˩46�kt�U:�?*�&��J�F�� �Д*?��iE:OM�j�M:�r���d n����M�^_v��a��i �s���ˮkm"����D瑍b� ��{N
X�S��!�J�}�����,&g�Pl��g0;hV��D�Y�{6.�B�<+F։0���2h?�
i���:���|� Hg�ʥ���?7n ��`.��"�ڕb��bʞp}[�Nӓ�&ik2�!��J�d�_:�4�;<�C��eck���ߛ�X6e�ؒ�S���67�x�;��{_������w�w���?�;N�o:���Q<��'Q�FC�EV]f��5D��ǓO����9�ퟬqm��X�^Ǳ���c������.3�̗"Y5��I���i��U$�K8�VÓ�)��q\~�^�^F��>����e�0���Ҙ�����
�:�<����Z���Ak�ɧr���������0Ѵe�z*���B�l~�j���2��������C���>Hr6%����{��Y�Y�	�(��A�n�:ƽ��T��秸's&��_�����Z�b�����D��S��zvu���:���U�G�zĚ}y��h���^���x*e�U�j��hRB�-'B��`9��/�8�:�����FK6��@��|r�F���#J�;�-�F_�%��gU��v]C!T4(��N�>���D��6���m��q��p�L�{���[@;7�E�>����~��t�I����ًQ���f?M�o�w��T�����>K���9ۆ=���K2p��#��[g�W���T�AHT�G��'�q|����sx��46���O��ܕkX�����4�;�u�!dT�<v#�S��+bf����7�g<�j��u��;kXݢQٮ;:�~�ʳ��}՘����?��⮓G���X��2�EVb�7��R������~��ߑ[[&���0���۶iJ�m�sx�	�e�d�m&��8pL�a�Y��������W�f�l~UO��m4)����AFU9�G~zh5ͱF�K�<�S|�WPWv��'��a�ZV�� @���iz6?>�ka���h����$Y(�2=X�cu��<d�0�YGzk����縍4���l%��,E�LP6�R/f�\6�+3#�k��a���ѐ�O���_؇&����y�j�Q�7�یrb�fO�z���/nv0{�����%p���P��5��}����ֽ���a�+-�\���;��^CI�з��`4��`���.Y����i��Q��0�r�5{��l��d����{b�W�/mVݵ�,�US>���$3��@j��I�����O����O�б)�Ƨ\�~�b���Yo��_&�}K�a��������3*=)��J��grH�
���N<vW�&G�v��{���y�q���l?ba�7�1��^-:�8������EHl�s�cz=4x>��n<z�D���ndx��7�r��|��z��<���beiŪ��gƳ�k��k�_�q��p�������e}��k�� O��M2��޴�Z1�����6B}���I[�h|�	���a%f{�g����csy����xxs�h�*|�(uzX�U44-��+?@ce�G��W��B�p!t��O�?H�CsX	��2Lm�yM��yV~���u�:"H.]8����<j��dF��U�F�^3I�T:�������5��~+Ͽ�O<�<AJ�V���U\�v	�$��->��P�T�e��J���Ε�\��d�W7�7~��t��e�kU\T���^*P�ƌ|X��2���(���^��0�>y��UF1%��,R�I�:ۄ;�]Vv�/�J~�f+PKP^��14hۺ��WIS0�i�V �;��L&���q��Zp�ӯ��j���kU�T6���6�#ʝ8�'/�2%��>9�g�����NI�Z����L��0�fL��8��`��љT�1�U7�\�����",)Á�{��6W0hK�"�\j��:|V�����F?� ��uCAa�
�.HJBՍU����G�H���"���ʷ��%[x;U�ݏ�-0�k:�ylϽ�ɉ�L�ח���ࣷ��!�U�1V�`u���R�S���e�1����yR7�Xy{�p�"�cqc���o��o�Fa�uQ�X�aj[�ڵ&&cy<r�Q��_p��;9������b�O�0-]>d�փ��Z��ұ7#��ף))�t�w�8�O<|֗�Ca*��<��ֹVD�s�n�Ux��"$��]h�i�{������G��X��bՖ�q��vxԠ�9iT?�T���*����������g��jt��1>6�l��ܔ���5��fSV��U�h��+�GD��*����oRv��IF=�/&�R�(jj�
:��u ��[���I�����ţ=�C������v2h�<:l(�m�F��iE��_���Hf�p��I��M��p��R��������T)�Lʈ?�il�Ty�d�@a=��b� 7D�LG�����:�By_eI})s�;%��ˠY�r��!�S@��M�+GGJ���ێ��H�oh�C��^�auz������)n�nW&j�ZáF���ܟa7]<���{����=��7��`*��H��1b�q3�����N��ȃc]G\Z�����6j���I���uVn�s�S�X�r1A�sH�v^�����ENػ�\&b��$���"�9�^$�8�$��J.������	��,�G�&�Y�z�d�m� �����_�"������<�.�=G��pcq��8XHa��5�g�"�20i��P��*5�u����΍���6	.rhi}�FW�i�')K(��}�&(E��$���h �o�:?&lb�@�w'N[DE�S�����(�71A�����i{�=Mƪ,�ų�)|}N�������Ugqt�-�c9ԫ}\|}�8�x��sx���=�݋t6�{k9�?�~�?����g��x<=��J�����}������?��g���_�59r�2h�b���q<�̫��Ul�u�o��7� 04��d�`0�����q��ILƉiZ��n�4�L;�� ��+x��8����J6�}&pE�6��,���k,��R���?f������-t7���͙.������sܵshb�N���gE�����2�n�47��9�oR�.�U	[%�h��F�U?{���ِ��e�?��t�(��͆�W�J�����7�T��}e�J������|���v��e�՗'��T�v���prD�d#UVP�9?���s�
~���z�D6O�0�6^؉�>6KU�ڋv
}���D���.�_1 �3.P�u�;�C�߃|��쵟7`�s��ͨ�?����68`����cӨ�{�<z��e��?z��2�@��7/.3x�`j~
�����l���]�Q1 �8��{�;jP�� z�P'����)r���<�c�?s��]�כX���ҕ,/w���p��9�\Ϧ6C��ݍ[�����>�����F�����)��Y����ި�$ �3��'>�d�n�{�Oᥗ.௾����4�-��#�Ԥ�?蚢���~i�`'�~:��$���X�C�)M]���r_��}���F # ���%MC,ф$�.��/<x���μ��?��i=��InɌ�����K��2#'����f��C��e,�/�-��h4��Q,�]:/5��ߞ}�i��m(��ѵ����r�t�&���������ƽ�w����߷�T�.��sLy�qo#Yz��}�����Xr_j���.�7QbS�DiHqf�3�F0<O��^�d��O�� �!cنmcs �%Q��El���[uUמU�gFFƾ/�^���7����ET7�DWeeF����?�;����gI��T;A^Q@���<������X�!��8"�RD9���H.��\��
ET�ؼw�����A��a+��={}+��Y'�)é��ZZ�6���������ό���8蘁1?��y��f��g�L�I�;��翅=Ӄƌ����4��N0z�&�i����?����;"?�`2���x��²�,d��8�>�9�ЖCza�� )�+�T=S��f�%�z��I�Vkk�99��.5�T�|B�P��CAɎ���1��?�� Z��e��gf��$���l�5��05L�+[H�QL�d� ��m
Phu;ڸ<a���{���w���BkPW�_o�`e�f��x�un�H0$AQ2-@��������rHfMA9�~���!%��u::e����wY�L���W�^�fǌ�Gq!͈r���cm1�Me�<S/�KF�Z��'��/@������-�/�7��?ĥg.i��*,L��1���&�ߔxa����w�{|�;v�RA9ǝc�|��w��K��by�l��PKב��tr��n!�������×1�u'����P����YP���*2K{֞;����������p�1t�	�$a�������ӟ�|⹫F.mdd�������Cv~�L�x�iAՆ��Ħ���>���������::��}wL 0(!�b��Pp�be�}�$P�c�����ے�4Ocn���7q��	uܧh��
�ZA��ҡW�h�0�;*'6�O1l�Qv`&O��f,��w�F�GDe?��qs�:�$>7TDa�S���sT	�R�<G����fl?�5�6S=PX��v��>̂=��ܥ�~������W���X>��CD����M��8�?���5�3Ofh�@U�#~�W���xF�9��KepV��K(M�O�� ���؇e)�/˺�si<�V�3�)�3e4�c�a���7����?�G_���`3_(�r��bԑ��a�N����G����s�7���ܑ�j'b�Gq���#��2��I?��b�<&w	�z��%�9�.Q�TA�8��n=V���^��N��e�d*��NK���O���C<�w�i�����"V�d�jr�v��x��<���}[�rH�AW��`JJu	�P�y@�8�7IK�̘1
%��j�F�eV��L�7p������^{O3�e�r�c�ě��C.�:��"��S:��� �g�$~�p��{x(ǩ%��-Tۓ=��~O�����h��)��
��q��C��l$���B��L�9�6��
sZ ��"�X���Vi���l��Z�F��>�h��X�~��"���@e��2B<��J^{6���4�_�H"*���g��M�se�BK�#�-� ��a}�7�[������Њxh	P��8�+{�KP,ّq�T!c��6�+�keS�Ņ�ɗ*!�Q_�C4�� ����c�,�'f8A�!:�i	�y�$���5!��&	kٴ�P&.�9+?�{���&[vʗ�Cy!�|6�\:$�8����9G��Cق�M��hBQ,�-Y�z����`U��������X��M��c0@���|K%ی! ������L����,V8�VQ�{G�5'�)>" '��!���e�0���1��WA)�Uef�9�A�'}V�y�TL-����k�N��D��.{��W���@�mw!�b&��!L%P�LO��bY�h�5�E���r��\�����}R����z��w�`Z)�C�x��2��A|���1����HجW(� &��e&=�~{�w߹�>u�9��c1�a	���Pʧq�}�w��cW �f��ww�bPL����`���������GφCT��:vx��S8�������������C�}�~鋟����ƭ�r�*jI�)If�/�Cj�,<ܿ�{�s8~���� ���Y����������[F����|��� '���{������<3dH��[Ԡ�� z��)�����5S��8%�8dC@��_��>UhJ1�IaҪ*�L���4:�R7R81x��t���f��е���ё:9y�$FN\rH*�/��6F ����o��;�2b:�d�~�p�-���2�(�ir܉/�o˙l!^^@:#��|K�l��>b��̆5��G��nЗ�vk����_gL9��!,�%���rڗT�$QƓ�8CĢ'XZ�q�B�<�A6g@V�����66�ڨ�ؾ�q}�{S�[$�o�o�YL��>�R��Z�d���������Vix��O=���q���m����3�e�N�1�!���|�Yl�\�����u7���9\���7���._\���<����\����13���i�s���'��|��q�|��=���|�hv�)��Nd4c��eya]6k������}J߀�8���C1=\ܴO�L4���y�Ϛy����¿�w�����?���D,��p�l��)mɠ�%!�� ��N0����㈹�J���t��@vN����B$ҍ�����o~��\C�P�N�N}���|�y��Ɋ[ց6��g�Y�CO�6X:��֝;�?�j9�fwj�;Yje��x�>w�E|���ə�	d:V�����֐|�cᔀ`I�%QG��{<�f�r�i�?I;'�|�QC�Q��qT�bqi^��s����e<����nc��,�3�%�vB�\��c41Q��p.AY]��X{n�w�nb"ηQk�n�3R=�A��4��ݾ8����H��Xօ*l����7}�'�<'Д�j%'�',ׄ=30�3z��L�/�$f�gb���=���$�%mH.m#��Oa>���D����'zX��d�=ia�!��q�Q�� �L)�|)��b
qY�즒�Q3A�R�N��s�ۭ�Ѫ4Q?�C�
���3�d���g���@wʌ�Ф$'���{GV ��2ql��s���cۄ��/Ϛeɟ,�0�O��~�U0/��j!������]]cCQGt��+�x��E�4yV=6�+�o�։����@�v5*.�J�8�&{�%�"�=J�$���ߩ�9���ߌ�0'��^('���[�Wֽ%vSv�-��㩋��} ��(E���&��'+�2?��L���w��a�����$0x�{���ݛ�q�����	��y̔
c��ݝ-��p'|��wq��!�hpr ob��_�##�$���rfg�Gk�K(K ����{�XZ�:޹�r��8��\{�;x�����>^����u}3~��'C�m�cw��v��7��G|��[�S�=f��Z횀[_���ۚ��ʺ�'���.�Nۃ�o��h�\i�l�Xk�+�A`���-����e��d���?;��T 4�6�i|����%a�2�~�V��5y�mOd�W�5��W92�1x���%x��7��)��x�LPB�����_�{t�-��� W@���?�ܤ!퉘�#���G�kk֜U Ol�S��������������d\�T�{�ϰ��Q�Dl>ⲏ,̯$�V�╫�R�S�M�qg�� ��1��;ح$��3:8e���>�d�I_�НҶ�F�ӛ��%�����#�Ol�������8��}� ������?����t��p�#�{F��}�Gm�-9;CD���<y�9bD0��5��F�hH����c:�ʆ��� ��"�|CsX<4ģ���������^���9���fd�� Z��,��eG֫��o����Iԇ�\*x��;-�22�!chxY$�$��3�2�g�:%�����x&�GA<�' #)4uqX�aQ�Z{~�)9X+O����M\���Js1��S�NP�$Q�/#/>\�aW6�_7wPKʚ��H��S>H��^��k�G��+`��I�pXgq�}��������`�ղN#A;�M}mv�������EM��%��cz�HȭM����iP�\+�Y�Q9`te�P�R�r��
6o�����w��s���,��L��
 vd�j5&�U 2	��).���\��p.6��4�3�]�C5�h���?+���ڳC�>��Y�}���O����.���!C�CC��mA��6��6����,푍�����LD-���Q�҅������U���C�$��n&�{�2Y�{�lQA�Q�j�BF�X5S-3�b)ǣ8�j��4�bt��8#�ti����v;r_}y�Tg�����c@���(k��>T�z:����ΐff),�R��2|u�������uЬuqҬb�$��� �	�T(jp�R�P�'e�rB��ˋ%�ySf�H$s:)�롃�$":Y9��3k;5�̽�H9u[^,������m�7�c�wz#�!ݺ��ϯ.��F�;'��x?�d�W@9{1N�0K��a�pf➣L�5� �L�������"Hm�j�lfJ��[�*��p�cP���w�aS@o�!�Y�Qg���n�g��{�:r����&p�P,�� s$��k��?h�a^������7oɳh� )rHJO�ʽ���L&��rE���7��v�����q8D���װ-�Hr��
��5Φ���}��w�~�(�r��ؼ}����'u,��L�3B�V�>��YG�eɱH*�_��$t�Y�e19K)�x^���x�� 2�"q�R_�@�!�2�-�m�>9Bi������V�O-���06���V��i"�Wf�����H�'|tH�V�@�M�	�eϲ�ٚ���.�L��^l6��
�8umOرgt f���F��!ŔhI�e��Q�9}���'z}��E�=��$I���;�
�*�zDt�(N�����{i�/���W�LYȐIy1y�z����4"��<���8x�V������e����?�������Gqx2En!�Z�?���x��ە:�|�5����xpg㡍��ed�����:�sד��|r�b<�aj���㶢�pd�D����"�mN[6WO"Ĩn8�O�Or���.���M�����5C�,�i4�hK��@�.h��3�4z����٧e�,|���ڹ�tyN�O�(� ����g4N<� ��|���i�:�`��BR~�V6p.��CE!/N)2��;����k���'�(^� �����u�Q��p��q,E\��2�&��$�ᵚH��V6�Yy֋blz,i�#�i�T��|5��_������{�埓?��.����̖�x!O�E���
�r��K���=����x�SG��J�01S��#�����jm�]��Z��h<��e\��*6V�`�x�nN������Rq�TNd��CD։���nK� �D�:����.�Q�'��#�+�c�#c�w궺
p��bD�Gf8�,-M���H�N�E� 5TU=$F���@K3��=W��e\~�̑ 5��i?X8ji_'�9�%Չq��e��a�EcN .�D��cfAVc�W�@f&R���g����:�7�UJ�{��3x��%	dj:����� q6��$6U�a+g�9: EQu_�T>�E ��瘆v��y,C3}LI�	����6�i\>��k��V��q�p �/Y��ڊ������-�Mc�-���S��,<u�<2r�X����t����{��h���:�>u��f��M�W��Ӓ�JN�
�Z�N߽�������h����u�4�s�\��4�zG��1��g�'88*��u�w|?���5g;E\�D���%NG��Q��Ao�cd����#�%��u�h�Ƙ+g�l��uU��/�R��tj��R���|���f�c�4�n����
n	PS�@Y��bY�/X���	�93���{��J�4�k���r�-,��@D���l/��<>����wޑ3�ƅq��+�p�}M�/��]�ױw|��?A9>�=�Fgz�b�TJ R#���m0���9=Jh�	[K��:S�i��p���k�cV�D��G�=G������xZ��-Ι���]�.���n����*�{F#��I����c<�r�&���	�ꉭ����{0�}~��R�j=h���٩��i[��h?�E��)ɳ�6\)��GYF%T���^���v�6��5��������mB��Ȉɻ�~ď��yH���^���"��<����ڭ�N>Î�x��c7�l;�G����L"s��ĒY4d��ۨ�#��c�3H�zuQ�`�ӗ�5��Js�n<�s�n�(�n"BW��R}�'��Z����\��F��㊦$��X:��Zm�Ġ��e�2:wy�vY6ɼ�K2��v������Xk�)�ڧ�?���ɫ����]��b��?=8���q�a'ӈf��VY���n���~�"<Yӭð�o,������|�����S��.P�=���P߱bl\pR�7ň�a�����Y��{̉q>��~�����kx ��^������_���>�9����.
��D�<�5�K��K���E Fo4ƈ�R��Q:���_�"�/����;���G1r�n����a�A[{���̺���8�4�Vn�����Q4<�Đ\.7�z���t���c��+�˟:iWj\�XDF���Wֱ"Q�T Z$:���y��WD�u��4��W{>>��@�1Dz��D.��*��f���n��#�|�s)Hhn�oa��Ǧ�0<y^1f�(�&���i>���H
*N�l6hs�X%��xgC�f�|�HY�:�8�Yf�?��D���5YѸҼ(Τ��ɖ)`c=7�4�yN��A��\e���GfO���X$�㞍����v�NC@]�N�{�ܢ�Uٲ��s9��������]4Ũs�����3�(UBqL�F�J�cJ֧Y��|p���'�F̊�eo&RYy%BM:\8{�fw��øG:c�|p�'���tї )bE�r����Gb<e��(��p���HΕ��#�pY
c�H�A蜨��sH3{�̎ŁR��yܳ�DX�b�ܹ�@K��\[3���c�G(����{��IE%q�Yw�w��I�rk�{kH�aV��%Y�~O Q1��5�>zSj�$�cC��L.��'c�8I�p��I}��{�-��,$�r��g�h�Q�B�|�C=�j��N�O�X��zՐ�ʚ�bܱz�L"gd-C�&T�yڞ ����i�;p�}�MJ0�_;��r��;��+U�u`���x�{��we�mD��CY�1-k>�5t���������\t$�5'�:�T��wh�˩@��o�^Ee�G�#���+Ј�ϣ�	�G�*�[b�@Ӳ�{�b��ᮬ`���"�R6qj"O�DS �-*��Zh�`/�:d�@�Rv���e�pa�r?��З��n��v�H[=�:{l�P.-jM�<���V%[�v)�H�G�2�@�>��l��r�m�f&�$�oz��O�J��6Jɭ�Y��mӎb 0m�;㾱�Xrn��R��B!9C�1����3��q��S�M��V����HΘ<ɐ ʓU-����e[?��ҁ�'�n�\kA�Դ��s0��{�g>�j�YK��}�%�U�AǏ����7�+��~$��khnt��{�a}um��?��[JI���˸�`;�8���Y�'�S����0�Y��4� rc��	����2���F���1=|e�ݏS��&d�C��� T��ʡf"/+84?��^�����)rI\���7���X.���_�ȏ�_���ދi�۝B�>G�-�zo�'$n6���'�6���ځW��AT �0I�$�&��8�"y���ߨ	��ŉK1p��lH$��x�o�PCl��L��hl�&����<�����/�����쯾�e�� V�2�r$ ����Bi1����T ���z����#�:�hT��z]�{��,�i㩯��
�A�$\��l��:A�ˤ���b���^��tV�|�~	{˸xo�����-�:t+Q�]���WVK�d�(yl*��F��)>Okql�|!�h��V�]^�Ƶtv��c���Ơ�0�U�u�VF��=85L�D~ݾ���3���Dm@���N�G"úL-�$�d�cziH֪�,��ڍz���TC�\yΖ hj���&�,���xՙfr[i_�8�Z��aw�a���Zy[ۨ<�!��ϟA�( H�5�1�uT�)���B�u��%�C2��d�3�O81��e5}��F��ɠ�I��V��MZxx�6�)}8L}\8��$�$�m6���$޼��Db��_���@ *)��?���ϪrB83�\�<`�T��{�C:)�r4Pa���NʿgsN@	}�>��GJ���ʒqc���|��׾��py?fU���a"�1�!��o?�(��KimM�8ڟe��Fí�$l�̘���>,��Ъگ�Л��@�s_@Ǵ��j>��k��z%�d%��	��z8��)�����i	Ƚ7L�����ru�������O>�}��8~�w2�G@-Q[��V��&A� ��|�������QM�m#5��֎�sN�����|��V������l%���{��\����t�l��2�\{���3�v��$h?����J������5��רy�H��4���bHd�%s���ݛ:Qy���� GԆ�=�DMH8#yD�@���Ɲɠi�ӏ�.��Q|�֣�G��:�����X���T\��xW?ତ��!�P������������F�Sm�,3nz�&z6gr����ه�	PVf�&�*N�^B�s�}q�ۑ��!���RN�Z���#;�QJ��3X�y�cE���e��leE��)EFV����><�X�B&%�&)�B�߯��=m��-۶]K���G���HLOƈ�PQ�9�a1>Q_7�5e3wT?�SKjx���xlHIa�?��d�~��gӳ��L�pj*�/ ��k&�g>	͆g���x|�j�_����q��M�� �5��D�wd)����H��6����q����y}$X
���S�zN":��̏����>EI"d�Mc .�e&B�����/�$F4��woI�¥˗����v��%4�5���w������9-y��ƌ{����C�����i�e����R�=�6d9Њ��Dm���{�����N�쵴A�C'�u�����I���ѕH���'4��L���U��S<�%�������o�'��є�\k��xX(H������K�$Bcme�c�o�2�iz2
w��W3�9u8���f���T7�f��@jE��}��˾ɰ}8���c��IA������i�NS���#{�G	����2���p�Ku���gK{^��H>��	�:�� 6Y�~�������������cu��XIaa}Iq�y�|n�3�p����iO����i�� ����J� 42Y`N�N�w{����`2��4��^�)���\�t��*�w��s��{�ʢf՛uW��o�_,#����/���ª�Ǹ�ф�����"� ������R ��k֊Y=�D��pٹj;YF+�������B�����/�ݭ#	:���c=?v�A\��[(@�z�Hb �[���u��R'ڗsͫe�����D˵t�F��Wpc����k=mG��y\^YD�W�T1�ўX�9y��f���hXm[*ؖ0�O4#E'��獵���$+��fٯ<�&
��r���J�30��t���oW���!9
Tȵw��|�Ͼ���M��⋲�.�̚O�.��ˋ�,���VY�}	��Ø]W�q�4և�gԒe`�Yŀ�*7�0ȹ��Md��N�z�ޤ)g�
+�	;�,	y���C	����c���nM��yQ1iٻ	%rYc$��@�-���	"�
��J���Ry&c�� [��$�?����4��4h�r�Gr}ݚ����`8���+u�1��̧g��@�̩-ar�s��1#��,^�+���0�Ùj��
�A��e?Nm9�o}_�`9�l��g�Z�zk��^���^���h8J��E�w3`�\U9���I���A�#�%��U^V9�:y�ʝq�0S!�����q-�ʶFW@�=m+=���?��M,.M��V�G:����v�J���Ρ��%p���䍆}M���C������y?%v5��J��B��S/ޣ��^�O����g��l�G����lHV�#�%�3�tq�d3�d�C��X_ܻ����� 5/F����/!�8�q��?��kh�h���� dz��5�J��<UG�]��A���V?�]}h������*u2���	x#9(�B���h�T�z�>ܒ��i:��%d2)��CXX�8��;��bumg��p������ZMU94�C�`C)3>JMM��H}.�!�Ű};hr�5#C�ɒX"����.ΡX�W����aC���{2B��5���b�����sk8����_{���YK"��k(�Cx�'�]�7�İ��%F�n���8յ�(V�8���r9�R.�b.�d�G���K����VI�p�'b�\�Ϧ�tzj�|��U�<��d�܂��,3IM�'k�~����N��@4�i�s�G�s%	�\�aض佦c�a�h���쭉!HU/��y@!�N,E�?U�͌mWr��	���<�!U���댱]m�՛����:p��:���H�0�5r����>��џ(�">AI�ڬG�Ht�3�A��%�/A��W��)XHɞ'�/���c�\ ���h�ڲ}��كSTc��䭭�`����Q�W^�>� �ڇ�za�d�:�!Kg[m�K8��Q}��l�Hv$�! s3n(+�ypd{��k1[����l˶���wk��=��0?SzO����49��4݀�L'ByV�4��f��u��U,�Z��*:c��Z���W1щ���8���X>n��3I�&���9�c�#?3(hTN�	�+Ob�S�y[�ج �d܍F��6�YQr,ZS�ec#2�<	�Bb{��#�Ǿ~�^�������q�����;��;ȤR��?�x�r�N�*t$�P=��I����o$y��cO,uk}C8��(�?h���?�,�#`�#�rh�N��˞��y{����݌qr��)�K��p�|\(�r�'��p�0:E2�A��P�^	ٹ��0ڲ�]mc�l�j���PL�C4�$ƙ�Vsl'%v�U�rz۞����g]#eG��S�&S��,�� ���%�h�t e� �h�t���O1���4�D�4[I$�1��T|!��\�NϘ��>dzP8���%t�)4)is5�w
`grd]&��ªN���ӵ��o*6�++��ٍJ�ۆ���}_p����9�#��k��nJ0Or�md�`�%wMo�w��t�9�����e1�ql��Eg2t%�cC�D�^L�nJ_٧�Ꮒ��v��*�'�-�Qo�`����E�ã��{Ixx���w���M��i��nF�S����ׂ-�;�>����E*�r4��Sm�k���^Ss�h�I;�$9h��H�5�Q��jxCS���4(*/��I:�ހRS�ſ3��ג.4p��-�&\�X�2�͛7��Z��7��ӗ�c�X���K�ZR�@:�\!{J�I@BP�)@�KE���3���YV�{E�N�q��-�P.��G-�S;��P�?�~����,D!��a��J�����½��(=5�� ���Pf���?W��#�FS��3�l�Z#����qy���t���#H��~-���h�[��$2�f��$d��M@�|��S�h(���:P�*Fo�ms<-JX�0 h��!�iP]��݁?�[�8=U�!�oJ�H��yF_�mԑ��/��������Þ1M��B���w��-q���>�����]L�R<���/�Yxἀ╒XqP������Y�tU��Ӈ^��g�X{H3w*������`�#�����Q +7$Kc\��(Du²M�޷���:���%�p��q�5��:�D�0ݼ��T��X�x
%�֝�c�ܔ�ل�e��)�q�,�[�TЄMMUJ'�y��l�����0C��(����(���m7�h�zr({��T>���.n�G���d�ϮɞK�#g��@}��.b��?���a����l|qp��a�qK&��&�y��=x:�@�7�k�4������n���jE�lh���'mͼp�H����J�B�j��~��eC��5v*d����W�-U#!Ș�\���},�K�(�p���_�~���r�r�s-eW*|��_ś－r�(�؂�!ٟ�uTS��ܫ��{w�ƹl� ���_��R��ca��t~$�&�9{������)���!Ň)��o�|��Íf1�
��dSSQe"���H����i͐��HX��k�#4$�3T�3D�̤��P��q�b��bf��V����;.�G�E�@B���9��������[A��g���$M������� p�Dg@&�V@����Z0�(ƾ�@�����&Ɋm_���Ǣ�B��L[�r�*HrV��P�X$ ��*	9j���a����2����y�L�N�~@oFS��~�(�p�����Zd{�8������-x=|�Q|��TG�_��M	���g�䟉]����רQc!�ƀ���1�9K��;0]=O~�T9Y��H��L2�̓;�r��WSJH���h'��%r�љ��sݚQ�e���H؃��C����MiC��:4t,k|�/���$��]�����[�	�V'��v�J��(s �Y�T�C�L�v1�0=�q�T8_�a��������L�Z&�E�XF���q�����?C��2~e��P��]�gϜ�(yg{�QIri�b��`}e��	�Q,���A��(�ԝ|o#w]L����i$7�g�mȬ����(���?�9�%R��<���C�6h��c�i0�a
�b�b�vfG��9�������I���{�.���v�[D��.�rUb�6�M4��
Ql���9���k("����b!��sy���RQD�}�@S-Z��G�g3��*��2�9��[�����$Z����g�
�&0#c���9Q�Y��`8��<U��L(�75D�$�u�;n)���{C������8��'�7�Pm�Q�8�����1T���G��I˹�@_p|<���'�dp���0��s���Q��T����:0�������X�R"�S���\Y��rY� .!�D�1��Q#V�~d$�e��I����5�V=�ٴN�E�M$1��1��	�k�"1A��<n�v�z��H�Q\=�����$�)��g4V�`�Kwj�z����8I>bvT�k�VW�C�wʘ�%�=��b�o�2����<��NPF��v�����b��Cof��h��AR��R)͐�X����	�ܙ�9�U7�(�=:8�u6 �v�*34b����	L����/�DT�MKi�,���+K��>:�N�z��8�a�� 	@��]�t1�J5��P{{9)k��*�x���l�<����V��گ�u�>�Y/�,�cb�	�H�����/�گ��_�s����>~�󿂌��h"��l���YT����K�����`�I)��W��ɘ)YN���08"ߝ�\	�O���ѡ�-�3����ٖJ����/��� -ʙ�<��˪O�sF���6�}��/���U,��ij��qb�Rr�~X�A_�B��T����P��P�A "�I(+=��+]����f��5��=$����x����(�c�U��`L��<Ʋ��)�I@(ς �-䒴B�V0�洭7��g5�z����U�6��6{��G7�����򁆰{�G��������K⛀���}٨�+�xv����E|�bZ���~q!��n�񋗯�ꋟ�7��{�ڪ��!� �,�����<��c�wX�N��d���T�%��ď�F|l��د�F<���@W�#^�G�d	�)2=�40=A��tu��?��?�7����Yq���)��1`�=G��T�� �6`Hu+�T�t�����1���P k�#��q<�Xq%
N��ˤ�谷G�	�������Rn$�� �~�4	\y�

��fϸ�/?u	��n"?7�+W��տ���e$���Ī\s:�8���S �L�Z��`���?�?�N�� �O)!�����l���=Ff4vĔ��d0����Itr�`��i��_G�f��X�;F��J���
����O����D��Xn
ȕH�a{��p�6A��y���r�nV(g�X*�QH�X�K���ˡ2���tT	�c���8(݆��̀�41Z�vĈQ��P(KՎc�1{0M+�m�c���:�VQ�r,��d��_�71FY�:C� !x��'��W�>	���eCrM	��o$�C�ђ���K�o��!�3d��`R�W�RLM���\�ڸtn�ϔ��9L�(�UPp������BD�7��Ң0�ٷ�6���Y���y:<b�v�	��|�-{�#�LN�[��{�;��^ƾ �所9*i�gq�$�j.�֯�/ k8N(�;KIyv�'5�Z5��c�c!ղ�,	|�1���ٴI"- �SUO�%��_M'me�����@Ya�sإ#gו]7�BB��8�X�1�W�ehy��}>�����=%�էډ�*�o5[��	%Q�E��.��Z� `0
",�N��F�JK��f���_�l%�xZZK���8��������Jɒ��O�&`2LC��J��h�rc�\:/�;AC�A2�P8��53��β����`p�!�t�
g`�Y@gk)	�{��̸�VϞ�g?�Y�(UF9�� <_@�K#�τ|F�Xƺ�����Zrgo6�I\<�33�����3ioq����qUs�Jݍey�&b7��H~KV�9����m[Җ�i�W�C��RleH�5���`�Чΰ؇�#�7^�X���UC/ +ʂ�(%+@V0|�=�<=�(��K�9�����t`��:d�%[~'��딒����p�����3�C���䚩}�в����y�	�ڼ�����~Oɏ�_R���T���2`�2�w��!A�oZ[ȷ�6�Ph6m������G�����v���:��/��K�& ���D|CT�U!�l8/6���<�"�����0�o��o`u��@n.�D-��<�t(�I$]�'d�Ncl�C�Db`�P�X����J����_bO��X]��·w���p�x�|�Wщ�rry�ڛtbU{Y�����I���?ke��<����<^z��Gإ�����z�܉��b���=k�q�T�]@�4�g�z�*�8�da�q_����D�G��2���A�66p��D�`��ѐ�=yY,1%3q�~���u��q\���g�b�#��)�uW%�ڭ��Ʊqٔ�6E_��%�9�h�*x�@Ȍ���i��\!���WQ,/h������������4�k��'8�
􌤚M�g�Pk4q�٧0�\���&j�d���2FR(<�Ͽ�9��=z�@��������ʢ�b��w�Y��rr�8���_�	�+�Q�˂�we���%�ir��k����'!��Q�?���]��	t�܀��"b�z�Yze&�B����`*U@'`YB��fi�t?Q����B81LMԡ|Q�?p'�֛�%�5���L���g��М72Q�o1�Y��Rx�LW>����k����1����o�������@$�� ����ً�X$|�P��Y��~![�ɕ�Rl����f��A.,�A���B���=��������P?ԕl�[M�~a'�6��'�X9��3�FI��˟|N){�S
�g��Sji,g#�׭@e��\�]Q����i����t�@#���`�vN�2�s'�s�Y΁�l�Y%Y%�i4;my�I�$�oU����TN��w�P���'}L���=S��#�HW!җ}!7�6t�$3WC��Z#헌��l�J��ϛ/H *�d��L�  K��ةf_��,���;l٩�Kϩ}��48	��������{�z�3��YNT��d{��ϝ���oba}����������V�}I�3�ӷ�|7o�Rp���|F�76���b�G:����v�%|�ӯ�E����ilX�c&ϊ�e|���C�2���Jr��U]^w�j_(���.�t��|�z�#��	��~���(���YΤJ��fU�v!�4�2�	w�?��h�i2�^7���Ň�<��G
��\�<�����S+Yw<�P���-3��Q�\Ur� �K07&Hu#y��&P���F�Euq(���<K�Cޢ�/�'>ɒ�B�Fͭ��Zݻ$�!�=��}�'�����^L����s��p�9�c�5���&8�������-����g���J����C2Af+�ZB �
�4/��Zl�/~�����s�4��=n��2�ýx����z������~|�G�&k������	��0���J�؊�Z��l�����Np�����%=T������n��p���>R0�V���#�1k�)��h�O�0g�������Cx����r�O���Qm����5����3����i!#����I��`6�d�ߖ�0��)����r<�=1�|�8}��*?W���jQ��z��ٖ������_��|��ҝ�g��T{-=9X������{�xB�zww��h,�����=�����sp�)�PM��=��é�*	,�⸲�����щV���A��Yf�Eu ��P��(q���*֊�:(�y����X7{f�����&����$�ثI��P�b��y-��l�PP��'⍈��H$�KO������5����
 �S�#�I{���Y�	H��X
��]�jś�JǑ�ߣ�k�rR�i ��(��%��<_*�6�����R��CT��1�%�6�]��8���8!Fq����-�����MT����q3�*kJQ�K�PJ0�y/�@��	Nc>�ā�ɾ�c��F����^|��������q��0pw��ŝ���Gygc#�J��1 �gVQ ��-f���Jc�P�C�x&����^{��AK'�d�eĹ%�b�*-��m<��E|��#�>�#�l8�	Wj��.���'?!φz�e�X:s�l^�\�[:F���xN�рN�򼰷�نn�iHb��!S�6@]���z�D��#�
�������'b9��Jg���sy��D:� �<���{u9?�X#���� =��\Z!�ޙ�*��F��J���O����R)��լD��[�՚h5
*v��7߻y��
�j����e�~�7P��`��h�a�h×�?<:BY���22Kel|�9d%��ʿ��0���`s����7�����
r�7)?ƶ��[oLU��E8�2���x��}<��j�T@D�� �q���ݖg+�wS�ȭ�5���QJ:J`��X�fq�� I�-��"�UBl'Ŝ�|/�@O�<�s�4ZnK�DO�7�Ia{D� ��@�X��L�ZǩBr�vfAlʼ�E��&j[��'5��=/�N��HiٹExNR������.B�1r8����#�����<�h��~40����P"f��Q�j�.�r���=qժ�ʹk�+��%��ʖ�!G�c�JB�Q�����K���8qJ����t�1�>�Ӌ-��J+%	B"	��6����M����8	�<9Ӑ�ސ7r,�I�3�hP�W�I_�K疬M�� �F��O|�H�{79�|�_y6
[K�s��iu�q鱟�B��ݨA��<c�c�T�4�[.�&;ڊb�����m���'��oS�Ձ5��e�	�'�v���]�nl�ܹ._XF&.�a�!�=h�M^{V��D�t7�����R�$2e�zB֬/έى���*/'m�b��C?�Li����K��LúD�#'JG���c����ɛ�M	 �t`���<|jR�È�ӺO|ޏI	��=�	{����E�r����1��w�hMb�`�Q�x�꫶籸�O*�E�hLz���j�~��*�e�Ό4�*��M�*�D��;o���W����?ř�3��W�"Nx�z���|ce�uq<)���#G��d���ơk�'H�����ȿ��B*���O]}ϕ��bA���Ad��Ky-��������[!�\�|Y!�zd�2�p�,�⌿q�n�LX=�R�:l̷ "�9��M��-�9�����߼���q�:�1n�*�C�W1��K��=�?�)6��\8��1F��냑6Ug�q��X�a�X�]mJov��UTF�U��/�TfL�?��.��A̜�;�#p�A������٧C�O�%��(3�8˳&�# ��,-�{��9�������/�X^�0c3ie3��Nљ�4w��P!���8A��|������+��.!�����s�BZ�gm��;wqX(h��$��Rjڿ�O���8.U�x̰�*=��P<ؚ�S�@�������@�� �}���Y�p�
��=��ϑ_@�8���� ��L� �'磸���%�$O�2m�����(j���+<��~e�i�,0�S<I�i��=U���@ �H �p�g62����dyMy\�OAlL�YGS�z���'�G�8�ᶀ������p�,���������Q`_/'m�M���&�f�q��O��9XP��؏����s�qF@�T.&z�&���D_�������_�q��`�>�+�~cq�1���Q��禐(���yn�>��|A�+�9� 5�6�?~�k���������Fuo	�u���ihك���9�.��W��m��1$�lH ���2����Ej_YY���؇��,�Eb�9�:�����.��k�܉��P����q/���kP�0�h��i���J$��'ZJT	0��P�S�ב�ȒY����ۗ��bj���Kh�u���!�I�L5�Zj��)q'ד�`/����[@mOr��pf@��&:�q�%�svL�N,��*e·g����vk5���8{#�(B`��9���\D��QS�@4�}�:�'k<�zu�K~���|����]D���է��ܕ\^���r��@˃���{�W-l_ppw��_���[�[h��H͕e��Tu�/2ɬAZ�F�Ɂ�g%m��p`i���,GC��7��?��)�b�{�����Ću:���;,~�mX&�0EP��}P}٫3�mAa��Ӄ��f�S�>��U�,�#	�n?����:6�JX_�#j���#�Vh?s:���&�O�|77� j$���d�d��(���H4���YSR�"H�O�h@ζL��C��x~�">���{Y�2�n@!��Q*�圖�6/���Oýä�T��8����{�)O���Dl���;O�Ų��%W��/'.�IH(�ہ=6������&�����X3��xV��Ve.Ɇ���xДh������|��%Ĭ0����]��Qd��P,k�($�*&��,ה��+� K?�'Ҁ�QS�����_��[���W߀Ւ�WX�յ�8�����!�Ĩ^�G�(c����D���ŢfF|�G..��?��.�h4Z�_X���z� �W���?��La��w�h2�KyD��5rg�̣�D��$nm��Ǒ��SZ�t�/��y\t_��c�z�G]��`�7�ns��ȓ�v`J<���ǲ�,��Ѡ!���v��T=�#�:�����)��1w�dj��L�|3?�=7ZI�� �<��A��=�&�HI��$�H#%�b&X�%'ޣ���O�FTNI��o�N\�%�2>�Ds�s���������^���WI5����a�:��^S�O��{����݇�79���N? c���u��6RrL�>촬]���Cy^7.����}�vg�ŕ��u�kA��d��K�z�1�@��]l�F)�DG���H"�6�H�$�Is�Pm8Cj�Ӱ��餭8�dĔӬ���� WR�'@���-c6��F��� �H(�*�Q��A��G���I����]<�:F��vF~7.���T
!�"T�����#m�{x����wp�W_��t&)g�-�
�V�W��U}�����#U�bn~�M"	�����M���Cu�؆f���ў�ַ_�W��?�/�p�,r�8 ����M������2�+�W���\cR��Ć1��x�ނ���Ok���h����_�y���*V֗����t�Y)����=�G�����{�ޕ ��s]�_	�Þ ����rn����{3�ա*_�a�O�@���޿�8��/��!3�c�8Pm�������f�챀6jg��FqC��ɹK�SmHD��_9ުw�\"��o���I���9p4/{<'��>���� "�I�DDe%'>G[���e�41�2kX�7���>_Bxñ�u��a6�<pMZ���p�~���R?�t��C	��і@��B]������\�R�lW��؍���փ2�;��X�4ד��Ƀ�;� +�<���\��d�8�+��;x��-���<����Ig�Յ����02D�?�����2	*?�"�d����}
�t�>��M`�Si2�C���?��o=���|�y��Y��,���C<�gi�$E�8���l��r�n�r�k��x�0%�JD$�*�n�u��	3���N�`-���2I�� ��pW.~��5?��
]�8�"����p�`��{����yf����x�}|�;����eS�?���Y�$_H��p2F>%�<�A�E��*�(��hS�W�Q�DF��s"O�'["_�\B~�nn���W�Z�#��k��	�Wл_Gq�,�A��A��BY��L"��\����Ͼ+q�4�� O�;bPi ����"]�\�ַ��[kq���K+%�e�X_9+��-�[p��"i����:w����/i?ރ;wU(=�ϋ���VF�u�O��LƇQ j�2X��ij���Qx�i���}��*����-3� �kZ�m����B���{�;�$B�=�����ֈkN٪����F���BA����x��eŪ"%c�c� �ܷf_����Ƃr�9�>��}��^4Y7�g�i��ұyfEJ&ޣ�a"9�����T���2Srfr��D�31�?c��!2�^唍W~�)\��:�<�g�W�O��j�8�[bX��?�Iw;�A�/��ݙ����� �T� W�� ���\q<$O�5�|!�p>	��R������B����_���[��R(--#&V�b+d�l�b����E,/u$�-*U�p�3��b6�G�=C��e2ܠS�=�K{'9�����~�jQ�%�=ˮb�8|[�ʹz�ǆ.G����AC�E�����JC{^[�f]X9`Ϭ���9yQ��z�b��U~���qe,@g��*�e���(iy8n��i�8�[�]�	�1��-Lj��.�c'*]�����yD����B���_{O�����/aqu��#$����;J�]<�`!dw�4�@�����?�BI��k����~�&�
9�W@A��7o����Ւ��[��y� ��*�4{�z��r��=��`�\�c���7A�1��l߻��&���Arp�o�߀�`�~�d
���S����%,r#:��M⒕�TNѴ�0ڵ&�Gm�ɥb�eJN�J!Fۖ��Cr�$A�D�#�-UGRhJ���⤍HR@�<����pB3ꩈ������*���c�S���P��ik@X֫۬b�=V^[��P�Xla��������RK�8���ȹ!�3+�[7FcTￇ+v�����R]@�=�Z�J�c�)�p)k֛b��MXg�촰������ť4��TkU4�x��S�b�nҫ�zC�C� �&2�Il�%]5j�`�\��>f/�Zه�*����1W&i�Y��~*�J�l)�۪�HӖ ����rm�9~�2������O@��i������Ν]{.v�c�'ԚC\��l���|A=޻�ﾶ�J'�� �p.���F�	�G��e�}�f�LmZ� �Y�#g�h�D=PM�&���{�'���:�ܛ���^��:�a�$@��DQ��`(lG�zq8��G�/��f��a=آ$�ERm���l3 f鞙�{z��*�rϼ��^���nV/��.9Q�]]Y�7��}���m�l�p�Ʀ"�B�<e���2�^�������j��n���?�������?	�}���o����LZӍ=������c���M�Cӯ	w�6��<��󰩇)
�6!���
N�=`Ty���nR:PR�5OG k����j�M,c���gx��l��������S������F3q������߳��B��zf�OS�������_~��;�k�QD����<�-:���}s�yF��k5d�!���Ư�+بn �{�θ����f�s��t}���Q��I���X����h,�88<p����o�(>>8YnX�t��o��;EP[La���l#g��}�%|��|��5�����y�:!|^��� ����:z'�߾��-Tpht"!�N�Η{�EG?���$�"��&��{��(�X+B�&��fO��o�nQBe��4��=׿��V�\yɞ+\�7H2���h�g��Q�6t0��n@�}B����hb����te�e�����3�
�kC��#������x��&��1�H)0�;����ޏ�0�N�K[|��~�M�I�����,h�N3o��eTd��G*)�*�>&p�~Y�g��X[���=�J�ø��A؀�.�xXW��I�X�����,f'�N�l`b:�b�0Ʈ��|`�Rθ�����^��	.�P-/���H������Ǭ�-e�st��i�q��9s
���V�U�/boQ�h2}<%}�)�Y���_X?W�`85]�R�M����Eq�M!�K5�	��;eH5u��GY��W4�`��i�I�`�o����be����k�ikP�SU���o������/bo{��O4�8���|�6�>5�������ҹ̐����G��������x�~��{��+k�5���kw����ץ���|ֶrEλT@������_��7�4(v�wYj!r|�d�{c����+M��`S��t������T%Q�Af�d%i/�1��"��@k8O<�a�Oj�C0M�z3�xUڮ�uLk!V0ȶ�R�Ͻ:���Fg��F�w�fcUq9�G�B)Σ?���O����B�~uS�gL��ӟ�{b���G���{(4�X]# 'p��P�VPX�b��>��ML�d�"��\Vك�ˊ�ޘ~��s� ����x��WGܻױlc��yya��b��I�A�QG��a�ࣴ��x��{������S+V��vվA0� �������FYR�3ˉY���F���������@r�mܽ�
��hғS�����ϚL�]������X�.�Ӳ��Y߫�j����Ty���2�3�Z9�:�*���O�O���R��G�!LС}����vG-s������-�{�Ky�9��r3�{7B<���;�#+#���mH?&k&�*����R<(!���F������4.�)���!9�(���Ν}���J��,��t������^�_�c~�.r���J��W~	_���ޕ��"/���Sק�����9T*,"\��9��t�e�ȯ��X�	C+�5�*�p��m��o�56.]桎-
�C%�C�.��D�V�3�uy�3���E��H�I W�Q*�L*1n�q���X[4����.�}k���֓�>�C�댸�[�p���F��_ɞDDg3���m �T(���7�'��Cl߻G@�`�����-����0��@����ybWB���� �n�$no��V��>��s�'C���;x筏,;r�,����E\$�Q6�^����U��p�x�N�x���[��頜	��Dh�M�uCר,i3�L�̅	��(�ygr�.ke(�qÙ�[�r�*\\�j�s�v��z۞.z�e��6Y{�TBS�(	ġPH�6��ڰ��t3�St6��*K���P�])�z��F5K�]��>N�����d��葴3��ţ�?|�4��w�@��J��a�E�`�H�54~/��#�?�I�^<��BB�����MP�2J���������K<�(�z�T*�tJg�&����	�L�Y*�[���n��.���2?�
�����F&�����K9�4���-6�٢����ݾ�7q�iW<�n �@T��K95�Y�xhe#��P����F*�Bl��j�t���t�T1{�RV�zv�E�w��)<q�����UM��m�c��P���˗��T�����Q&hDm��r�4���ڗ����5��|��0)3�o��?� �*��G{��;����+XY_�����>�a������	_y�e\�z�k�>0���1s���k�k�����=p�<J����1�٩�_4�=q�k0��GT�u;�#��8"���O�{n�{��*����dʽ��XVK����}���p�Ek�p�b�G�쳘��P3���l��A����Mc��+���N�{�H�"�����D�L��i�����
$(3)�8���3;GS��G�\�;��d�ש����K�\��;G{|N���� ��M/��4I>��P�Sӽ�x�"��׹ӆob�3x^���P���.z�4d�	r��j܈��.o��k~p�2�^P��;`��a���lV3�4�����:B�h�N3p�F!×��ן%�����1�����`�����_��X�CIh^�{z}��5�]�Ω�{�U�!��f��(������ҵ`6��'U#/�a��;���uj9����>���IE�:1@�y�X����3�[��{w͌R�D���J�/[M8K�P,Q^���X�pf��W�o���:��r6e�%��dǖ�L�]o4��c�����}�&,��l��F�8L6��Q-��[���a��5��`�0�R�>֓�o��(I��0�\�E�b?F�`O�{x�k�z��S��C����6���p������C|��o!�-�B*7-��&���--,�@�w9�,22�ڨ��{���T���J�������}CF�jĞ�u?�!Ȫ����_���+�c��!^N�q.W�o4Ob�M��C�c�2�y8 �{x��}������~��
��^�$;�f�aTV��CY��~u�� �|�k}X��ҙ���k����ݧ�K��2r�MPŤ��\�ee�|�	�6^��[\��ݻ��<����v�1�������*�S�Ux'�������8N2uq��%Y����EO5U{���#��3����n��d�<G�#-ڌ�����ЀJ/|/�]��1�e���K�C
C+�5��O��Yԗ��p�"V���5C%�R�����47����v�=ܼ��n�5���&ץ��~�M���U	H\L�V�{�Z��szs)7��V�9�����6���%=������Ƨ�_Fee��FWO�2�t��M����\:k�A"�'.i�O,�z|��=��c䵺ǳ�����rm���L%[�*���41^:p&�9"y��!�9�ZH􈦑�*��W��z�D�L��I���w���,ed�Yi�J���~��2��1g"r�IA FMTA�YtY�J�>�쑸D��"��N��}	�q
?���`�3T���4+�;yb����9^�򗑯�g40 A���#��U���£#	#.�l�������7���0��n����Ool��G�(��]�M�fDN��7^�o���?�z?��[t�##�Ux��ȢZqxp�/l8@�_��iHf����^JM�!�i �aY&:��q=a�&sM�+�z�����ݷ~���3@c��,eYNѴ��m��@t�s(N8����2kozdC=�gQ��Ҵ�T�.����~I\c$��l��e�#��~ǒ�Ӹ���4oK5��	�cw,�w��LQ"��X�X<��IY_b��u|�r��X=�@�}��+�E?����(�h#{�Q�U��́����.�O- �q��>���k��9�y���з������X�p�6�<U�z���<&�{�v=��Z�ȷeyNO4�8�k�x�\jA���j,����5S��'� �>�H��;s~��3Ԍ�6�!�v����`�f���݉�bN�ښ�yZ׌%�"�q��'�<����a��3���F�.;)��^g�����2<�������p��z��<�k{䩷a���ܺ����g�8{���5'�RX.{��u5-dr�La�D�!�k��L���һ�ec��#��7�ɛK�<=(�����������������G7������>��8��֫�)��C�{XM�eFc4��tZ�`�#���%Ida|UӇtӪ�N�H�eqce`m������Z���hehL'6�:}��������_�����&~�r��B�g�+`��C��3��t�� G���{�9i�X_d�c�����CD~�9F��^,6�AiԻ;�<�F���p��9�oxK�6�&(�Mc5$HזMbJ�X��cn'� N;��!��>��
��8O���wa30�t�<Kk���w�i��G�pb�a=1�s��ʦ%� ��J�W.���xfs��=������#|t}�hV�FS��2<|c:.ble4��mPc��(�[�c� m�q`�Ƕ{>�1O�)��R�������3�u�MD.P$�Sof^{-&���R�#����EN��D���b����eTyOמ=i:�������-���'���-��1��#���5ܺ�� x��WM
������SC;��T������fB52'��au�D?.���i2J��|B}x�A��`4	m�R��
\E߂3�)c���AA.�՜�SR{:5�<֣�;�쥓	`��ŗ�̜2�~�8��Q�wҽJ���fk���{x�b ��$�,���>��ě7N�]%��pj�H�xH��3]��S©���w��D@�o�-�[j.`}�2ʥ4j�2m�*�re�������/���g��w�c�2B��e���"���q��_D�����.�?h[���s��I�b�Oʺ����>7���^�W6p�L/��"��!��v1��>M�GC˂V*�	�\_|�5��;1V���=t[x5����1�swvq������!@���g����,�>�K�^č�7�:�۾1 �}�;	��z��)nvw��{8�$���H29�4J��Ă��m��]��k�=�ISw*N8�I?k$ĩI#6(��
�O,{�G�Ay�����=">�/W������;Ҽ���?#L��exg?��B�~�&������5��*)K i��{3�/�McSL��l!��\�ː�����=� ?9�/����	Oc��WQ�� h�x���|�\�(F��G12�%,�%���#T�YE��h�r�k�&��ջ}d��0�I��dܺ��vg��F�ӳ��L��Yq��"�k �`��-�thS�8w�d��v%��v��y8P�(I׹��g`:��Г��2�j�XXj�����Tq��5-*�T*������8���V����M��xD+���(���Smp�Ћ�����z?�IZ+K��^YZ���9��ʵ���tn��5n�#,.�q�T�F>c�ä�"E��&2����pd��L�QL���d�M�����>��NH]т�?���z~�X�s����]�����?������K�O5Z^t����E14���e8��=��	�R< *���ֲu���[�`u��]���12��}*�it�ַw��C]R�
區���JEC��L=�N�F���h1�-&�L���`�H�cИ�,��9�F���[8I����2�y �ϛm\?��P��<��t	��/���*u��ϗ��<���z�Cv�Ő�����xb�כ�	��~F�3SNpڊn���\L]��J��;�Q�-�����퍱�>���],VV���/"�.ֶq�O��|�Q(�O�'(*Z�-3����w�̅���!V��q�6���v�p��&��1i1���6���D%9��{5��@�ix��v���+��>W�t5B匉��R�c�����f�%`P��i����}��(�D��B�Q2�9��T>+˶�$�U��p���+n�����"t.ڎ�L�	���!������]����^z�,.]XB����Wvqw7e�&)�k_���y��%ue���Bˢy��$�����Ofx#'F����\Hb��7�ф�z�N�C��X�]6�\�`QrF�2���^�IH�K�r�ʣ��+	�
%'���jk�r��t���<`S�;��-I�+8�c�e[���ףGd�{��Ws*��a&t%d�~)W4p���LK�/�N1��s���R�!��4�*ɛ�IS�̤��K@�Ѡ _o����_������<�x�C��H�S����[{��ë�6
�%ܦ�_�ǿ�g��p4p��kx�<4*ij���Y���r�Ti�\<�W_���Cښ=MT��˯�n|�}|��_G��D�n?K����`w�j���c�+�N���o�3Wq8��?����ܗx�+�u��4P%�t�Ξ<igkqe^��6__���c8PO2?�@��y�zVg��4���bʄ���[���H'*4#ț�d�5>�`h]���f���7o�s�k�92k�H�sA��S��a8Ĩ�I �ǀ���Z�q�bS͸G�~��['��U�v�6K9����-�)���%5��������%�����s5dg�2���1���+�BT]���P����O�3)l4G����G�����]�'�@��m��j��!��L��4�'���;��5���lsf�f� �׵����J���k0d0<K�3����N�W#��Ԛ&�=�GV���+�)H���@1��{0o�o�v�?/y<�F�t�����zr�=����m5���nT�tk�B��S�2#��2ϫ�|�I��O*u��[UUQ�?_H��G-���}. ')>�98�btUD��Z���h+��9�1���:N,�4<)k�"�%F������O[F4
<T�!	�,��$����2�Q�{�����Q��ɇ�_�cG:*����x��t�h�~��-ew�l b�9^MG�4Y���w�r Ey2�\�n�1O��`l��+4��.��
$F	��tO�^��*c��L[d �	θF�'�>��hFPG���������2�z��B�t|�/p�����,ξ�v�Ә�P��
S��D>_[Ev���|5'��)�c�R��Q�8���K���v0m��R��txKi'}u���IC��p�|EnI��u��ix�
-vxZG}�T	$������[Ǵ��:��g6,��w����w��Z7j��?⚌"3����&��tdj8O����c��:R=;p�_��;6���oYϘ���w���v����B���!tWk3Ê�lz4kYcF����iǗ����Ĥ���,�?	��%�]YX3��l9@���P��)ǒ���z�e�5N.�q��'���^��[��W����}`%�~w���.��=Ã{m�>��^����9������t��Jʊ��'��`����<Y�r�|i��Z��'P���M����"ȥ�������+��a���J���L;	*ߤ�2�R @�ɾJ%=8��T��r�wp~���?e��t7��d^VOv��pb��x<H�	�H)���@j7H����3�սV�c8pe�L�da}О#P���SF�o����_{9_�
AΩZ����0�����)��`(���=ϼ�
V|�W��Dg���,5�/�	�ȗ��� ��QZ@�N?3����gx-/»{Qw��8��X\�eS�I����Ơu�F�S�iN}T_�4�evg��r�<U}��w�Z�ZК/�l2_O���>�W�П�dy�&h�;{X��r-y�!N�xe�����M�	�4H��ZS�L"%�� %��	�F�3��z:��0�`4F���ɥW	>Ƽ/��o[��7ia�`�'"9�h��:$�W��P�u�J��`xH��%���d�d�D��S� �KY������Ѣ�L��TJSx.��>[{O�$��u�E��������u����D��be��2���8�&Ē�SG^�:���a�P�=�-#��L�/��������k��I��&�i'��I�X3� �ϗ��X�(˜+S*u_�m�����)����^iT[�����C��}����\�g�%cGc1W�����ç`V�DW�la�}�2w2��Ԓ������3��l��i�A=ޛr�����G� y��%�Ӭ��/tȐ��)+�X��~5i�6_{���\4.i��th����SK��QI����~dT�&˳��+i�3�Y8�xr�}���>@�>c\A�4ϑ��@��!��A�Ԍr� ���Y勝�M�b{�go�T��Pr���Ǌm���s���S�}��Y{���L�S̳`�d�!�/����n�{p����ѷ�D��e�ט�-c��o s�YEj���/]Ħ(r���#5�������G�s��#��/?�ՠ���6��>[]�o,��b��[Q	��fXg�sy�>�=č�V���Ұ�!fzL���zc�=ad���1m\.���iFX,T&h�BF�KY���޺���������8{v%q	�h��T�&@R�s<����/��5ic�d��):��
��s��x.xe�����CsD�;�ÙM����b�l ���44.5e�߿�ne��ʋ)� ��`s�3-��$�*���'����:u���#���(�76�vM{�5p@���1 �;:a���jE�>�p��}���5�/��K��5:l�ƻ\����������i��5�%��i8MR|kD1��3یo�ѷ�a��t���Y�^�����H�@����Z	$����=m݌:��皣Ւ��I����>:����L]ğ��ys��yOe��G�B��s�d�n�z/��r'�2y��(���̕�|+����th�C�l��EM�"�V���I�ʱ��c�0x �<��X���:��;W	��t���5*VxKq�ν>�\ZD�6""�̈����,Q�A�I�q����W&�Ԭ���ϝ�`Y��gPf�P�>���2��mO~��J��M�.��j︖�a�~��4���Wv�D�m��r
�S):�޻��*r?�;��:��#�2��s5�ʸE���t�Y�W�K(�3�#p�r�V��t�G
<"'K��뛭6Ln��a��@���3�Sf��kg0�+k�K-�q��ؿ�0E;!V����נ��t�BB@����i(�"�K��gW�/��;�{\��mZҗS�$��	�5�������'�mО��Ey�SD#j?���KX9���yvnf�:�E�Hm�V�Aqv����.<���e��
l�V��^�ק�4��"��<l�n�'ܿ+�Sih�36Q�x{!v�x������qрP��NN&N��
\s�Ds$i�)�I�@od�-j\�[���	iZ�U�<��P��R2(�D�L]�^?���,�����_�l���\C�h�Y�Υl��ŭ
!���z6I��6��<o���
*��� OQ��@��E�
���M���ІLyi�]�A�s�^�1�J������#s�</��-1p�"��k�o;��ŏ �|����Gx���s�N��>r�z-r2�2�k��{r��}L��l��l�N[��m.\��U��f��� ͒i�Ƿ���2Ԕ����1�ˈ(�A� >��pl)�<�"�4_wJ����>��"ڌR�B4Y��N�e�r��m��h�)ڤ��>�R��B?��˃8 X�xH����k���54+��z;t
G�	v�j��::�)�h�A��![~�$�6��)z4�C:���kS���"��	������E+G4E��W��.2Ҫ�ʕ{ع��RL��jC(��,U=��)'�D� $3���b�+(0����	2U}+��8,{�w`�;/3�*��",�_=��Z���~j�j�zj�!��׭Z����Tҁ���)�{� �^��zL�����	��é��H�ñ�\�n_�r����7���^���{{0���^~�<^}�$�>�>�;����;�mO���$�@����;�II�]YQe3�t��U~W&�ODe�y6�i�B��L-#��zyzr�ʤ��h�=�JY��:������1������<�g��Y����z��tN�{@l���eN���T�H��|���=߲��eܺu���^����d��drW���3�+��K�{�H��}�6{\'qi�#���H΋{Tӫ�i5�X���_����(�V�H�it�zO��Vʎ��O�%}�x�PCc���5�)���ޝ�x���ŉ<�o�sͼ^٦.�GGC�%�Ѧ���w����l��|S�Y�(�I�M��ZFa������/�z^k,��ԑka��m,��|���W��R����OP�\}�Bu��6��b��J&O�"�UG��<��w�PE��s�sC�U�0�4	2�h��Azaհ�$�5+з�zUN�@4��N(����e��G���}y�M�*������f˚6]A�_��!���OzX!Wz�'�cR�QYZw<a�z�����AV�/o*�륋\�E�.t��8�s�����K����m��u䖗0ٹF�O߰�������<I�=� �8<kS��S��{��ٟ�VF�mU�K8�|���x�����V�5a>c�P�i,��L�J�+Sרe���%S:�vy��ʮJ�,��ZF�/Ig���ؗ@���S�m�Ȉ	@�s���u�T�����>���ݷ֚�6��h��yo����$��
�Ο:�ӧ���T\K���S�	�6�k�h�o�;����EyJ�Y6��RU*Z�XLC�:֧c��Q���Bύ�Z_��"�_l�MV�k�	����)��@�<1)so�����\��?�����M@�َ�z�Ҟ�&vc���C2�&o�I�*o��zU����N��,�Hfi�i���is"V����晑89(s��h�������&C�4��:zt��f�sK�u� *K3e�R2�}gƌ��fKu4��d�s钭��d{,��>�X���
�����w�yjx��p�F�{��8u;�Z}F�Ҏ<��w[OFj��@��-)9�B��x�m#ǡFr�*k���s��������:����\�������,��i]<X}x��x�`a�ƟU1Y���Q���6]�I�A�#i"Dd��4�����GY�Nx3�+"� ǹeuS�6*�T�hf�ϣ��j )��°��CqN�p�aD3��ɧ����=�X&�  E�2��Z��BF�����zܓڗ[���c��~o��Ci�L�d��jڭy"���"AoƦ���]l1����V��./�$,*�k�ӱ	�{�2�����R���^o�~� 0�/���4B���"C"���GC	F�f!�f0�Kp��ZINd��@�ٙ{���S#��T�BYSQi�R=P�Y
LSV&�,��3I���W���|����؟M��>�y�91�`Თ*צ�$�s��k{L�tFі�ݣ�=O��:ߑ��z�E��T]^�3 �:��y�Ҽ�q'�w80i�T�	L�y�60���Ď�U nI<�i�����9���I��k��B�ah���B�����%\��/���K��U��Ջ��֌�����Tk���C�ō���-���l���'x�� �-/#sr{�c�=:�b��F�Rb�q��!���>��)�<s�Y�.v�;-��1�[&�?Dk��pP��t�F%��Te�!*fY��T�����Lڷ/��
T�"�ʄm<o�D:� ��L_Ɋ�7{��z�>�8����U۫�T� ��W�Vh"�ZDz�3�i;���IC�H�����);�jA���㸽�{kZd �3h����Q��1k@/M{8#ȋܜ�@IY`Q�����JeD�9�����q�����W}x�ެ�F������2p �o.���)������>>�M�����j��J��)Ӱ��W�?���
���V�F#;;�w�Ǣ�c��S�������m�C� Oݞu��[mK.���@i����v�X��s�,���I!�^}���^Ew�j��륶�����dc���~o6���Q�l�vncy�@�%F,�}�Bŀ7M���C�F#Q�&Y�]��Ɵmh�3)v���Q�i�Nx��H�{�r�2�^��_p&�o�%�>u�@I :������o��6�q`Sn&�9=+Ǖ&��I-Fϴ�ZI�oʟ��8F� �?��Ä�!�u���i7q��rO�os Q2����g`R��<�l&��;sS��iJ�Ω��2:�l	��"^�|�,E�������70�z�GS\r�Rɜ�H�u���M��Ԫqh����t���2�B�یx'�=4��6����֍{������Q#+!��pdL��P��s��$��{JC�G#���v5�ȟIb���-�|r�����\������s�c/���.��,�ʕ��p� na�aw�B�R�b�hM��j���#29�"N_��Z]e��\SF�^!e�R��s@m>���"��������S#q�~
:�(QF�q��`������,��5X̬?#e=}�	\	�N�!�xF%�511�� �i��^��Dh��>1qȨ{@C[Ԩ��vr	��,��F�|�;7�S{�q��#��Y���ب� �v�z�L�X���8�A�Q}F36����m0n��>�jM8��e�8����~d������1�>�5ާ��/t�	q��+���N�Z����f�{�c���c�6�������M�����i��=�IO�2��+�	��2�s�'+��~�ϼ�B6m83&�n�2N�(�ӱ�b�bW�8��Nsi����9ʩ)��C%��q���*���ܐ{+k�Ⱦ�rg�k��3�M=�J�mim��Ϳ .^���^��� �N����_�"^g�u�_�Kd�m�/q?etf�&�x��[�� �X�c�����ke0Ò@��;Vy9�1P,�����	��:�a��!�}�'�H��=0i`�֡�2�0�evS�����e?twhM�,��o��j���{�@sf�S��܊��]�xU�j�k�Lh�J�j��J��� *LC��1xv܌��{*��,�Z�&�'"ҵ��?��}�o��X��M,����e?a�D�D� ��<�{8s\�̈c��IT>�q
?b�{��5���<'+���h��[�������b�v��5X��
���
��Fg1}�o����*ƃ]�'}fh.�]�,�lW`:�3�V�)7��	g�������2i��WϣM�����8�5�]?r�KKKV�m��O��OzXf?�dy����X�UdE�N�]ō�1�9��x��L��ri���hn"g�}F�$�M��g��B�qL���S���K��uFS+�L
�	���_��2�sهY01i��R�J�O�4FاQ.�P��>��<�������=�����\��8��ٟ��֎M0fp��9�
��)��u����&-]�μ��/iJ�i�� ��E���Pf�*~:��Sd��z�yB��gQ]�$W-���t��F��R�4"�aUB���bo<�E���k�.�W�� �z��Uy	:�ޘN,#�6FW37&*�.�ҥ����^/7Q�!�]<�˗1ȥ�=�!�^�� �vK>��=����D�B�bT~�MK���oR�vaj7Z�~B�1�f��p�hkwgk>�	��`ws�����յ,�/P8Q�s�������+wq��?�8j�p��C���b��j�Z�l��Z�>��kn�1��X:e���cĮgS�p@�ζ�$ȿ�B��̸Ѡ˙ڟ������I�;0�5�L%р�>+�$�L���է��6�S��'��	����;���,���߆��Id5|��xMԫ",%h>8���S��l��E��vqОل�q�)�t|"�HD�j��gT_i���^Λ$^<����z�b:�HgC�Y�r�.�}89��2�1?[ڜ��������4o�ځH�e�2��$'��Ӯw1f� �L:4��l��kO���\��X�X�Mr��u�Ց�c��[B�������j���&�Ģ/�7`���o�D�2���2u.�������+��B����E�X�v����]�a�5�j��m�*�)�����㙓���eE�V8eY�˶VS��?�²����������Ɨ~�W��ݿ�:j��@�ll�+(%R��,cg@J1F{���3(�N���Zը�F�*�5�"-�m8����j�|�6��jm��*��~����=��x�Z�j�j�*����c~u�'�-;SIy�>قi<O��QMaG��i� �&2y��z#3<�#�
����0U���a7�#I�j�6=F)O?��f�� gH��b���4�@�)����VȑՍФ*���=z��L�����OV@��K�Oy�I��-�����Uh�9��8ԠR� K-C5LR�x��>���v�����8���Gא����2�����������7ʂV���+�0�M��|����XW��#�K���OE:�B� ����R`܍�Ϟ2�i�@PV*Y~�ZY�6� y[ ����'{��d<��z�Si��(�xj� r�伟���iz.�7���Ly���x��=[+i(+�D���fg��Y U)W�:N���ϝ�g_ze�h�\or�=E��HBSf�3Y1�/b"�𠨯�O�3�ɰ`j�i��CT��&�eX��6�i����ׄ�����/��K����D/�n�4�߿�1~�����U;/�GV y�4T��N��l�q���l�j�\��3����*J��:ǞʤLsP OĲ֋�H��>�iM��U�$�g��M�����J%~��/*FY���-򻗺j|kҵ�P9v\(�R���G��뫏,����T�ت(�ҧQ(w<���v4Bw��#O4��Eo��`� �(tZ����T>m�.����#�j�HV$�'�`��m\�֙��Y� KC����h\>���e���q�!j��)���5bT�W���i�+Y4�j���ܼ����]#d���N��l����`��R��7�}�S[T�R2*M�Y�5�j�	��ROdʕ{���2g�u}��^@N��r�2W�W-c�3ɏT�6	&q��`d��&�9mE����[��(�Χ���A�xn�F͵<���E�#{� �����h����G����pm=v8�\fj�H�Irh0��9ub�Μ���jՆ���]����mm�����,M�QIVI c:%8��Z��|��� �=[,��g� �J�قgY���ASytFQ�rd�*?:����>�R�`�;�~�{��(��M��q���Q2�3r��˾��&NV)0�8��A��j��鐎���s��	�q=�)��3����W�*�=�6��_��+8{�4R|��߹������e���*r��^0"�r/�M�:��?L�bb��My���`��z����>�Z�h��;��G���~���d��o};G�xf}�g�`�l�:mg#�+��9��C��^i�aޮ�u�ԗ�����������x��
�湸�uQ�΍�È��c,�i1p,8�-��M~�<������W���|�h�ة����^5�(y�J���5J���x6`��+�_H�L� 0���s2�;˳�mq���NWX���sE��ܾ^�}�(@�̶�� �L�*F�{V+��2��&�J�R�Oڒ(�.D����9G�;
x6K�f��w����5'�!�\Ǵw�6?������/��g;y<|��&�m%t�S���9<{�"���c��k��E�E~��!m�Y�l�:��*/6	8��:h�Sh���OC�LڔXf���BJ�e��Ʊ�~�՛���1?��1�=��3_��&�����Y*�;�I[;��Ӥ����Ћ��JX�\�N�e�YOC����}	�'��C�h�ɥ�z}� ��y�;u"	���_�� ��9��F��S�>\ct3 ��_Z��f��<]���z6ݷ��"�Q=�����^�n� ����qz�J'<����9��-?�2�C�s�O��O�?JHVU��?a��ɠ��� ��2�4�:̒fy������?��[�t�5���-�%����Z}��������6��
\�s�
�-/cr�� 2^��|�N}p���1h5:�*�e�����͖�SV��E� ���'�='��C- ��O��P7����2�k�"�Z�A����SX\��ޫ/����b�yʁ�Pe���EV����q=Sې��N�	i_Ν�!�����ǒ�/�t���D�C��*��=4D�KC%�eBC/0�hD���J���x��zfTn��z4�U�_ZB�������	.<��Ã{�N >��t��	���*�]���'+X>S��;��G8��cw��� ����ᴽS<��;rӮ9r�1#c���cn�Sɾ����w�'Ұ��	���C�~��VN��ZB��a�`�2G�)o�X����)��G��R�v��%�@T�.I�ZF���X��NEv�T�ٻ���=�~���^��зV�>��z�|���ȓ�^h}!.�V �����}�G�p�4V�ϦA�.�˔��= �c"�YQ2yr�.,T��g=G���跆��2=~��qǥS�� "_�Y���#��T"3$'`*�m%�$#���\�H}����z܏�l��"L3�{���Vl�GF\�RvJo�w��{��8E���Z�9�|����=�]9�.�(}�۫��e�����S" ޼�i��8U���>�!���~�.f~g�Md	Ćt����7��O�dfC?:k6�"�:�鼁��Ħ��`#���>Ϲ7j��d���~���B'3���R��{�;��e����yFR{�4?7N� �'��p ��);ԧ=��q��K�	���=��Eڗ�`���d�^��p�����km�1k�̽Ϡb��V�8��f��l�t4�3%�WM�OE'�l�xj�#c W�B���	ԥMn1eٱx������������]���z6\���C�M~�\�Iѩmf�8�ejc>���\���q�h&[N�IjM`ԌD��IJˮǳ�4�*� �i���+S9�����]��u|��]���q����<�'�h�q�~�&��)3ȧ�(���E��\ĳ>$���yD3�N�vi�`� ��P'��/�	��<��T�aP��VDlqH��R:�3�^��i���P�"�Y����3(Q�;��7��:�d/>�K�������'0w<Mx�8>�$2��_P����m��}�t������c`=�]���4v�0 �:�$8�bŤ3�������1��"�h�abmFÑS(/��v��ZJ�Q�X�����;}����C:8�	C8]W�8~D.�� �|��f�2[=^Ѐ���퇛XZo�(�Ht�������&�~x��?�������p	��	�������i���r\6��}zug\و�uju��/��?��Y��i�������$�Y:�V2r�SpM>j��A�A�TNq� %�F0W�!M��d4^V��VjU���-q+%�VV�2��Z݁#�I��6��F"���6K$韥*j�֑�������D�߶I���B��`Z��[X�޺j�������5@>̘�zĕ�U�%�K9�y������E^!3L8:���|�L��;�./2�XfP�b �#E Y�9�)!����;��A�JQY9���z���4�d���3څ�{��z��>���(��.���O�R6�HWsX��I��`�q��a����]uz�>�F;t$Q�艮y��R��IG"3+��{i�����L�VƱik�YkT�~��T�.e%��>o�l���\f.'��b9o���X��L��]�S$�2� �tT�)Ct��������h�v�A�1Z��e:�'��۟-C,g�f��w��o6��z�ӡ����%��:��x�3���1��$���*�2�����b��p<wH�B��b��1��3��b4�ɕ�c��Fe��8��ؽ�&r4Y��	s�EMS*�	�s�����`����O*�5`��w�LT͋M=W�/�S���6&�>��LF���Y�uϦ.�����h4�kV	F�G�QU`�vrl�f#�������`M��KU:A�û������?�w�޷���H�mÎ9e���T�c��M6�g������ݰ��K� Շ>�Op��K���wnb��X�g8P� ��4Qq�-r�Ԕ+W:�]M���z_'i�~
�U��F)�s�w���u��B.c��A�e�<i8�7d��`l�@1 �,�m��<:�(�@��I������<ý7pՂ��T_Tִ�5߁�(Y�9eU�ز���<#l���y�Jg�$��$�,Ǝ*L ���d�#J�L4���?	F�}��h����0X�f������\��q
%���m����*��8>��&���ʹ"
���������k���t��*���pNpvc��k	�ܚ�l!W���r�����1<'�JG�Z� [��W�h4�X�+�S�q��\���ֳ����3��[�����x���߭��g�Td�L��dROu�=����|�X���������M�+���0�e���G=��6�gi[�6�!nٛ}��������ǐ�0�m����U)$p�38�>K(��~2�v[�Ԭ�s/}��S4Av��ȑT����y��_��������r��me^Χ�;�خ-h�H������������w?R?@���ݷq���}ꬑ���n�(A�.����X�S_��ϣ�E��|ȍ�u��i��`q��*ZL=�i�E_�3��y�����/�8�q��C�A�[y0F��Q/50e4�K��fk�2SH�1��!L�@OQ8H�D&�����Њ�6���^=:Q����:9N���������"�t�ê����cNgrz������]�	(Ճ�FY�4�D��u�i`g�1��Qi�UT�R俽�!�����g/����[��h��.S����rg��d$=m]:�Z�~o`�mqW���F�����.���>}p{�&�U�`�H�_G���Ĩ�F'�FǴQ��Clױ�`�m��N�*@���ctX���ԃ*rJ���`�h��wj�/n����(��.�'�+-v��1�g̹*�ZZ�^��{&���h�W���XB��Lp��j�lF��?+��i���ԣ!���툠E2S���A�Q�Vk�3����� ����7�����;�����v��+�Kh��g�)Ns�-
�U�Xf����K/�j$���G<^�UZ{V%T�@җޜ�&��l:ul@�>�o��d�2jz�� �&Ac׫h��|S{����!���Y:.�*��]�XrΒ�u(n�A�z]��U��2|�d"��ʒ��~C�s�J�<�s&P:��v��������l�NbN2i�w�ﾋn�ʫ�!y��G�}��6*��?-���?�+���A������8"�l�a�JX<tb'MW��Mt�h�+�����x,�:g���y�6���Ǜ�����N�|<f^���əH�=K~��u���o��b&y��^��M��U�/0�Sp!0��Ɛ�{{����}����/�Cܻ~��Gܟ����6����6j�\�N02*��IOU��h��g��� ]�$�?��k�}FP�9=S�O�nb�G�~h71�L$�φ)�ڐJ�I�ٲ�	��Ɍ�v��������"{�g��&�@��pm����0}O;8��;-��6���^���̢׽�8�&��k�D�u��rK�_ H{����1n�Ĺ�J�M�Ţe�Ǉ�X��Q�pcp�x�����M��j�bmj���DL�.R}y��x�����)���}�_�V� �����-��ɢ%V��	��I���w���c^I���3�$"�U�$ֶ3K7������'�{��ֻ���苨UX��{�q	���hﲱ�؏y��7#�Xh�㳯����cfCS���1�皎��Ydb��iTJg�헌XT��岢�2�E��Y��A_��-|��v[|c�VT�����@�-������uxSG�`Q�q�VO��]�=�0�P������_�>�޸�յ:Ԏ��|FwS�&{��C7�(L��K��+��>&��Q�T3ꐑ�D"/\���+��$��8����r�B��H����W?�4yq�L�Vb�X���B�xx����Ʋ!aв�b�Nk��[����X�2X^]�>:�����F��V�0%)�(Sb��|�םS�!\���c�������}�O�x�+%��:ix"��+��|��e8t�	�� Gc�Ҵ�_���'��PP���r�v��	Jy��[�s'�_~��-�Q��|�pG�16Z�XX�>=*c�X@��\/"�XCy!���\\F���=���7�ћ�qΈχ6�L�ʫ�@TC����pC1�ʓ�#��i�ȷ\��Ȏ�'�e��5%% �1E��}��5�\�V�(U��������9ǁeu|)|w;Hp����y�b�<��!A�8�V?���ctl�h�E���!±��		�y��ِ�Α�,��6,}�N]8K㳄��84)���F>鐔usm��A���ɳ�������/�e�F��� PrA����#Wu5�q{f���t�M"I�?��Fd��X��E,Tj�Բ���ii����F4�����9���C��K�VC��]���k�˄$ˢk�\�۩�'זN �����isG>o��4qZB�3�����̳H��y5bt���F0	]Ka*	�����^��ԛMi��9�������J���e�y�s�&��Uh(���-�.�^?�ʵ�b�+𑚇�߇��<����bB��RI���M��~����E�b��N�,���_whDqG���q��:nݺC�D��  n[�fƯp_�,g9���ǀ����� z�c�FEfҒV>�1�G~+���D����������^P���`���T�sN�-۠��w-*�ޚ|՜�R�<������r���#z�E�;3j���3�:�2yR^B��H���aT�A���no��������l�hť
����!0~�ճ8�z�4�������}�{�$*�s�F0� t6��h0���2���"�1n���`ss�@qc�k���� "?*���rܣ}���-�q��*��>�.㵗.!����=����eSۊE����~� o��s���9�*k�d)X�M$���ܟy�Y?�7߿��~�]�{�##�O���m�>er��y	��e�Z�b������s�룑���K�qf}��z�O�o�ә�e)ca���IL�:�ۨLţt
7>��?~�����+7�M�h.��;�%�[4�y��
���w��;�O�.-�3��c��|.o ����D������&-�L�ԫ��i^qm�	�k�����wߧ��0M���Ѥ�Ģ�g3�ofN��z��t�R�D���?gt�u�@���"EeDg���a�F{ߟa_�/WB͛X��F�Q,d��ˀV�t�ݑ�w&)995E�|En�b�l��H=+��u�
3��h�aRY��(���;���Ό�tH㒧�^^Z�1mm^eI�*����hJ5��u%�6ﱢ�"���ʵ8hb���R��0��U��!SJ� v9é2��Cr�<5H4|9
y(��Ȉdh�fi:����	.���G�r� �͕z%�qɑݺqG;uL6VЯ��ZG��/2����g���z��4JgsJ��i�"+�yO���*	o��!##:K
&�d�����zGRżت�j��ͧx��yX����sN�Lea�u	T(��Қ.����!<���t8F��.���a���k6�p�g���>
��2Rp��㩑���\[0CZ?����w�PiM�Ne�Z���?P�{r��ٛ�i�ml��e��R�~�̠��N ���'��g�a)+a�ʛ��>R�p�0��s��@,!���va���:
�9�c�P����kZ҈Y��ܑ+�{����:7���po?�?f����Oh�
?N��#�����A"���	keT*���s7<�G��@��u~����-;�+�������o� T!�	P��n�������{���~p�i�{HC�d�h�ԤD�	$A�P��B����9����}�" Bj�`n:a��[k���d��� �)�ߔW�~�@�}��X��R��63>f�e|�?�\�\L����
��pFN]N������g�Rݔ������E�S_�k\ͨ���յ)V���Pțf#t����S[�h0�'� �� �c&��m��|>�D�!E� ah����exh1���c��8S��Ų4;q�3ڝ�JM�w�#��;�ܧn_N���}%m���q�}��4)���)vR��,�ͦ��bp�#�t��3xf������|����"0ru�,�\��]��Ȉ�"#F�L����!�1j*3�<������[=�����ҝ�-��S���& W�o߬˭�#�]y�TJ6�!���{�e��|�w�?+�h(�]��Α��BZ�AC�IK�æ��$)	kk����S����sw��{ �A$����9�S�7��ue�`��~N�c_>� ���޾�um*{�9�@_����ߗ��Km��i��Ï�pI����
T�^8��>�<R+rν_��~׼�{�$L@���_���s�5�pB� �:����u���7��9Н=���D,�?�M�F�:��	�74;�9u5��g_~꒼���R*���sm.?>��>��Q&��ް��5t���ݡ��ڑ�wD^k&��M)V����uH���pfC9��~���E����we��1u�Ne��?�����h<~�D�Ʃ������)�Ƈw�������|��d���F���7�7ܧH�O�=�P\P�d![�~�ә�l��{j���A�W�4�D\�#�F��8?2��ҳ_�SgN˹Q]� �x1$�4b�_ɥ�ϒ-*H��I_JUu�����0�����?��W�6V��.��\ 2f�ɀ�@d�@��xi�M1}�,V�ή&d2�u��F�
:���!���؉�C�.�O�
bx��;�>8��l�R7�$;MC�1��ѰͿ���`;Oe2��!0�H���2z�A�.ǭ�t\�=]�l�,iu��VW�1���GE�W��ʡ~u�wi�E˵"7':�r����
��2	[.��F#���:(4&��LLhKqD7�cB��i�� �9��5@'�l`��ф��)K ��}c~�Q�r�K����k�@�?�"����Ce�����?�0 d�#�+����8X8���|QJjTP����ӆ)���p��d�)��"#��.�k	s,��!SK��τL�Y�9 �y��w\ۨ�{
Y`��ёt�ko36��U��� b�;�#H�/��k  ��IDAT��� �����3=�
�'���V<���-1k�Y��r�,2��Wr��5:gÔC;aK+�������.`�c�3�h���ddV̽��',G����xw_r
`�N�W�蓓;qf�P����'�G������V�&Rr�iP���>l�����Ҫ�+�J���y�;c{��f��8�� ��-2z�Z�C}��$c��!8��`uaE&��Î�d��$?�����Qh� �~��_����<E29lJ� @���t�|:��&��iǴ��ьt��,0�%2	Sp��x;�C[u��tqf��?�����b��8��F�e[� w��7hh��?�/�Am*iK��6,�,�\�f3Ϸ�k�e]4�����W����q�d� ���dky�ץ4I?��Q >�+x���hg$���reV��oO�=3��iJ����g�~Nv�g���6VsH�˼ݐZ!�F�7?��J-cİ�u�+(��i�4��@�q��V�A]��W��J�ɻ=���r(o�7�O�V_�i�Y+�:Jș�=9�:F��;ץ;�s��s��yy���-�i63>��ޥ/L&�Ě��l.��;:��Ԧ��I[���o1�7�u� �2e��ev�O��XAe4_ ��[ܫ[U���"WNo�n�O?�Ǯ�g��b6�,d�;�yP�~x�����r�����-�'�*�?P��gto�Q��(������1��?�)����y�����B�K��_XB�H������ǉ��W|;�x�9(,#u^��������R
h����1�^��P(e�`f�j���{k�;�����r2/�hD����7B��'5�j��Z�H�"���hJ.�veU~���ȥ��8#���b���#5�]����f!!�fV�H0�e�E44�>��:�J.�(�ׅYZu��?���5̈₱����83��~�ʘ��"UB��8�����+��#���!�-�qO��`��0!Yo;o ����W|3����r�k���*�?pr�GqӾ�<Ȋ�d)\��c�B����Nܪt�܎�]i���s��^U���kjd��f�#�VA�J)�]9L�$�yy-2�L3�1˨i��"�$C{��dK>;�h᰼��,��t��L(Oo23�wa�A�Ո\Dt�,�0�nʒ�@���0�#���+���|�@#��@A��S����赙�^O���`��đ�y��0	;kz���H�쏆^'tE��<d��{Ŭ&O�S���rT���=R�l�BU~�G�n^��_�Dn%f8P#���c�K�
��9�o�Y�D���V�=�Y��/&���	y�þ����4��zN�@�<+̉���4���9�%;�����i��8�v80."�����P��dX� �S���~~8	8�9�r8sg�k�� ������xN߳�@ϗ����o�5Sw	gpML�yJ�z�3���ٞ� ���D2��X����că���9�4h����Q� ���5��d��ץ���k5�M#Ľ{���v�e[��:h	�D��Fv�?��=��ă���!�Eh�3�s�8�f$���'$^ZjWIE�@��h�����P�#Dc	&�D(�(������G�����/��(�I&�y�s2���f�(]�����P~�$Im��d/M��1���m�︴k�~��&h�ڽȢ�OL@���lL���J�6vB�o�fR9[��x�{w�$��ʨ�0������F)�`�3���rC���O�j�a-@+X�� �YS��+h�������f
rasSm��F�4�h44c��2qdk �� �<��n'帑�@�&�ޙ��G���8����,�Ҹ;�����͑��o��5�������c��-@Z=����?��F�=�5��'qC�� �uX(���7A�1I�XYT׏b�;]���D^{�]鵏(�CnA�� dG�*���I`�H�W�NG��_������{5׀����.��O��&nֺ��*�3�Mt���>�_*���+r��%��Ҭ糖��bǸ"�M?�V�҈n2���j��������{nh�x�WR��,݆���x�/l�t\�c_�C�|ǱJ���8��VO��������\ACO��2;@�7�[#*d$�(m�Q����c�Ц�T�=�%���L���y)�c�;C��1z'��eZ\;'�0[M��/���|�Џ_����KyƸS���x<�&t���R�8�|J]0)�[e{N�@9D�$aJ�zQ�����O�	�ϧ�n�V�	�m�]ypX�)1��QN���n�p��b�P�Q�]2��"�s�B�VLv:�{9���D=��A�Dz�ꑝZm��8g�ƈ� dRi��c�%#xD��"A��;���sU�|jU
���P��H�a�p y$Ӽ@

�r������j�
I#�RN��è"'k�����X��!�AB<�G���
i��44��!�2)���̈́��C��������2��Agl�,���:���!�I�Y�B^�9G2E$����f�B�t�Y�dj�H,`X�������(�����Y��1��i R��pwO��|����I�b�%;:�=�~\��c��^���uc�P���@ω>���'� "4���Bj�ݛ�����p���&ʖ�����N�#	�pD�\�1�=��6�M#�fv�ރ��`��3�������}�Vv���@�2yz,�r�%�$\� d�v�R�7�\*1�����QD)@|;t���U�F�͐��G�������J�����bM�ךt���GWG3��ΓF�T\�ߕ��)S�\a��������;�{4�{�c��0���$���-�<�{8��Xr�T`���ަ|?\o��\��.Y6g��a�s ���;u衕cf�5#��a��4�)�<i�F�b�mC T����9��g��vu�,�LE6# 8�[�}7\4x��Q�`�*�� 1�}b�<A^H�A6�ylP�L -���r��Ɯ�����\�}�����X_�l`F���:3�&���&����n��W������{j�U鶚�AY��( [��?A��0A�z��`&��\8uF6W6���s^�{(����Kd1J�%Ӗ�o�k�����|tБ�.�OOZ�Ҟ���V�ԅM�G{�j;B�7_�6�VkE�ݒ�ڒɷ��OVW�4����!�'��fj����/�d_a�7��>��o�Ͳb�g�V�-������&���8՛q�����/ߓ���5~T����A[��o�G��Yy�Z^=�f��aS��S�jo �̥s��m���m�{ ���xҌ���q1dq��)FL9�����U�,���*�_y������T+�6�������+vW��'���5b�Jw���>����/9t����%��祈�Gԓ?3� y�����B�Ԭ�/���q�c�ɱ�S�el�Vң�d�QH�M"�����?���[o�N	$p[��Y��|u�i3�H�{��yYY�Ƞ۔�=5�})zsZ�d�Wc�JbU^���:<b6!�;-��ß.(�RSmQ1m� &j �����'�`W6vɺ�����1ϡ���3�J)�Ũ��3:B�zNJMy%�׳Q#xp$E=7�S���f�I��1�+�<ʃ��m"�d�4���Z]�鱛�:�{;!���hڀ��=&�bC#��'"~?�Rx& ��lVƌ^�
b"r;��T��lq�$
P ��1g�:ì��P��q���ր�L�\�y�:�ʄ灌,�r<֍���=�볌�f�D�+�r��m��4�<h*��bB ��Dy�����u��(�!#g�M�=���mQ\�����q��rjS# �9.��sȼ��qI YO����'�6Yop��Pv�k���)f����`6+�t	*0{��Y2�p � +����o3S��W �"���u}��gd�J�є��u��N8Gӡ�	DPq��MPc~ �H�98uUH��gl�
8��t�� �x �0>m��6��h);B�R$T���(E#���)�;���]�j�T'D	?�~A����2Q_�V�~�p��Bg4�Q��kY��Ԏ��m��ٗ���'�pst�D��A�Q�ɲ{G߇`�5�t�2+��<ĺ��{�ŬK�9��(+�Ƞc�Nb*٢+�|�H6Q̾�NXp���� e�AM�Қ�OI3�<f�5�t�^#(ѵNl���Ӻn��gdm�w%��B����(x��/�Ze����E�k��29�z�z���՚�߁���1`2������6������7苨S/�m�zK�=`�*�狒x�M]#])�sEu�;�ǜ��^��2� \L���6��2�3\"����#�S����	'�8�!��Κ�(�����ց=̈́��g�>PRP�w{FI1��ݦ��̶�piNh(�cKP�8�q-7ٱ�����A�fܹ�[4��r
���?��x��/���B��~�u����L��ӫ��&������T���}V�}_���ퟮ�ՏUdk������r��D
F�;{rw�5&E�����L����{rOA�@?#P�R]�Rޫ�1���ki�0�8����@޻ޒ��NMj�S�g�ߓ�?x[~�;�rj×�RG.l?%�.�i/(Mc�5���,5���C���u4����EvuY��ΎtdK�b��2�&ު��H�%O��Վ�98�?���ț�_�<
�+]=7H�a��QI�S��AoP�@B���g�l<�!���s���c���]I<�MӀ�$n����c�:E����t��o?�����ҝO޾[�vN&XL
.R�BG���LM����G�	�o��<{����֗�n��^��^9/g�y�t�'�G��,�<�<�iV�Ll����w�b����O{����������
(�ِ#f�����G	�kC��h�� �h4�P0����:˳S]v�c����F�6�"�Cnt�8�ֱ�"��dG9�5E5�9�� ,����S<2=��g�/���� {j��!�XZv��7�Ć:tG���?=��I#@��l �hz<u����K�%])�
)7�(h�u4���=�$̸��;_6zYh��d�����%��0�P��4�Ȃ�������yiKa�qC���2M����*���L���R�1*Gt�S��3�ω1v�gJ2�����䴀8M�����z�3ѵ�<���1q����vz���rw-0r;�J�u? �6�2J0C�L(�$��!KgbS3��Ǭ[|8�<��؍ju�|��t��T��`$����^h+ A` �R�D�5&es����m�QJ��uý�w�i�t��
:��}����*8Od����5���ng@��} #���.9�Ls�QE�	N�������$�c�S�ȝ @��g������n�	�������eԑ:p[q�p�C�l3	 M �S�wB�Y��)��k�@�q���pt�j� `q\��i"BF �Q��"�� �Z��+ *E�HCB!���g�f�5И�`D�i���6	�Z�o�&��u]'3�\L��IZA	�"/2YZd�\KІ�RS�ó�|Y&(=��.BcR�6 �VC�ш3Ф��`�ҵ����M3벫�'W(JC�s�����ɭ�I�롫���,��ިM�#CW��Pm��
i ������S�H���CF�H2/�>���U��W1Y�V
�shi>
@z��stj�$�Z�2��a]�
.Ƴ�n�X�Idr���������HL�@��@d��d#F@p�qlhܢ�
�-P9pft�X���>ˉLƑS2�?�=��*H�-a��" �䤡g9�aֱ�?
U�i�
���k0bs��#��uJv:�� 5�fD����g�9e�P?4b9�w�� :�:�i]�����ޡ��q�,6�d��I_���Q�d����\�xV�j��rV��ǻr�ޕ���
�z̎�PMB��À�g�?���G������Yy�JB>�uW��"��-�^zJ���ߐ��{V6ky�5�E���k�g����|1�v?j��R6��3]ۏ먀��#����#����[�o�݃�-�y�#S_`�`�P=�i���A���e�}��3��dskM�v�)Yѽ5z��$v�%��<���L��a祹6�BK���aS�˺��3r�u_�����R�#r��B�C��n�d�"���$�v�d�R����ސc�s{��|��ru�Hp�ı2�j�0:�"`1�F8$��,�G<���E����3���ޠy����޻.��ߗ���T��P���<� ��F�����g/�cy��{(�F��h�F����E1�K~J�԰�6,
��7bg`¨?�V|_=�1�kƖP�}�=��f��-y��U�J_�mc� �+�׿ǉ7�>�9�ADVM�eVw}
��%�z��x�c��<#���*hz@�
YE�yFxp�x!�����`:�&��E
�V��eV�b�0_(a����L����`�S��+$,���26�a��+:��j�����c��b��.F�28c2�Q�k~<1+{��Qz*��<�:��B�R�J��j<wn���l���:z�?�2Zw�n�X߃�-KEV>&�0r@R��9��H�3#�La�l�ޤ�`t�k:4Y~r��Qh������B8Vێ�����иA`�N���S\y>6�)rv`ȇ#S޲�S�]G��~-��\/�r�Ƽ�,�R;�%*"%\3w�	)I]O���\�d
ss��Za���)F���A�<n�0��s����{a��Ԉ�zV��`�It���ͅ(u��?XCp�WFG<�gȶ����b� ��\[t�3���,�8���������rp���������#$�W�!u��ڢ��-Y^~��K�
�p0fپ���iCT���tVM�Nr���ݿ'ׯ�`4[L���j��/�=|[���m��=i�����R��٫Y�6p��p�u�=�s��k���ܹ�/?��um�Tu��
<ۏ�'@2�Fi&��)6rq������l�l�ӵ�@ֳ/)4e!��l��@�xh�W}�Ӻ��3>��/>sE�=�ڵ��|�f�v;-]���49�#�,έ�6s�1�:�fZ�ϤE����z��YY���Iyp��hNBpK�����`	��R�L�&��j���F�j���1I��ʖ-7"Y$��c�F�G�@��ޡi��8����%m���]!���z�:B9�	82�PA� Sq���LE�?gt�d6X-�xj����zg���ǒS?R�Ϥ4�˚��rw ���`����Ƌ��?}��Kݔ��[r0�ep��$�!�H��}� ��ܓ�yG^|�$�������wߕ}ە[�-Хz�����#y��?���ʥS�rz-K:�2\RE��B*G�����9�z�m�2I6@�L�c&Y��	"?@��r.��'?�vO~��m���wd�~��gH��jQN1���	B:T&INmc�M�z�g�6f>�F���o}����)���D�ێ�8�1!�ӧ�.�R��Ix�N5t�����WR(�����GO_���Q�G͞��A�c�x'"�Ѕ_�i��	���(xi:��?���uS�����K������8���f�[h����ȋGr�#��e.��b�Qg�~�x$���O�/������������#��`�HҞ��W�Z��U�`�H�6�({��]W�}i:�S�,3ݑ����:�j4Ɯ�9 �#��l�E��y������y*��:��u�:Uv,!+@R&af��}0C .W)�� �#)D���
اÉ��͸��j6�ql�q�D]�p6HSzn�����ມ&K���h�V D��
��s�B$�90�r��<��dJg	@�@�'��2��;�vԜ�p8�k�P<�����
��� K(�yz=�=�;��:D����$�p<1��/8r��q/3���w����e4'Δр�dyA����љ�Q�+�����=��|�0]�R�k�A	HpD�]�̌��g��k�=��$�&"��-��ی5'9X>����3��������-���g�Y	
9r��	�@(4_��Rg;ì��X�Gu��_��4Zu9{��l�=g@&{�b��yH ��=�B/M�E2��!����N���P���Q3M&��1"`�72-x :�k�XC��L�-1�5�l�m<#{��k��Y4}�p�0N�i��9�̖�fC��l�E�����N��dƒ�=�����]^��J����r&�'�~7܈X�@	%d�L"�T ����sn��l�XC�\B��o��C9�{$+(k�����ўk�Zm=g����Rzx�� l$�n���w�U�R�2�E���Lsz>�ؿ�5ݷs���/5�I[W�z��|ɑ�Y%z��-2� <������MJ�q�$x�(�!�����C]g�~�{>���󯮬q���vo�f�\�rBG;�r��u�{:�B@ļb5Ǩ��!B���<;Ron�z<�:�!;��r��9�x�ܽ{W����~hL�x&�)��kg�g���>	+r�B�;e tKQU0n�W4�Z\��'Β"�Nu�`�T�tc�K�BMG�e)B�l���e`q?���_I;� Mw�<Xc۰��&|p6��R6k�i��je���kc=�����R֠���@8���ǼV�H��'����ڂ�l�����s��z�:pF�F�]�ӈ|r�i�������������gd������Fe����e����H�5���K��׾tQ.�ݐZ>M�-5���<[��X�-�ױjG���+�(��6�g$���^_�^��ƍ���7�ɻ�?Q�����͸�99�� �Z��.�����õG����{/\�o��R��+�7��
�]·#	�~6&z��s�h����^��w�j����<��ߑ���/��P�;���EV���,(�#�:F�F^F-<-Q��N�(ܓ��¬�����5b~��#����3g6䥧�*����HM����aT����\�_�h�X-)i;�!?��!��r���AO��oȏ~���;��@�R�@f�=4	!y��
>D�-�K�?42
��{
y���j43�+aJ�j콁�dZ��r��o`o����`f�:J�E����n����J���H7�^���g����%^{ ^�!'���Y�hqjD���@7�P�v���a`���uS2@�P�`\jD�\=�����
R�9��xdƐI8�*�d2`�����	(3��?��s�(���=��h�k`8hw���A�Ѕu��|�>����I�e�B�44��|�
Np2��Y�qGT`��f�m.�a��5pJ�ᜰ~p.	^��y"aGEFs�q�*� r��%n#r� Dv�3��`���ؠ:t�r-c�&
�C��g���L4��� z����q�| 1N+��,���,2OQ��e,+kU)�?�42�rr�����`� h�s����wU�j�A�#L��R���L� :�)^�k	���� �luXZ��J�F\t��c��Ie,�3��4E��!0+�{��)pl�����%
�>�_C�k�ɘ�w4�^��:�� �ԝ���aH��rlSA1J�x����/C�xԠ'���ù��u:]f� t�jYƝ��Lp��} ��s���N��2.�g���; �Z������������4�XM\�c`�?��)�&�+�M%{ؗ�\I��7�q�CO���<�j�#t�}k�&�@t��t��1dRH�u�{�a�өgG$�@�3fvq@��D���fY҄�ɠۗ�;�֤M�����N�YNO0��������ѳ[���k����N���u7420}\����g���b���Y��Q��1�?4�`o�ӉLtGz�I9��cH�k�Hg]C�4e�as�ig��u�-�>�b-�TG����{�9b�����A����lY�v�R��$��S&
F5D����W�zM ����(�G���1���.y3�~�FP�'��R{7�u��`�R'v��{�h��{ґj>#��%��.JU�Ov��+j]&o$�ꁜ]]�V)˺����}x�B�]�2���&��,]'�d*��5�qבk������֪|�ٴ��Gr��{�֛�R^yY��Mz�o���:�X~~�\<�-_�zY.lk��-9(b!����I��j��6�ǎ��!7b�����O�g�J�!M�]7w�r_��=.n��X�t��%T�f&�Gg;�3�6�RS���NF�0�8��Q��x�'{���X��s�����g��$�~$�GG��<��h�|~�ӢX�o��ݞ7>���-�ݳd|~C��w����sG��"E��2)��I�4�ɓ�@��c&#�K�����x(��ܕ�g���Kg��g�KW�ɩ����t����X_�r��^��}�"K��(�*����z[n�ߓ�����c�u���|�r������<Z�� \���D�~/Ac<��L"�M,�G���RP���(7->5�BtI���!�(x���帶�����.]�� Sh��rR׍��}�~s�V�5�p�$+ЄT�k��p$=50ǝ��Ӫu��������4�G(ob�4�4&�ل����m��|D"t���'�ɰ�0���#��j��2�F��3g-�'W3p~��BF�zy��r3�����,�̈�N��2����������i��/;{�	�Т��aC�6�r m%t��� �e/*�GfL;�Qr��$Ӎ��EY����3��^Q�襡��H�Lt�DV��݀�W0n���eF�a{¦f_ű��R.L�*��-�# �:�.����u�[���V�PO���_Sc�F�,�:`�I�-�����c�r-�q5����h�'�� 8��ؼП<�y�%N�%f4؈`��Hcp�3ă��T�F����0�՜˦KU��� flK��CpFN�:6t��]w���l���<��iǳ�8`��P�P���jU�^�c���>J�E��*;])��H�Q�&��J�ϳ�i��b�'ʶ���LS"a��[��b9�&3�җ))�,o��3:�쪘�q���?�#�CO���e�
�S���NV7�<�l�z�\D�3דAu*9���l&e�#�8&n4a �`��kP��Lj1�Q�0U����)�m)F�`Д[�3���O ���x�4���R*K�w��~6�f�B�{o���[M��G�G�՜3��[�6�A���e���sitF��)7�\Y���d�
P�:C#��{/�[		���f�x����L��&�;'Sy��J������.��$P�!�ro�6=�e�|ې�������G���맴�|����yV�检�hq�Y���ߜ�.�i�P�H}x�8�2�M6L�;�Q�a���P-�heM�����Kk���\�~F��)�#�'�
λ�6�=D��.��n�H��YVV�=O��G�rQ�7��&_}�)���ؔPm룽�u����{�S��r�Ѿܺ�H���#�xv[�y�=�9�R��۫lZDz/d��GXh�b$N�(�����F�`�@n��X6�����կ�u���`�D@��e���8%q4�^@-R\0��Q}H^���4�Z�'��7�N����i(��<��=֤Fq���$�>�-������Ł~�
�$t�D�(/�\Yݮ)�xJ~xT�zw���'�l��&#(�愒>�|�%����|82A�Q��k���w�[�������5y�̖<w������ɐ�փ�@�� M7�h����m] ?��q��AjFǧ;��^\ �aO> ;��x�\ɛ J� N�>�7��CBTWT~�Z�$�Ҙ���]}tg��\���(0���X�=,��%���1�0��W��{��P�����(��I)'�&���1��1��k����J�8o0t��#�#@���D�&�7��}�t�ZA��Y�>	�N�g�=a1�2�P���$�>�q�j%���Qw�z� �'P�E�-[2�kjT ���A��i��Ǭ�ll�(7����d �D��q0(�'=6J �0�����l��p� m У��Np0�S� ��;̺2��C�d�l6M�nF���Vlf���&�S�)�A��LN��k�� ��I��xƔX�U���ѢCvO�v"RC�켧�ҋ���0�7JЉ��]�v"��n���N��
]��'��No�ə��Y��������`BC�+��(�	~@��� ]� ��B�sf����=�Ǜ��R.��p���/^������\f�؍�S'f��,,��ɧ�����$t'a {<��+EcD��P���(`)�@�H�PB���sv�̲p����@��NJjxO��m^@�����5�xB�1�ZA#���y�<�v�	��RS�5���֛ �w��3I��1�)�T�	0�73WY^���	d�@@��O����B^�k�U(c]���t?�T���C������
2��f�Ҝk�;��$��|�!
0���w43�B��FQvO��j�N�)���c�	 i��kxf�Еu(v�:}09&g7�S[�c���z������if���!1�re{]��ɬ��Ukz���፛R��'1thxxK�v���|c�X���5c��욳3�#�o��q"�"RfȖ~��O�ޢ��k��	*R�M�N͂~f�H}D�w� 3A���5Pjo5�NB�e��{��� �_��t�:�B4��0����9��io�d��o<4��R9/9��U�����>�P4�#�D���6$_8%=)�&B� ��'9A���Ӗ�nOV ���{x'���X���K�Jz.��rxؑS�j[�n�*�)tÏeO�qo>c�5�둛)֐�T3y�{r�/��[����\�\����.����=��n$�t��ofW��g��l˻�J9��+�������
����'���%UK��әK�i�{�HZ����������qKM�A	i�:ph�Ca�E��$��j��o��:��]�ّ�z�wD�f��׷��?[Y�W�l�+��=�U��j��G�,(U�����L^�ę2�M�t���x �lYr�8�n�U��������'�����hUVV7e�K�՛hI
��`��FHO`|�.�HӺ�`\���������7^~Vʥ�l�7�X��mi��cn����.o��x��=i��9j�n�%o}tS�K���@R
Rz,8|QF�TJ?�r��z���@���1���[�8�����ɍ۷�ZWzz>�gݼ\n�e�ёTt#��3f��@:*u�d��3\�c�؄C�d*eZH�Dj�FٴFG.����8M�b"����>��T�u��$��.��n��LN�?\&*~+8�4(�4:�T�W�1�j�%	*0���(+�F���32Ug�R,
��^3�\��ρw�ײUo����5�A�eA� ��#��:��FE�ф�aʏp6_D���S��cI��qn��0��'�Ei����f��d�0�],?ϔ�#��6��Ap^���^���څ��>fF�|ILxȠA�g*<C8�3>�Y��j!��H�#�d�fq�	0����J d�y�1BVI�q�D�$�׮��,J�N�hD�$76�8f��vt���K��T�@�7J�$R,�@,��! M7ɌL�7����D�� N�����pgGZ���q���
�����5u4d <���V&�1�7�����8�E�� �����)�b��x1$܌r1ڔ� <�F,E���)��X'�!_�s	gC&F���A8���в 8sM�	�h dx�� P��m�Y���10�ŐDy��YPH"��pF��#�|�D`��o��̖hc�=2�C��<O  4�� � ��]�>��){��20 �1"kh$8�������T�[�AFAA����wӜ�q�i9�ϼ���\������ο��T|�-��~d��k�ϒ���5�9l��Q�x-� )S#W*�J8V=�NdttcP�׮�37#4��+��Z,����6��4���ʱ� �Ȝ�J�ʁ��iz�P����zBfٵYǜ~���%W̳a��vś�l)D�1��A	�e�LIH)((ƞB5��%eoFCr�K�X�X/)}M�~$�ŕ���Y�M.���&0��Mvnjy�8d�`�`Q�w8�v�����4�Q�Ew,(P�RV���Pkt-�s%�7=UY�����6�m�z��|���.>+{�;R�p�F�P�N�����k��e�'s����`C��f���W�SI�:��uîl���q�e\f}���gm5���}�\ےRyU2~M^��V�ɿ(ddk�)y�kY�����פPβ|>���v�5NE���	�Cr�wt����;RT�T.�u���Þ2���N�=��C�*��<�['#�y�Q���G��45��\���4�kX�TN6�֤y(�o-�qC]��ÿ!3:AbC�o=��o_>%�dkK�?h���->�	��=���Lz@�xC�g�<C@t�F�1ë�O���af���O�썏����ʷ�&E����'�wԖ�D^�H�4�_�F�>`��4U�N�\��Ϡ���#�$��IHEI�����d�Ԗ�̦�*�d�#�|EtEP�dtD���v���S�5uJ	�]_�[���a
�^���U�B�BQZ#�Td���Ad�=ӵΥ����� |�٧�@��C�ˍ�weW�v�*�/gC��jU~G�z�#�HP��S�B� lOo��7ēՉ�P�����N5�����H}]Z���͓T���z�ok$s �.ʙ���ͫ]ӿ�Y![�w%��Ӟ��> �d��V��H�"�;=<�jڑ��D*��Z����M��MX�&���,b��~& �%/}]��pG�kM�@X�9�޾���p<}�)JA�����.!Á��I�l�}G#Ad�#�
#�Қ���>ϔ� �n�f�/JE#�"���^Z˩7����х3�ۣ��9I*�� 0ΤL"*�j���)Jศ�����5��qM�$�43��:)�9����%��
�`���C=nf�ء�cJ�� 4�|FtF�q&m���7s���1Tg܇Μ$Q�ۦ��8<ϔ��>�*h�V��d�X&�4BU@���A�,�9�����"d����5<h�?fx�&��V ^����E��h6Y:��y�r<�>�$k����i ��n3��(�#sk�aM�:���S��&2P��۴�_ȫ�hфKN����MP��ed��>Q¶_�}�j� -8] ��f�HGp��K���L�v�<F���Kpt�aRJ(�gB2/���t_"�#��� 7�����a!�,��Q�;e��n[�!W&�mB�| S�ϥLv�ͻ�{C���tT�(wcĚٵ��م��a ��*I
&z�~����`_h��h�������Uж���Aʑ���s��?1M���"˯{'�Q����wh���?K@�)��C�)�2�p�p,rƷ^�֠Oٗ���>?G��(�dX0\K���zC_��2��Q#��:�����w�e��D!3��}�!��<p\k6��F�ͳ��@[(+��=FP�v��$��s�)�v��5X��Ș�-�ٷ�\���Y��l��z��!�\�Z�����k2�h�aS
���L��4��>�4�X�ph�>'����޹!�LC��_�g9�A��H�(8������{gl��k���B���Z��l�ͭ\�'К���x��/��ɺ��ߩ�ʖL��QG�5@�60U?�h闪xk5i�߾�ޱb�-y��K���}n�*�]��4V������(�╤��@�UA��t����4&c6�M�C�ěGE��D"	���������K&���:�ٜ=q��!ǅ`(l �=u괜��&����{r�s̻Q+TX��m�T�ra� ���!����ڵ�U|Q=n����&���wdhm��y'��q\&ːDd��ٟ���L_#�kw�7�~�)*��wݐk;�ȇ����:��!��*r��4d�_7Y�󂠃<�?�P0���;��AS���w��)Y�f��6���x<L� ҆ *�� D1���uw]y���흁�yT�C	��V����a`1��%�+�بn��6��֭;���W��˗�I�t[�߸+�����婕�<SJʶ�{�ݒ|���/�Z/4□3'��i$4��d��-���)F��S�#�)�W�2��Ҳ�E��a�F>��rR�΍g�#ʳ x�x��A�~R&E�23'5J.�}B���L#�P�� ;�l���|׵�/�t���^�1f�T$�u�kd����U�^��q@#� @�Qޠ��JQ�J�#�L�n�L~�u����4��sLTX����  :F:D�mL����_�B�Fd_�(��i|��A�F���L�XL�mZ�E���C灿޿���� ��He� &}���5�X��h�/��vy5\Et<�3�����$А�{'��2( [Ȝ�'�5������<d��@�����[�ے����-��I? �Y7|��fƺz��ٲ�9m@�#'
ư��n�z?P�7� �O1�W��{�{��(�<�N�	%̈́�Ŏ��X$س`��i+�u�{a;�(�c3�x>8���-�^�����Gj�0v�m�8����:��<XdV\�����?�V��Q_q�Z\,�7Ѥ�5Nfߚ�ǔ��<éĽC5�uR|��g:��؁-������cv��W�UY-W�dj����Dy���1n�w��*ꠉ�x#����������kORl�@���`�F+� ��m4�qW@/ϟg�Ww��jF��! .˭�$B�i�Y�:�?��&;B�I��,��#���TF�#*-v�
2�	�z�X��
��[>'ǀ��m�D���8����0ڔ�9��(�;��Ԕ�a�ͣ�f��9'a�o	��n<(Ǝ��hԑ3��]���&@��$��ɍT�	�t��'��ɛ�E[$�u�R) Ŏ%�*ܳY]#/�߹��k�|�'k�e*�U%�����
���
|6T}F=�(c^uJ>�ؓ��o~t��|N6N��~��K���.�s �2ˎe+?T��{��D㌡���'�#mE{���C��%�t��RV��u�(�6���$��C����Qm���'Y���&���M��ɡ"�:%4H�����9W��7�>+_[��٣��������#D�����3��d[";��S�}�g��{��}��7M���L�:t�Ѻ Wt\����T-!~�y��}9کS�zumS*�
��)YϯJ:���5�Ǝ�� R���Tˌ*WRR��Ϲ��;���yr��H�V�RB�.�l
��Hzm�قj��O��;�r㬶��� kd�fb�g.4�hk �	�"�D�@@V�ԯ��-�:u����7ޒ�w�(�+E�9{&�Qg(�7�M�Q�tȱQT���a�ܐ�I�l� 8�|T@��,�����Dv*f�F-I*�ۼ�-�a[�K��n�B9��JO�3Z�91�"S�ԭ����gr9Z�P[9;R��V�9Jj��#?�tkw�[C��'�ɣә �#ӫ�:�nh?�(?���4�I�l^666xm�=�'��E�ƱV�q��ЁZ��Qn�Dޔ&qMs=$e���47�(��N�9��m���2]�pJ �i�a�O#�B�e-�+ d)�R_�u�!ͬFa�(�O�ySV4�pf�׃��y	��QY���A�)�6:x�{loo���1K��{���C�Q�V���O�a�)0ˑ��q8б`��Y���ڡ��Dd
�ɟ^�) ����7�䔢���ϭ�p܁�f��Jm ہ��qNI;����$��0��E� t���݌K�|~�c����y������:<#��2�g7Y07�ϡ�g�b9�Ie��[�Wⷲ_�E���fQ`E���%���=&9kl���&�^��㝔`-iО��q�ۧms��Y�Rʁɂ�Z{˳4�%qO�Ͼ�	R89����ns��M��ӱ�8��� s�)RA��cJ�r�G��Ä�W�SR�C �K����܃A�M�|&c�S�X����6<P���բ
����G��<z=W�=�)#Q.C�7�x��`�cd�&���� �c<�.&�����wQ.������������=?FXs1�^����0�ln�㩟m���١$�s
-�m�?+�v����x��k��8Xl��O�f�O���S6�������0_�b�MWs� bj ����s≿��kӖ���K/���}��hWj�]95TV�ȍ�L>���4BM_�	nW�~B�:jGAGM��dP��hLzQ�"Y�$+�#�������/f������o�rt4���%=��~����Qu�	��F�v���R)�r�#�������O�rt���]���a�C��l))�Om1�9�kK�ޖn�C� d`�EF�s�,�8�*_����}�߼#��$����Cq�4�xP�oJ������~��A�Q��4�iL='HH�4Bz�#q]y��g���~U�x���[��A�)Ё��O�[�TiUj5 S�!F+�BO	D~�Xq`�yS^~�l�z�ƛ���z[r����cI���]���V�ly���7WP�7)�*�\Sgp��*�Kѩǣd�T2�a�ɤ��\��]�v��@ᠿz�BG�~��|p�:I՘��Q�(�|B^��q�)ä�u�2s�2I䅙m�ޡ��K�����Dg��[��fy��*GljN�._�����άH�V���U9��HF�}B�Zi�F�c�|P�k6�mq%wh!az'`�ohڻC=���N�ǂ� v
AE�^,��xt#61"���n�?72��P^�Dmlp:?���f%��9�}���mP �o���Y��t�4����15�S�P6C�8q�l�E��GTogݺCE ���sl��-U���:)*S��mH��Y��<8O{�yrνd�<�-�%���E޺|Y.������|F�%�'R̬[����(�x����43�VF��E�Dw�}	i�|A�֪�"yF�2N�l��C'�W� ��� �X��c`������n��=8-/��cL��[�w�M���-x}���a��c2�q�±�JФ�'�	�a%n��Ž�١��F�0��@N�����|��[\�t/>�scE~���/�#w���a���8��I�	3zA�2�g��#+-#��b�����՞w����!J.QO-ɲ錖
�;��ڈ�V#�%��3�/r��:�"	>h䆏��'�W.��P�I���5Y��i�2��A��qN�9������d�����+`��d�c�9��}`�(M��뙐!C����ה��(ɽ��ɬmc�;����]-���"��yr�,8��:׆k������q�'F�'��0؟,�<y8�V��3���<����j�Ʃ��5�]D+�2+.�k�QV`�e7�-����Q�r臩��ڷK�|E���g��ޗ\g"�v(�ki	*��II��[�9�!��t}B�Y
r_}n�?��Қ�g-ɗsRU�X�?��NO��V%�ʪ�I���<uiE��3z�	���z=P�����+z�'Fv�6���� /�>�si��dFn��M9+ݤj=�����a^��ˇvdo�H�#4C9�
ۈ�E]gJ%ya�$_֝����w{�=<`s����侏L�<e��6��� |��ړ_�� �ZC)u�G�Icܐ��� �Fo��LV�+���#	z���������ʩ/�[G�r�(��nN�qؓAp(��9],Kb6�7��
��ei�;2�+��Z�P~�[g�٧=)������#]_�
�c��~�@Q���ۑ:,wlf!���U�Ra]��rt|��m*U���ɥ��)i���Р�����R��T(��K%��Q�Ò?�9�{����%��ބ�ހ�NJ�����æTuab��^w�2`VA$�iA�+Lg$ m/���M3��>�y��F��(��T^�|$c�q��|�}W.>���\�(�BU�}#���M����?�^M��ɉ0���]�^ #tS%�>�ʻ�k�c7�Ԩ�&X�m5~FB|#��"C��譔%�{b:��^��C{D2q����8f
Q&�p� +a4�$nk��O�i��\��ǆqf���E��F�H�'���E��k�#eɹǆ1����=���)��S�4�n9�1����otJ�2qv�gFk���f�� /�M��ʀ�v3�Ձ`o3M����8V�d�]�� 2�t�v��#�1?�t����X.��XȮ�TZpc�1�����!�`����-T��쉛�8.�{{�9�9��Z8:�\3�L'���u���C{]y|�\y�]
���g������_����#��㧳�'��K�䘿�������߅'k~��9t�E�͇ >2j�C���x6�`g01��'�~Lg���~J��j6����ܐ����_n���@��G�6x�h&7�`4}r-@A��/c�X��Kˑ�Iy�򲫜��$�@��,	�{}e$\ F���eN,@����ѣc��.��^�H�`���������	�{|��%^
�#�37�@���K�Y��UQϋ��\�j���c���O��6;�ԭ��\��ʪ�������{���Er�_X�ˍ\O�/x[�X�砐t����%يd��=�����3�_��1+sJC�o�T��L��e��X �I���2�D��b���m|�3��z��I�aNɚ�?O��pS5-%��'/@��.�I�|V��)���t�Ё���a��0�D)L�r&�H1�*�h ��9�R�$ɟ�����kh�[_��J^���uٚ�z=z���wa|?]3-�q?��.��/��vW:�쎏A��� 8 �6�"�I(ED�;rt���lɕW_���ˍ3)ޗ_|���7Лӗ�ސd8�UE��krjmK�-9>���N]
E_�}�Ȕ��RI>�ɵ��d�^GV7�J]�uqo��2���޸���+e�;P0ڞr���Ԩ�]*�� ��M��H# Oz� �}�y���,gA�l��rxt$��@�CS��������h.Wt�_�z�����i�qܔ��ڗ^d9`2�J_7�]��,�Q�^�IO����`��V+���_׽�H&������Ʌg����du{�eC(���^\,�*�,��e�G�������킟ᘙ�x �.�!�
oyhs�W��F�-�br5G�ah�C�9�Gt�A��M���Z�<�x�c����:�ص��D���,��WMal�N^<�I�8�B��Q��6#ط3e�Д�8.�u>�sO�'\.C����[>�h����f>�~���O{��~������Õ�5��n�y�T�=��?�^=�F��/v<O���Dh�ߢ�H�7V�7Uc�1l���y_>yp�rm�'�h|������o�yt�ϼ?F�?Ṟ�����#��徃>dh���_{��}ˏ�X�O�;���豋�&K	.f�ۖ`f�"c�Фm�nC��Z|�c�~���Wֱ|PP,��3C�@�W\�DV+�ǃ�賌T9��q�-���fs���1��)6�����d	���Z�/A��k)M��D�����=9��J~}E��ܘ�e߅p��*���v5���ߗ�{��hȹ����rxP���q�zs���z$��T��yT��KJ}���g�RҀ���`���P��l(ń��͒\�X�Rf"�N��wS��;#9n��е�n����2#��8h�Jw.�+�y��Y��`��)�����߽.;m�$���y����$3ܗ���7��x=�a6rO'��W��?h ,�f�!et5=;;�{��\���q���Km�Q�;z��d/��/�(/��Js"r�;�FW���AAu�$ǳ@��S�Q?s�Tv��Lve�.�?�ų+�_�sE��[r�AC�� -��(��0/QB���#�
�RYIR4�L�N2�~�d�j%���J=�� �����'��{2u���P��b�L��lN���?�h�f�/=���'���^��l��R�K2�Τ����X
ٲ8�mh�%W�H���m	�#�f[2j�*+E�:S���_R|��җ�+r���e{c�ݵ��sf�\fN�e�ؾy|O��ً?È�H:<��E6��%rO����F��)� ]!�~���ɢ.;��S������c����28I�Z��?�>�xH[ !�i����_��av%���S��1 ���s���< d����|^�N�g����2c�N@I�<	w��?뉇c���8'z� ��ϧ?��{�g���L�;���r�CN@ $E�QeY��h˒,y���t��Ԕ�����������*�=�=�M˒%Y�s �^N�ݜO���>��s�K ���z��������������2�T���G�UI��pg�On˙رn�\�]�������պ�o��i�Z�vּ`��Pآ{n�!A�ژD��n���7]�8h�����]�4OR�������z���M�.��<U޳���/8p�_�ł����(t�	D�6�I���8��B$fhPY���m�m,Ӵ^���NP����)��ﰉ�Nom���dٵwz��-�ob�$bє���=�������Ѹ��p�=&��;I�lR��,�CL��ęr��<�OLJ���C,�`�!�zC#�����!;���<��e${��TV�����CQ<�ผ�k�2�L��gf0:�C����Q���{`�X�vZx����r�lwcv�Ud��f
�)*��N���p��ǆ���=���]���E��uKϡ|q��!8�� �^��r��h��H<*s�pv*�|i���y������5�m:Z9�*Y'�T"�DSJ���ɡ��$�x��CZO�t����e���ѻ	܌�|����*S�V+B>y��q�҄pM�ر�/�1�W
U�D�|���#����hڻP���ŏ�K�T%a�+`3�B-��o�`~��7��42�|�Tb�G�a۶zM���-\��A�X�� �m$�1ad��ޡ~�4��׬aG!���,.��\# ��'�?p?�?�ILέ��?�|�ġ�(��%�caa��?�=|?��1���0q�2��A}���~z&�_GilS�B�I�.���D[�����~����@i���E<=�Z�����*�se�%AFH���z��zkI*��r�6k���q}0�+I�����6=�j����6�"��������kX���1\�]=������-?{!>�kj��i�d�.;[�s�ε�����o�:޽��V��� ��)f����=��׊+{�p���G�u�,��z�����5�������7k��zTI*�������3T��3��0�n;�w�W�������z_(��͎�>��|��p�@��n����=��?)L�e*�u��M}�7�n���㊜G�=O������c{+Z��W�����f9�y�?Դm���"��*��Cd㸦�0�D�VX���[�ت0���~��]�&�����l,��Q��1�� b�B�:�؏�'�����0;�ZsdkݫB���GZ�ì{aG����I��U�0�.�r��O�ĥ�aD��
o��ihÉ8F��8�N�H��`��mU��<�<v�#,��w��_��Z���>�:܅lz4�,(�GƔ�F-�U�%y���Ak<y��k$�Dc�b�LK��^�W��������E�.�,���x�a2H���&��QT��.]ŝ��Lci�.��_�eB���RױR�������<�x��a���`�����m��,b�N}����`u飣G�s�WYB��*V3��2��8p�ITib�$����]{䄰@��ä��y�|Sӳ��2`L�ɡi��������H
{�G^Π�P@�R �^Aծc�I�ھ靇�X��W�Ł�Y$Y3��>�z�Q:q�{i��)�<��y,�h=]B?�f��N�i!�����Ea5u),!t��"B�H*�,u�Ul9ֆM��3?����t�B��
����ōjOu�J�n%�zW��8ؔ�C$�CtBSWk�C�4�@���WS�f�����q]���sX3������m��[ШMp�lm��7���6g��D���кˉ�f�Dl��x$�%O�4�gǧ␤%h^�.�-l%Ev��Ӟ�;_��ý���v����N�`������.[��[��l��7mt	󝂩.f~�]j�{��0�߸^�V����-N��/��k��}��%�{���K�e��� �����[j{�]��������������BW?p��鳘���6��d��C�>��z�R	y�g���J���[\���[�ۮ�r�0�+B/ԦZ�Io���7rͮ>�����*���Z�r�u�,�`����տ���^�~�m@�>?虄�^S�(J���$����**1 �1����<���u�7P�K�l��e4q>a`�q���~,�`"K���Q�X�UQ=y����3HD�H���&%�����r�a�b�g7�a��W��
&�."7{��u�C�8� ��ǡ൹:2����F���.�H|��X�E��<���h�xH�|06�Q��o����8��Ǳ�5QY�Gbt��(
�+ՠ����ฉ<���A^w΃��p�>��zivHS�l�8\�	�{��#p�$�\!ŕ�1p��,pe
�c}���9܃�{��1MԕH9���
��_�-bQ/�H Jxr2����	<8鈐��i�4�gӤ:�|��]?��D���4�G��^f2I���ə��h6ќ���q���&1B��Vv0J��@@w�@@��p�,�2�_`*��"��	fv�8��ݴP�+��W��?�>���]{qbl�+x���x��3�H��ǯ>�	�5�z���y�3聋���)'u�Z��q�\ ���+�>��"���3����wcM/��4y���������P��d���)�N�8y�f

U�/��m�H�7���.�_=)5���(�y�8��
P8���mR٨��߫ۦ2E��^��� qQ�M8�:B�-�l������pnЄ#�]�>D\�&?+�ǭ��>c��}���4]�s�)rrw�[�u������|^��k�����v$j7��=��~ϛ�y�����۳����6-�����܅��X8.\�쩥�1Ky$N4ËٙB��A���}դ.�ZE������
D�)!{m�^�B/:X)*�=��ڬ_܃��uԫ6NO��ޣa䘼=��˓��ӷv����e�x!�Z��f	����ݶ=v}�$��8�1N�z��X�Z���l:h+*}d�>��_�-�K�q��G0��/�b!P�� ���(�=�(�4O�/��������+-_wHeX7�
1�"�d�+�����F�)Q͝& D�����"~l:��7F����V������&�#�>���m��$b�JiX �7����YX�k\̙�9c��糘�ձ��6�e��2BaV�!e&�`p�Rě{03O�q�:��*j�����"�d@�=�J�&^G_�Ķh��n���F�|��$3NW�Й�@a�m@7�,���e�GK���FANq0��@��5���B儋����W�`nq��&bG��ٷ�ã�8s
�_x��S�x2��SA��'���X�R�;��J���D�Au�Ź#_�L��P��<v[��kE�	�[���V������y	�>�~�_+��y]���2�eͯ:�u�Y�N*�ۀi\U�U�)&�O��2�]ͫ�L��Ju�������d�(o��^��J�
�_x��7Qϸ�1�P�� ��|%	&�ު���\�_��m���#�2��jMIQ�7&s���^7����6Ӎ��/o�[����)����P2�*�Ő�r��^i�;}�@�?�^�٫K9��z�NX��l��D�h˴w��|�QTX���1Sh�k�V�6`��+E�ŋ+p�%q4]���TaV�C� <��H�-Ӛ8S�3���>�kb����J�J�OĐ:�g���~w}��(��Y��ÄI��PǙ���&B�JHb�?G�pp�S��4�F��$ݗ��Ɯ�\��*�:���ŵ�ް��䰑7<fy����%�^xF���B%Ͳ>��X�ů���3����eV�\]�k�o���p���P_
�4eDKl��,ez&��� Mb��2M�^����#9Qv��r�����&D��i13|S$�X�#I��&�s,��I���;���h�l�BQ�K�|ᒃ��|���R��P��0�0cH�����=�F�)�9q+��o�]�>�)[�
m��.��d2sHٍ����Ae`3.�R�ćzpd�1�x���gQ,UO$b��-��g?|�{|��PM���� �pom��6�~N��<2�(KXA�˄���启e+Wq����#ŏe{�q��dx^>�SσЕ�EW���M�Yszn{�T��2Ӻ>����
�����#��nڇ�ylC[����x`�'R�Ն�GC� �W]���u���9O*.)�.���<	�Aܲ��ס��m��� �z�C�����./� �R|���/(K
fH�����߇|4�����<�_>�)�N��͌ ԓ�ΣG�k|��w�GPmj"�Y,�'��4�H����mN��^�+/N��[�̣�^���8�Ǉaج�� �f��
bY���Y��
���+�j�k�e��gp��'p�W>���"J��;t;��}����w�����Ǹ���:���� �����0�V�#�o�C�+ٸ�ͻy��H"Y�3�~5��*$)���œOVUM^b�bF�8�S�IX��Ũs�Uc2�@��"�z`�ԐM��8(���G�ʍct9k ���݃��\�͠T��%���Yk�&:�_g�z����'��U��76�����XIVP�8��*�+y��:,:ڵ����u���F�0Mao8�����	�B��8Ÿ4ߥ��đ�.���T&.����D�(3w�{m
Z�>XGv!����~��O��b���_��8v��^��?�k�ńUm�$ӭn[m��'�n����L������g��U�U�F �s��϶���l�q-��4(E��|�5q�y���H��U��n㦫dn.f��A��*�j��ڟ��9��Mw�*ՉHr�8���=��9[�%�S�PF���
/�L�0��}Ț?����y�I�  �5�>����X-��FaP�6=ih�h�c�{�4�gO��X�	әya���=��z������nԴv^q��^N�z�Ɠz6i�	���2�p�c�l��P#�f�B*�����@��S8�[���%,�Y.��"�#�"��c�.;rN�uz=h�-��y���Ӻ)8�e�^C���u�(����J�B}8A�A=Y��:T("e9ؑ@3K�9����Gã�#5� -���D�k���b��C��aT����40|� �TtSM�]��!������r��5࿓�O�q��$Be.mv�r����ج�h{m�2\+����a�J�Sr�%[df�i�@U"/~ƆJ�X�xa+��:Sk�&�)ۈ����*�L1�^�ʐ�'T�0/������Ц�s�H� 4�;b"GSh���L�5G'��C1[C���(Q�B�������*.U�b�������6�3k�&#�`�QiT���p�4����`�y��DF�*�ʇQ<uNt;�y��$������+��o�&�R��n.�p_��p��	a��}�~��u̞<��7��.���#�v��k��;�n���&�{��d�)o��;�<����=xtUx��	��gve�=9����k�ےOB���6J
�������HSk��%t���)U4� &�,�>;����Cm����д_�t(��7�v7�+�R�p,�����/H�En�y���m�� ��:�o`�R��~z#@�����Ǩ���7�do7Ȧ�^K6ϐ�:]���	�t\�Fz�.̆���9��4���Ui_��Vn;pO<�i<�����GR��*TQ�\��͡0s�]G��|]S�Iq�!��"�D��%0>���NQo��O�\���~��Na![E�����?�[ƶd�B,2�%�P%�``�>�fqi��0��v�p3yd�N��a�.��e��(��*�W�`ұ��<��_Dz`���S��#�૯�-º��r��Z���e(o���ta��0h�7O���%4+W� �V� �%���$�ڛ�r��%y��j�@�@�ALK���1�0��א��E"��8A���(M��{ph�ܱ��g�NX�4��4�ͫ5�w,�Ū �&�O�T�w㮁�x{�>̮,ab�
�]C��!��H�j����**X��P�D{���f�%ԝ
�#�,��a\����WQ�Sȣ'��4���6��4!�T7.�U�LL`x����^y�0�T��8���D`���|2 dߤz� �]ߧ2�'�R�|U���r2|������;%RO�0=��%�Z�7�����~~�+�x�4��x�M/|���
!ͦ���cM���(�'^����5.�&�3����1p�v���A}��n��d�t%�s*U�A��V����ƍ5��q��F�v �`󵫥?7 �|��{?j]�]��6ը��2x1��WO�,�<�xg����L6�B�����_�2��;�q�EW�W��<�����d3��t��L�m�Ӹ"Q�ȕ"����F"0���:���>F��?�1�&�Ο�F�cC(4���̧{��ѝ�'�b�2��`��_��RvÆ.��N���*�V�,P�
gI��k%�X�7�¨�.(��^��$�^K���~�G���j��v�A����_�;�0.�l�+�fJyD���u��#��U��,�Q	�Z�Qd#Z�u� M`�'���Z�J�:�k��X%�]�=I���1�I����ayf��
�"m�d+�kz�\͘��m�va��GQ!�!�v��eL<�
��5���%����q��a���ۤ�e�x���&�&ѪJ���;�f)�l	��q�_4�La�W^�I"�M֜*�,����<Vk�=3�

	,��t�+�Ms;�T�5ޫ-�����]��zk@����lG����@몜0|i.�g��Z���k���DXM��2�[{F�A3�	^1�KQ��8-ֺ�Ӻ��� -���'��g I�o�a��z�*A����q�6�`�t�lV�%��|���V$�G?�$��@�O烪�@��xܺ��V����r��y���D�혀�[g)=��&�O\ ��t�����p*3����P�H�A������_�"���@an���1u��D�xN�&XZ�"6eӶ���Ǐδ:�rJT5��Y6bU\��09�*���>�G������c����]���|++���I Sϣ�)!L(�����`M�Q,��9��Lha�(��d%��]-ʭG��5��C���
o�W4��̷R|x�Q��7�u�34�c�7�x�Sp�J(�5�X
,�L�E��@s�6#�����K���um
7���J���I�nd1��e�أe���z��X<M'P��a)N �*��r�%�����;F��g~���!ܵ}"�>��fΞ��勸x�
�
���T�0�fL5�����b�zz��}������ݸ��1��q\8w���^{�%�VW�=�����w3�1���{�1J�=��Q-ĻԠ{h�*+yHU�J��
-.�{qܚ�t1��N�M%Q�E�D��L��B��H`8v%��\ ��Ԙj1I�����_||���07GA-��.հ�>w�.��n�$�0���#��
E�ւe�4N�-�IQ�W�,u	�*Z�VhM��u�|�]�²���qm΍)'"un��i�M��㭳�LrH`*���ŀ����\q���:lF�j�hX��XK�CϺ�nD�$��i���ݮv="*?R�ݰ=�B)�mi{�@�s6:x5ϓ��-�������ߵ�r;�������ձ�&h�>�/R��P����t:�d2���� ���\����l��FQ��}Z��赿u���mi��o�mB5�'�2\� �ӀѐIz?z�
�D7�_�c���_�S~�쳋�N��+��ܹ�X-���n���*#� ���|^$RϸH���ʒ��m*T�XZ)ȼ�--bfv��+��+��7��@z|O��������~Xd�_Z�}گ��Z��Y�c!�	/16p\�c,)9\1S�V�uk�	�)i��8�0c�	�q�a3��2����Z��@�f�y��r���m� 1��XV�a�/���&����z(W�tQ��߳qeoZ;��d3i�
y��`n��|g����QJG�M�G�c��E�;p͹U\|�U4��q�S��:)Oٱ�$�[!`T5�fO��_8J̙�@��f�YX���B*���F�kϡ}��؝��C��Ï<��ǧ���/#I�IEQ��s����Ã=��OB'Pi�R����1Tr�TfrJ�U�蔥b��`�����1/5/֫�ޫ��X��rBuzy6c�U���C��'D=0
�)IM�u��)�� ����opۅ� .Eݷ~�٭0¾�XhX��\o]h�	�4�P.F�)�Gݽ����JY���v�orB��u�Jt�J�;8}��v�z�9��}���^�`r�mE�r��|P����g����[��V)UܺF�G��5]Te���G�p��=�]A�赅D|쓟�c_�ul����?�k��cqf��LcZq-���D(�*���a2��� �C�FH�Z;�u�/v<1���\N]����*.M]��&��_�*>���c0���_�f��0<<�����^��±X�~�X�	#�x�;���+Q�r�C�G-N�ZE�^�w0*���Բ��vN��8̃d5Yf�]Z�>��!"a��$�-w��X�:�C�'����8��`�nЄ�Al{�x��_ű;��}�<��'_��SW%ƾJ �5L�F@h���?8s����%�2��*��! ӡ�Ϝ=����'���������N�~�ydi�%�$�����S�ң�e��Zᦺ#�ڰ�c͕ܟ�<G�H��9��g6讗d�d{�nQiͧ���+o���R���`�^Κ��y�,Mͧ8Q�[%���_~:�8�4U�
�0��ʍ�x���6P�H�~Z��
d��I;4����e�s�c�l)j8��W�o���\��[i�s�'��̭���
wT��Q�05��ү��n*o\oq���/��e�\A���?����UXz:4���	(�0N-��ͅ9)@���<�ۿ��wƥ�_��7��W_����,�+��d%�
S�1=��8J�8�쑭��6��J]���c�_��\�Y��$ͫ֨c������)V������|���+����+�+� L�Ǐf'�ܵO��,��MD-屳[tP[Z���[�e�
�1r��a��c��7�]lJY���)��԰�РIU>,1Xx1� �J�z²��o��4du��|Xm�U���<�{���t��]>I(��cO⫿���Фe��i���1}mW��#C�ћFh�O���	��r\��Oy��pG�Y�
Q����P�\	�XťNg^���
|�q<q����;���1w����#��G���Xz-Q
a�P6���a�&osr�um���Dݦ�DӶ�p�N�GBI�0Md�PS��a�C�Hq�CT�N���/��OL�T�E ���W�ͧ(������Vp�*�@����OqF����:���|�(]�<��mC����f�kK~�a�m_��8ݔA��(c��`/��5��:�y�nw��i��;��R��}�ny�Z�p�^��B��ٸ���)D6%F�d��ś��i�v�`5���$�	8�0�/��Bnn"�J����݇/�����m�����s��,�&��X.�f��W�Sy��d��!OKq#�m� ��Ԝ����G��)�r���>�`]�P��|��y�L_���W|�����/��I�$O!�,�����b{2��.x�`����Y��� �ꦴr<��N)f��c5�%�0Ե�'��)�5�@�d"�p�}f*�- Oc���4<ѭUrk� ����g7E2a2�m<+�T%�7�9�1 �B��Ǳ�������������~�c\|�4^.�C�EG�\����Ȱ��-W���dMC�~���z!w�Qo@��h�M)iN�`.]�����~i
�}�Sx��'�����S3��'hQ�1Ѭ�0qOz�@'�X��	�,ɫ���-�An�"V4��	Gij4�`"���9�9���t%q7j������-$knr3q�p��̩�C4y�d�s�{y��)�q}� @�;�T�xBd�<I2���H��0o��{�����w������k�'��,g[mrX�"u��尭s�E��rl��NH�9tO�ҍ�x��_���]t,ϛ�<���Npn�+P�UH<juy
�Pف�����nZ>����jl�˅�Zn~q��	�� �!�K�X��ul�J���x?8 ����M������t؉a� ���9�/���`���X����ql�^L��f�Jd�'�'�DCB�19Ϯ.a�D8.�Y&זUp���[�ys	�q~8;Ql!^v�^@�D��[�1�m���Ŋ�?�"�*�������o~�/_���� �\��C2�
��eE��D�#�J��%�6����"DWq��ܱl�D������I'�9�!�a2dN���^O2�d:�<]T��n�ŗ]]@�ґ7\\�f1G �h�`����*��旑 �S���O�._�<�zL��0������;>����y$�MW� ��.d���k���b�����"�>�:J�"�?�;�ޅ���W�JJ�fM�jE��1J���+&-���S��E���F�/���S1���j�~xc��`m�d��V����ɮ�m��ۣ��$(o���]R����[p{7?O� X����|]��m �.=�T���s�2�{�>�+S��j��՜�74�i���"Iҵ��u}]Tԝ��6�C(g.����ڇ�����|�%���fa[�J�_�K��@�X��c>����e��M�I�4�Y����������)���������n]��҉�C9��IU�fC :�B8�L���[��,CQfIhJʘUW�Be�2��
�2-\����E|�H:�O����|���/�����(����_���	����9M����X=��V�"xA�_�'�[c;�������53�v-/H��Bl�"f��C��{�|v�"ξ���d��1�U���,b�VW�����M`�cx�˟E�&��?�o��:�W��,C�T�\�5�$2",n�W���.������D�+�Ń�%��;�D�eܸh�Uq>�귭.�}S�9��[��O>�˓ӸHhިA
'��0��$h�ش,KP7 ô�=F &�vᅇo�y=`�]�
$�� ��D�N'm|�� Ň��{%�:V@����y��7k9�d�]?�����aS �\�o wx���{�a��	2l�;D�{�C��� s�廎*HZO֭ř'E:��) ��T 1@;�
�����I/pq'���3g����>j�u4n7 cp���+��6����G��u��V�{�s��y���C��D��Y�h�K��q��,��sd/�̧�λ���(\�C����VF�@
Q��I�@��5,�{2��!�#1h���Nѿ��Zi��� r�V���h
��ҌtN1��>dsT�ӏ������C@�F*_���|�w�Ã@?���bzz�|�����KS8ܿ�$�Ŭ'gnxs����>ٻ���F9TN���9��)N�VnM��mS���/��%\�0�#����Q��Y�H1�b���:-������'�.��J�*��|�pպ��{��/�:�{��_���x�K�Ҭ�֛����l*���3e��.x,�E`рr�[��o����Tv�ѻ.���Н��M���w��æ�}�^�'���ԯ��I��I�XO��2����qZ��fU�-�I����H�v���!�Iu2&-(���]L�lU��}�9ޓq{�-6k����)���i��N��x���չyZ�K�[B4���J�6 ��+�s��])2���?����k2�:c����?�m{B���r=O`��?>�� �q76��ד/{���_�v��;j�ll�n��܎ %?�޸�v#o�8�o-�n���v{��y�����D�x�!�L#C6�J�"��%F����ơ������7N"�YƪV`^4q�X����=�<���(��:���z�j	�?�1��݃=�w���_��|W�^����X�8I �A��C���F.1�$��G�^����M�==����s����>��q�����۪f�1��a&ZE8%�B�\��x[��������0�C�����:@^;)Po���!�PoT	l�	�4����طxl Ca����V�}Kk����<P�dP��$ڗ��z���j#K�ڃH�n<���q��q񕗐=}��i�l�pL�[,n"W+x`V�@�QC�'%h���4��jM<�Fo������֊4�z�z�{��\=�s������RkH7�!�jo��*R#�x���S_�5<��'[B�'!�j�V�Г�ވ�4��F@2c���qbh�9��(W�DK�B��J��s�Ɛ�r���~�x�Z5�,����21M/�Xi�����;�����_�JU%]�u������wyaz<pTf����h�U(������x�����u��U�y�'#S���
�c�8j��5i��AR�2��GO%*҃K����%�9���ut�ѻ*�~^��sU�,�M�Pk�w��j׺M�9��б��U�C�~��z,u�t��e��gK��M�f��������ۻ����Q�gڵ�� I����<���f=Ofp�}m���"(����1��~^�VV�4%�W��D�n!B�v=�V�x/�ۆܼ��۸q:�xb�o�Y{Ӿ�DC@"���"V]��I,;�>����02U̝<�������}mV��ׅQ���^�m�Kc?��E�@����o~�װ��;K��k�a�P�V�]�"��
ξ�:ο�*N��Y�
zba��0�B���R�$C�`�Xe��&����~������3_�-�����x��z���t�mC۱M�C+�S�ǈ�D�^�30B�'ےΦ�zH�yE�U��������l�^t��6	X�!�� ���F�(7�k�@4�{p���F_��&'���u�q�y�=�3�{�M�OL�B��%�J$mӃQ��f���a�N��H��@(�`7¾�!�ڳ��q�36��w��y,�-�ب ���7L�y$I�:�����(-��-��mc�q��1�q������%tV�:�49���^@'��
\#݃j�Fώ�԰j�	$A'>����ˣJ'@#���Ru궫r,�s�p7��y/��!<9�K��c�ֺ��@��5��\��7�T8�۳�[�-äI��?Pn��#uW��~dv�|���E(���60]	}+W����u{:���9��?j���G�~�@�~��5��Ly���9����ރ~������T����*��n`ޭ:�mlN߻��G}0d�5�,��ҽȖWз}GN܃�� ����X�p�Z	�A&�;a�7lR�4�8J�����޹����->��_A��I��m�9��F#��uz�����bpx�����d6�#۷�G����u"�g��k�x�⮼�&*s޵���'`5�d�Cd���jeZ�S�������+�*�M�� ��/��r���Z�ְn6�^�X�� /�҅���W"�cr(��:RU�&����9��.�sd���8�l��aW��������Q�{�7/(y�FH&U�1����0�Rk�8B���f�Yd��:v�}�Wp����I�	�y�B���.�9�3/����G����Ib�L�'݇J�$F�F�@%s�I�R*�ڹ�9z7v>�8���SgނU.���$�@�3���V�V2a)�$�x�=c��0��0�E�j��J`��E�}�H�ch�>43E��K,3��m"lq(�h�<�L�{^���ZU�~���h�%���k��{�4��@8��m\�M���� y����&ysKM���������P�ghkȮ��Yy�߰�ޘ��~����6&������o����m�m�]�ꓠ�����!U��irN��qm�Yt�W�Mw��w�Ǎ�G2�h�ҔHAˍ���l�ew$�?��g������o���X܈~��������y,W
��_�V���}8q�(�K�x�udX���g1Kh�"Mc�ôa4�.W2��|���ϸ��Gi�È��RI��q[{=�!v�x����=�¿��q���.�.���z��ҫ9��1�������i���3x��~���	���߅U�J=A�T�lv�z�谘��ѕ�`><����G?��{���о���#��X���� `S�g;J�Jh/��"!8�&�ov=zlb�y5����ӕ�趒3kp8���'�K�M-�]�;q���Q�,���ϋ���a2kx�T�"���lT��$�JCO$qfv���{����y�Ah��R[�L�R�5e3�`<��q���q�'>���<���o�KS�84:�4M|)���M�&�S�a<E�\���N���'0~`��q�_�F����_ P:F���y�ǊNt߁C��Ydr��.��T�D��8"���8����c�\��t
����{@U���*[����xl\/�ڍ-�zI��B�F��f���>�uՋ�E�j��kkIJ�ka��v�6�z�<��J�ns�$XEI(d��}�nck�fU{��L5�zi,A�֪@��\ף���`���E5�gӽވ�Q�:�-��=��}˛��0��+M0Z��ۛ�נ��r�����d/SQl۳Q���X���
U���.k5$D��,6`똸:�������?����v�rN�RRHa������}
+I���B�c!64�/~�ۘY^ĳ�X��g��Kj}1���X�q��R�_}O}㷰c��{{�"L���m��V�%쐢~j���)�^��p]�/=�:����@�k+�Y�s���䪟]w�����b��˫�e�b�'��н��L�!�VX%�ښ�"�N �AT��+�h�
i(C�&'S-b�RE)j��J`ۑ�&�s�g�#G@���B�ς��QoԐ&pƹa<q0C��@�Ұ�_Eb�n���/��O�tR�A%�s�B�P��P������܍�}{! �'��ƕ�e�����lJ�\�"E�e��4����8�����{�{q�����!V,�_"�]�	H���0�M� ���qi��$+6½=���5�=�wb莃�؏��_�S��ª#=D �e�<Մn#���+gN��]����V��O�4<�����W�p#�I�N�w[v]�,�<2����ںG��sK�m�q` k��M/�l�uB�2��UTY�W�k_�y;<=���i�{�� =?���x��r<ڹx�/o�dw���'���{=�S��A�ܺ��}���M:��Ѹ�麗��q�Ê���8����%�!�q���{n�z��X�OV��`zÊ�T�V�<O�Ã�ҾV�N��e�ٗ(�S=i͟���p��哊���9�XZ���͋f�Q��.@��T�v�`(�VtK���%�	�O/�v܏��4ޚ�D��J{�%�j��C4��xT��2+y������q�C��n��K����^Y��ߤe���]#!D�^�q�|㛿���9������S�K�Uw���z�,������O�4y=#�عk?fQ�TP5����"���"����Ը��rv�{��4���5M�@��,,���M=y��eq�)"J�1��|
鄫��X6LH�����H������5Y�l�L�J����`j�\�$�Z�˨�0|�JS��'L=02���ăC���w���;��I`-�*=8����y}����(�v.�G�7�/����T��������Ɓmc-
��b�Ώ㇣^���oa��=�w�.�;zgO�����3��+����>�X"�F�����R� L�{��D����K�ú҇�rVX�Ȏ�C���PY�K��l��� ��Y��f��_.�^���u�ӼT�����l���2P�v:��o�����:U��\�R���v���������1o�j���V>��5��S��G�=mB:�x�����=zn|/s E��z�΀p[�q��`�Y�ɎfGX�b��-���m� (qա��r[�@��F��S" /dJjv͓D��!@�#�M�K��cHR�7�G��[�=N]I�����҇��[ ��"��&{�\ęp.'�gJ���Fֽ?��K���)rd�Qf����P?��sa2�ϝC���frȒL�ɂ�u\:}�[��#��9�E8�����Do�yw#�w�_�"N��9����Fa�g�S��m��'J�t�N|�7p��](�ue��a0����hy9���#��J�	����v�*hCn����yLl� �Y���\��dhh��^X�ab0���?���z��Ĕ51�4/��X$�~ǐێ��Q�&&Q�2���
��4��L�7XvC<<�x,��l�Q|�k_��#��dT>,:���dk��=�B�n`�d�ޠ��S_�V�f����A� Z�&�r���&!]�������+�0;y��4v�o�zE�{,.Ш[X5k��P�k(��t�54�R�9��/���ǧ�N�Gh>��t��*������0�G�袊:�n]��R���.�*P/��䝜�=��v��;l����e����v��'qT����a;:C)�l?[m�����E�ő���.���F����=��e)���hK��W��l���I��S��`��H8Y�4���9ᇶڞ����X��w{��8�{��o�m�C���M��"FXF~����t��\�8���K<�a��Cn[O[UԷ��[�>�1��y��w�yFu$�q�=U{�Y�!����$z�O�յ���赨Q<;�<�r�T�aGY����hпe��t%WK3�\����~�%b�xmnvV�� �X.�V)�W�I�@�n�ê��XDl�D"$��9n���R�%��j��$����162����pm��p��W��FH���L�hl���ǮO���LUimA�U���<S�G<|`�Х؁{>��y�����%���öT���i"x�*T���-lԶ؏s�$�&��)H�����ȑH`*;���pt�����^o����)��	�4/�F��p��<F�6�#d��b��Q�x�����3L�'L8���o���9~�)�v���ȿv
��Y��uRq�$LA��ݰ�D�yx��<���q ����h��g�ɇ���~�61zA`�+q4���7��3���7��C�R� ���h���^�z��R�
a��q�]�-/�ͷH�]1� #&j�8��ٷ���ke�_]���{q!}&-p�QB��w��J,j���oz@�	���C#���#��{6���O�ۙ��x��-*y@������t�ϻ���. ���Gz�/��X�iZ{̼d\&<t}z���6����Ri1��2<��m%�]IY9�j������3�b�\U�|����t��C��)�l�Gi�뛁��}� �v$��!� ����
#tzl��U�h%��_^9�����
������ת��:j�d�3��/� ���9G�� �wۜ���y:�#'�W��HNR4��_��|����Son�w܈���W�_��lH1 ?�N���4�X-(9?�6�ũ�~B&����[�y}7��{Ƙ���
U4m��a�S�䢒/�H`eee�l��,	4l#ܳ}�`J�1'�C�Ԫlϳ��k�fC���64:��Q-U�O9؅2
�K�-fШ4���g���^��܆�� �d��w*=[�7�Ѷ�7l���t,�/�+b��$�]�@���2��*��'	�9ګB����=��U��V�~�ֿ!�"T�U��U��sQ3���N(�j5��AB�H����J۹�=A >$���
���m��W��)�F<�>�	|���b1��Hf��ޔ�:�:,�@�F�| �e�e�_O<�J��*]��|��wa�WϷ�}����z�G�&��W�v�$�s��5u�ݭ�0�:�snY�Q;Kj�X:̈I	����d��P7j�Cl2��Q O�'���+=8�2	�ⴙ��Dp=���U���"�֤�ZZ��|!C�6�H4�R��\���F	�8�4l�"����/}	�O���$�@�d�t`x|�4�k|��2w��ھ�3�Ĺ�_�,m{ǆP��ma�Kz -�cΛG�VF"G4M'�%h) [.�H����Ч����G�$�.֮-�ܩ�t2؋��
�*��1�!9����pe�`a�0�A[[U=��	W�����E��=�v���f��a*�����|��ӽ�e���׶�W+d��^&���K{��5k��b�:�7��tݫ�5�� /K�{�+�3_�O�A�Ů��M��ϯ�*�4F�a��*�BM� �&6ݖj+�F���O���z>�e.�SWt&ż|�MC�&�M���`O���3�h0y�"QTkaZ����ô���'I�����r�4G��mѵ5�f"oL�u�7�6'�}�J��l��{�*5b�$�@�i�+d`�������22���1�$Y���
1P����%��/P�P�QS�AU��'x�$�j~m�"�F|:��b���������XG\�eL	g䋫��ѳ{���?W����cqz�S���/�Jǐ��!GEl4������^ezx�&�y`���UX�����$�ﵒT�:F����۲�������!����NޖG���l����`u�
Ȟ����^��- 6���k7V82���y��^�qU:L&�Y�mx,l�U���ڬ�v�ˆ�Y*����E�e�����D��2jS���y� �r��}G?��w';GA֎�!���p�.��堢��]YO�5`�N_b�Ξ�0q�#?/셯�.ý8��Ksh])y���Di8���4�]����1x�!D���{�l����s�!����M�佑CylK�R����i4B�|j
o��^XE�mW�D�D�� +�v2��d3�}>�cw����r0,�
r�z��H<쥚�s�>�v7�[�Jޛ�;��d-೧��K�?Ӱp�]GPY�CsuS+⽖s���O4{?����"}�0��d�Z�!J1��ǻi�=�����
�D�v�=5�"�ԏ���<s�o��h�}�Q�"�߃��޴��s1���s�/s�f���gt����F���/�o��NN�"���r�l�#+�p!h6�9H�3<�YA�ǔ��<]�©gNn�)i?�x�����68]0�����b@V,�}�e�x�M���V�JO��3ݨu�!K��m�5 �j&���z�Q��""8oHa{�N�C�N���\�1������#�te�R��	!��Jh�L�ըň1m0����]�'�'d+\:|���u僚]bbDySb#yvC�	�ˍ�߇����_A���"B�A(�͎g�s����to��ԉ��X�T��*˒A]�����P���듓02�qyt"���&"�5z��L�K�=yvC���'����T7��rLz�͚����KI�3�*S)>%����W%#՗������T.a)F1�%�N���Hp��\U�B@��4\]��ZK�����=�:��]���m�e�c
d����T�&a��!4,��"o���ϛ�O�B+ݞ>�_]|Pª������[��u:$�+�_^��_�p����mЎ@��=�у�\�E�
+~#���V������xa���X�����tڑȾ�9��K�ߖ5c��M�"L'ʡ���М���2��ǮOݏ�]�	:�m5'���[�"ZǼ��zy{�i�c!��9L�q+g&P�&CR��Z0lS��?�x�����	l�^���,��vaK�����d�fC9P�J"M{�QwQ�4�����"wq��Z�6�
4ڸY�Rg�$��4v�s'�<���������uI 4��6� ��y�����<��p+�/�|�*ҫԯ�U��d�z1��~���LҦ�D�'�m�A�~��>��<}>�s#��<�\���5q�G?ǵ���Fzw`dhh�B�U��E����x����2س��q�F��+�@�典_���NueG8���C}���gN���K��W�[�������^ݔ(Py2��s�~��w�����0Hn:�*ex)G����;��L�ho��:�Q(��C�"�Z��Ef����{/����_A�I����r��au�o,� �YΠ������н��1*���O�z��u����t�~Ð�B��+������J�O A�81�RʢF�F��衮�ky,�,�>8��~oqܬ�S�0��Ш�,C:�'n�:�$����GG���P�� ��������M;U+X��Q��zM�E��m�nt���O)�$���ij!S$�X��*,���H���/����ZB^,Ϛ�]��^zN�"�e�v�U�R�W�ۮ�ݢ���͏�	.�i���y�6���b���1�q���Д�3��DܓN`���7^���ʉW����x#:�8��Ѥ���f�[���` �0 ��	(����_>~����5n����;0l�Yؘ�'��>��݁��^#�N�F��ec��/x��L&�y�tJ�F��w9���c:��{(Цl��
Z��e�h<Vi����r���ߏ�ɵYz�C�H����D7pt2x��Z�~�3�6ç"���@6gߜFvu�Q��s�����N�:�"�<�>q�;�0<2,PLc��|���!>���Tl�ҭ���$sH�}��]q����Kߋǒ�H�؜�"���EerV�#�'E��\�SR��H
�G�A��C�c���P$��:ڸ���Ekx���v��C缱48��) R�Q����y�If����9X��G!���T�V�XE��Aެǒ(2��� ��^o}��x���!�er���gהV3��
��x��ٿ|�?�<�?~/��T�=�p*���(���ί 6��7g���i�w��[/�@�p�;,���6:��71jRX��p��#��t�`^�r�|�g^E��E�je�G�	q󆙧E�q3is/ϖp� �Qm[��W�5wX���2�k�4��#��a���5\��O�z�4��3�a\qX���@��5F�L��4�+��ދ��qD	�L���f�Lck\Gx�M.a�{�!���7���լ��z%O`���^����'�H 'D�I�Z�#G���gz���b��>[���(z�����C(��������w^��b)���v~�K��go���wE��f��%��,�Lb���~�	�G���4%jÇ&cˬ8o_�z����2�P8L���:�WP}q��)D�yc?�A�1��$�j�)ڤ��+��O�:��l�F��;�%B
�y�<���������>RX% �ח&Q��bͷ&1O�X;w��$"fb�8L��0ϭ��X���J�UB%������"�?��}���і�G��1���q*��fU\��W1u}��fP�����5DR� g,"[ؠ�:� ��h��Tj,Z�yn,/���.$>���~��c��ЭE<[ˍY*ͺ�Qa��U�4OM����dH�\�B��pU$�ݒ_�#�T�>�1�C)G�8]��8c��H�;�9Κ5#�)�|3��94�ι�{��w�W�9��$)O|��s�_R\�vJ�f��II5��#��|.��v���
(уI�	ڠ����`��3L��hm7v��!N�1�D9��2�p/� �xL/��ڱ!y���~6ք��Uzx	�zR�4��	l��������T��
����[����6Ua���hd��|�B�(Kc3F �%GT4H�L-�i%�3�N�b��z&v�v��!���� ��ǁ������1�,۸2��J���)�b]Q�(��, '����'-����ȫ6Ξ����Ed�+8xd�v q�8���gQ#�1<�Z}���׋�����^�Z��I{XM��J�Tտ�oݯ_����}EI���L��؊=$�Ffƈ�	L� A�3��8��dl�p��H�%�"�E\��fw��������߫*�ܯ�K�˦z{�U_}߽��{ѥ6K��c�~�@�K꺶r7	�CB�㯏��ٮMqI4������߽����T�Tp��'P��)��)�KRK'�|���o!��ú�Y�9-����<�BM��Y�o�b�� ��%,]��+���k������Q��;��[�����KH؊���1&���������>���iT2sѥ9l���� j޺E�u�|�@ud��.���+a��f<�o?��9���Y�ɺY�ܗG:R@K���X��)dv���Ij���s��Ve1BYA'v%��$!����L��м�������6����'�'�?v�9Dy|i�\J8D�X*�03}������ݗ��@���k��^8g�8/�5���kX~�f�}[��c��Jڇk�)#���7W 쀕�d��Î8���z�A<��g�E�m��)0��gn�n��!���W�cPΡ_]�L���'A���0<ڏ}�*e��4b���-�0�~�Y�T��w'���x���*~x��*��ã�4�f�SM̟� ���/L�od3�f�Q=�1j�/"W�*�vY~�R�b����ߪ�%N-�����o��-Y���I.>D9�b��_�ԯý2�t�����'i�/�mkF1-��*-���0.�0��ݑ/"sh;����bV�;j��%a�@+�u��E�(����cg���4.^F�*�����Ku�)g�SN��!�5��Y�Ϭ7*�=v��r���tT}
O?��p�v1�&`i��K����k�WN$r9	����g6-��^��H%�rb��؏���j�&@qC�n�_~���>��Ad��T����F8IU����?�omf���iA�R�A;t�i<�HQ�]�)�~nS�0=uΗgL 41��uon��!�Hګ�퐵����k^n�Q��|�ޟ��zn7��	|X�h9�����l2gdP��*nԋ���C�h���v@���tW��TyY44���P;�|������QCEnӠ,_�9�B"�Z�jR��ɸ5���=4�-���0�M,��n*�|�[�2��&_��1�8}=�4R)Uĉ7���t#�b�&������"�.�m��tMI䷣��m?�ی��%4
���:�Lt�(��C#�1(�ב��ГK��gO�����}r�,��M}���� p�\�&u�V��
R�ʱ�z��E��=Uc� V�R���^A�Ů�Y��e�%es.�p��%�QV��kU7.��l+���|�h=*`�j�������'NRiNd2�č�g06vU�_�G�a[S"K�$kY�/���t��\Gh��aX'.a)�� ��	��FtM��S�>��$ꂲ��`�Sa)���#n��i97X�Z�Ft �X����ߏ+ga����C�m�#2�@D��/�C���d'�+����Jв�d�T�{�U�]�K<�.�g2�	2��dv�!���Ә9~=��x�;_�'1{������ҳ(�x�/`%}㗮��s�`���+h�JHnBT�<���7�a��aI�=mmM:�`4��H �$Y�Mǲ�^tf�1��?���^Er��8�E��),�Ʋ�1�1C,'br��%ã�F~�����!�Ǯ���xl�t���W���V��F��B�����O�?���e�7�	6%��@V슖��ؑ�j��:��g��j7�ѱQW�ҋ/"���������D��gQ=r�3�ȴ�(���L�a%�Z3g٧$�664���}+�7��	\y��ٳ�?y��Ѡ�I	����^.݇�e��|ߌDf��}�0����͞���X��ԟ�5����Y��0׹���8�K3�5���J��Q��Z=1ܟ��=i���z�HS��q�ĄP���r�Y��hM�c��h_=�dqV ��a���_����0R��j�;e�YX�Rsb[Nۘݒ�ޑ!�#q�����6�2�l���YeI�VF��ty��z��W���Qf��T�l����R�8�Ru�U�
�|�rXsV�S�r��>�8����N�T
��{ݠ�K��+ڳ�ul��\��riYQ��/\���,2�Y���#Ymhv-��Ƚ��P[�{���3W����,Wȵ�u���k�^*c~f>�O�dlnw�Y5���YS&�;Z�ժ�K&�{�h��/��5������x�r�`�Z���g:��9���z��0�{�V3��s��z:N�3]m �ɿrL�J[X����u�o�z�pRG�E��TC�a\�x�� j�ôs[���r�D��Qko_z��Z(���O�?A�N����{M���	6c��o2{��a5U�8�wC>���X� �h�ϴ����;}�/�/�6/5l�_+:k�zw��
�T{��Ȱ�U�vX�n�4$����Kִn0���N�ʗ�*�蹷���w�#�*H�I��(ű(���?@��ILxE-c���S�Hk���&��ڈF-&�� �N<��}��7>v'?:�٩�\��2�-��UA�|#ٸ��磸���8������
._��Ͼc�.�x/A��� ��vR���*��	�E���1����~�*f��0R�u*1 �4Q���R�<K�Mqhv@���Q�H�+	L��6�����B�񃨓�}��P��^3~�
������p㕷��3�B^�-�_����èF<f����1u�\9z�l���H\�����(:M�����6�{����˼�V���X���wP��>���wN������ić2�.����.�����{ob�( ���3��0�f�$�.�L�<�<�=�#=h���R���A9fÚ�y�&��u�n��7d��?�on���WA��9�)B�b�im��Aұ/��0)9���q)�ap�(�O<��]ݔ1��掺wp�W� �u�3X�����%���p�#���<P��MO��2��9����ד��v��?o'XG>���9$w��3]�voؑg��W~��G���湮a��(A$�^y(��D*���iL��SD�v��	G]�+�h��`�匝ځ�C{a�c��c��6O�� S��g�����!z�iH �������Q�M��>	�c���٨�,`[���r��70w���]ۑ~d/Z)%	��$�g{T8�&*����VPʲ��+!�_s~����0,g� �;5Dd}:�3���9���6.�]��@q��H���c�������=�\
k�=lt���k��_�b��Zc�A��E�ʳE:u-�;��2����LR34�V�D{9	1Vj�-�P�Y@��nk���+W��E�
Nf��r��Ū6����c����gNaTl��<�\<��?�r��b@���j������Ţ�u���ԧ˛)P0~�ml��|y&b���A���͟��Ѐ�u,LϪ�/�_��̟&k�OV�kk'{���(,� Oh�`��fS��'���H�a���P9���Z�\v�je(�&u��g�r��
�'��1�G���n��a[6�S^�{���8���������1G��v'��T�l���	R�!a�+��1<�7F�F��G^*��v53�'"E�^k�jx̉jTJ�ՔȚ�QM�4��7�_�5fb(�<�l�HĐ��|U�M���l����C�e�ъ<:@γ%�K��He3Z��i#�Lz�5�Jt�Wѻ�"Ro!*F�)
dJ$�̡]�HA�&�"�5]�|��A�޵��A�Wg�⼯e�v�R�ɭ.�d
���-�>���<N�<���i��Xi,#����Ҫ]ؓ��n�Q��1;1��M[0:<,��`rb\�8�2޷g��l-oU"e���ًA�j���Y~��Z��
�?FvsYv�Ug0Yg��87'f�=,G�_5y6q9d�ꊬ��H3�Nr��N�F�"џB;z��=�{���-�8�	Y�8��߾���1r�ne��4����W��*!�Lְ��Ӭ����h����C[���#軏��d+%��j�f�Ϊ�	�k�z���F}�#���_�s���y����/��H.N�>?�ک�Hʾ�Ψ~	�G�"�$�#.'�{S:����j�FG|�NLU��|2	x�YY=?�y�o���Y��`V1�d�:j����	B{gd��4Ԡ���0�	T� @��9aʦ���Q�W �4�]Dd�(��J8�u����x��ִel IỌ�ѹWB�<��R�HZΓ���_m�����f�%�W�5y�G��97�B���ױc�ȧsrl��2u�8
ǎ#]XB�%�د(G��xɨ��#�`��F��梇\ےs"�����ɤ ����`�أp��sϨ��Y�F�T������Crn^C|��m���E	���eq蛟G��n�߀'�8/�`�#����m�M	#�H�b�otP9w�;`�bc-��D��,�J&Do%�v����X3��b/�"?W��9��h��<�rVZVU�%i+	v���_ܶ���<W�G@�'�P�8��c�$��W6W$Є�xG�@/����O:]6	Uk��O��X���`U��n�lY��{�9#��VC���� �ص^Aȉ���J�����^m�֭]�M�E�,6�W�W"�3-�����SgQ,T��Ob����Y�}���g��7?@G�;�"����;�Cr�)�_�ks��|�464�X�G����Ğ�e� &��Ӭn5���Q��ӱ�X*��G'����ّ!�?QΞe�B��ګ�uB�̆��M�֪x������i�>��O	m�	I���U�ͣg&W�PЦEm��좀�T\�U��&�u?��E�f���i�
�,M:A�8��KI�7ψm�C1���~T�����v;]K��V��k������-#8L��.�t��ǈ�c���u$r�iC�,"�4"qUj�0L�D�ԉb7.I�������̦n��,�-�:�TQ�RŪ�q���,�E�\�ηk�Kbv��v$�?���_"�)�{�<��y�I,o4�,ക��$�ώ94n��^���(H)�mn��D&��e�*h4oxy�)#�����c�v���@�Ѡ�[�Cv��GXX�C.����
8�Țǵ����#�b vR�lcN�k�Cy$S����\�g1:�1yo��3®�՟���lJ��AJTq���_�¹��\��M|Y�D��CL�ܧ '�/�:εh��K
��VP��TY�Csi	S�Ŗ�>?�H���;B?�(l���a����P�ҵqD��0Z�R�'�E�-Ƽ#�v>��PR@���
���z�^����SqX�~\�pS��ܓݻ�L^�}�;8x��Q��t̴��DE�ٕ)�O^DZdg��J�0�Zs�Jr� �s�u5���Uf5Ȱ�
�ܸ���Sc����<�S�dn]`f�o���y:�F��n��9,�8�-�Xq#?B��v��M"���6؁�d����Ѩú1���O��ه�tv&*�n��'kï��xgmm�oZ�`��t&'�Ӫ�K�ĵ[~���o6���j[vy��N]5y��գ�Ȼ�lۆŝ��(>�D��L������y�W�^��!��RE��)�M
��|�+�/�M�á/�k8��2Mã�}nr/�t�r�5�Oxoڥ��%�<;���$2�>�٨81W��;���nW)���}��$�s��?R[��A�dC�,j���	v��rf**}E����Z��Ͻ��5�B���Ĩ�JI�m˹��&�f%��������lJ����I^h�]�@;)�y�3(ƻb�n�va%(��5I��D<�j{���f�:�T�g��Yÿ┨h����6�XF�Wp<=� 5K,^��-�gА <Æ�5ks�r����;�c|���q��	�gq���=�c'?�9l��vrF�	�\5�Ύ�4]m�d	;tK��6�S]~8�4��/�S��"{�%6,�>�Ɋ�gމo_oہx��˧O�������$� ;om?�Y��.|'����q~���,��$�]l���gV=c��쫨�V���ʥ��f����JM�:3�$��]z�4o�����t~�dw���`��l�{^C7V��]��W�7q�aZ�r
�S9$If�ȱ�EQ�4Г�h�9�(� k��y����h'�eJv:�"hg'�v�,�ι�9U�PCuv�w�AvhT�&�Rmv*j�5�`^�e����,Zbp.
��UJ��j[�V��y�۟e��ϥ����	�0�Y�e�\����騣�)��<�H^aL6yZ��|*-�F� 6�%%g"٣�����%��҆;�͘'�֎9�:�9�I�G�@,K��T}<��R�-�h�xZK�Q�,]��m�v,�^ʸ���Prm����m�)ڔh .�?�BqNr=����'�!���������>س�&8�{�9X\Z@U�]с���3�|�"<��>K9f��f���*�N	�f�=$΋�ș���`�D��^�$JJ�cHeF��<(V$h��Հ6�S�(�m��J��n`��	l}�X����}U-1{���o�t��y��T:%T0�V���oO�`�Y��<V�mT��v�%51�L^�*ΗEl��Z]�'�:6�N��ݨ�Fس[�H��_�-=s�'1�E.V i'"�w�`��y��Ɋ�A	e�ŜP���qjeY���U�����ֳ�Ͽ Ӣ ic��^L��Yű����؁)	p�)?k�KD{C�.��ݾ�^�s����e�J���t���:�d���M�J�[ھ������l����n|Տ.b�޽@Э�I70�6�;f�ٴ�t�*&Ϟ�6P����JQˡTZ�=8ɴޔ�a�imy��)Aq�������5K3�r`t}�z#(ƚl�y�jw�GH;�|aR��Y��+��'I���*뺓��#YlD,�Ʋ��N� %�W�^ԗ
������Yʲ�3��IP���N��zK݋�S�\OM/*(�I�V@]��,VM���>��c��|�m�g�%��0���ҿ	��eX �+�%i�Q�
e9�eYGO�n�3��(8����;,(�1��Y�F�zNu	-��	�p7�����ޛ��Z�cc���I�l��v���j9k��� ���rm�;)�$��$my$��<S�<1��&�=���m3+�@��7.�����Qm�ˈ����bsE�C�.�Eqaӓ74clD<�D�3��<1�u���Q��Y�j������g0�<�m���p�����׳/����z���b���������Ķf8�و|NE ���J��� ǝ�ט�\�Ymj�T�/��\Ɛ�T����˜̧Qoxʓ��@"�Dej���gxi���\N��dD��yG��p3���-�7ʕ�GK�̏����v��ܳW����J�����F�:�����̀�A&���u�1�-H`�t�;;�5?[���<ϛp5S��d+��z}�V��D�ۨ�qE��z�:y/+�*u�Te��ܹXD���E���Zې�x���ͼ5�e�W�**c:S>�m�A*�$J�#'���|J�dT�vt~F��$y���D�Y�gr8v�� ��������o�+m8��f=E����pr8H����\;	Y�b������=���ٱv�ރѾ~L_</�bj�Z/h�L�����U f���\7'`���LWD�e�1K�ػ;!�H�t�K�Aɫ��.�z%�^]5���'��.@�F�͍����	h���BE����<�כ�ٷU�m�lVL�a��H"p��9��P,9L\�ۀ<�����D����J�����/��d.�(5�����&7�0���U4&� 1����i��|c��� t�0��(@x�/�ٔ�f,�l� ʓ�4 ��`i�G$�V�ʂE��,���)�A�����8�K����uT[h"Zz�aF	��}o5��< ؀4%�M4�=�#�(&�0/�f��M�}�d$&3K`��ꖫ�||�#�E���,J��ȁ}P&���[�ǵ��2�6F���vu�l ����������U�IA0����R_}ns��a�O{����^gf�}3m#`�:����ʷ �&dvQ)Rn����By�7��ʳGcw�]&���ޘ�1� ��of�R�)VgzAAqT��kU�d�3�����8�$S��		HO���ZX���=�����87!�!�B�w"l6`���U��{�� �3��ךZ�`��.�W0���g�eF�,?%?*-��${�^XV�v����U��4����GU-�r��Z)0�2���@9y�C,�2.f%Ђ� e��:��3�5���j�2BS�&��<�vG�f]�
�DMS�xA��2�n��b����^�T(N9���UkڀFʑ���H�:zN0����P��m<���r�@���@W֋�V�n��/�fL����B�$h{��ݷo���ݿ������&���SDujs\X������Z8�8D�^!�¸쟮�B�x���
�w3��0?3����D���],��f^I����G�X_)�?�>6�ށ�~�;f�P����{k����%�_ΫX.�W�ř�N����ϱ9�Ǝ�>�M݀���>f��#�&/ ���&��m�p
͍i&f�Y5�H(�#%�+'~=����2VoDJ�����"��k^b�����zG�G���*�wLf'��#?�\Mֱ�c��g���kY<5A%J�66RR�����sm蘘gX�#ъ72��LI6vU˵��C�>�DL��.^��7_y_�ͯ�Ie�����VP>�a�ۀ;�ذ&�Ѕ(ID�*W�8v'�zG^��mެƍ�$h���Hիeb��z��@�X4��)wA��t��3r����#��2Flx3f����@��]�~ t��T�|��Ǭ�����?er��L/��6��\8�$rK��g59;���ڗ�{�~LN�a�� �[
�����̤z�����������
��ꇵ��}�͐� 4>�F+v�����^�
	���i�-D�j9�DxfGi����J#��|���q�H�7���kou���KKHPc+�E%7���2&�i6d����;_�b�B'G3�,N1.�K��,��/��ӻM�� �^C��:���Ԛ̵I%�lw�[Yj �4���@B�1�J;y�LV� ԡc�Sk#'�(+��҉
�Z����Z)�<�!��׬�Y�5���۹�r*:���, GJQzǋ��P�Ʈ���@);�B��T6�"�r��k�7;��!��r9���н�F���Ŋ:�H�����ڦ�N�t|���v���(�0�cOY |����<C[ =�LM Q\AB�D�g���t������:�Y��I�G)"@#�A�uО/��+ &�ix���e��ܟm�*����lЫ
�t�,�HC�ˆ��د�����:इ{��R��2Q=��'\߆�(ť3q���}�ԣs�e�@��k˶jﴙ+�G��v���n�S\��4Kߌ�"�Gm�x�,�E����ld��A��z���q���(!���3k��"W�1��Κ ;�u�0��؎��s-<y�83> �����yu)��)��|rZ ?��#V��b/�k%��q'(��F.��~���5���?DV�o<�H��'ݢ���M�8�ٞ_�p���~	�$XZP?4ԇOs�n�J�5MKlPX^µ����/`�`��qq�u�1KI���8��b���}8y�#���`t�nly�a}�+�2z)��6�����d��1���p���?�o0~�^|�q,�M��)+و��FK���s��2��<���1�}:�[5�����e_�1d(�������X����rs�z3��$s���xȴ8(��9�������+f����xl��b3�M�TM�9��zڕ��CN���Og�΍]���8�l���](΍k�K�1��\`�t2)F��� ���|��������G&R�V�%����^f��y8�*`�ܐhЭT����K�N`0�CJAG6�5�h�2�8�me7#'���TµO�$d<�Ć|o$0�楘��I8zk��
�7F�]�h�[ݐ�}2���l����Q�8���Ʈb-q2�e�1<�׮\�v�>� �S�B�X©S'���η���{�cn~J�?y�9,�C�� M(a�\���r�;��T���i5d�Ia��v�f��H�a}�L�@�;�D#�����K���v與V����\q��C�qojj���찬��X^��î'����D:���М}��L-a�O�9���8Z'��U�fd��fQ����MC�:2��-��L�����k�\@#����Q=���J�&�Vr�*r?#O>�}O?�����O)�y|�ӗq�%9ۄ�`�[��&zߔMm핊��fX���}|�.�%���Ų'4�A�UL�[L%r��W9~�?A�C�D����M�I����V(�c���"5�v�ޕx�c��0�':wU놎(2C�M��]���--�x�
}�=Z�f�"#ͺ�e$`�Z D���Ֆ�%��2#�����n���͐x�VS��8�ÛQkX���1���'�8�-�Ɗ|Y�TD����[�A?�� �0�0��5YF���Ӆ��[ZlR�S����={�}l��[ka��{�۱��r�[�˚
0|���1�n�A�*]���p���yz$�w��{ԅ��@��T�`��-?��_R! |-����`F(��l�ec�~4J�Y\3nMv�ʺf����NkG��{&?M%w$0ɰRe;*��r2K�T4`È|���x1VAx/q��۰�*�U��I69P(��۴��f(��������\��f6�/�3*
�N�ub��}�n�8�W^~�gΠ/\of����P<�TE�����6������ ��Iyƶ��(�������o��/?��?�/\�`6��J�PǤ�1	f:�Κ?�7�T*��������m�e��\`9��8��ɏ���������"'�V�t�tZ ϕ�[�����,ȹ�q�~<��/2s��o�_��6'���F��&'����F.0�v�]�w�wP����f�� R���,�#�>������� �v�Ɂ �"Ὥ2� *��@��*e���1�	k��FM�#+/�*���О�Feb��{�e�.L�߀W�+в�u܌�b�[;�5y�i�/L�?�韢p/~�;��Zp�g�F����
��jL#B�ŮP���N��s�����+����d���kEդs��-{���];Q�|��2�2t�"Q�,z2#��A��b�(��Aū&�%��9��Q[�צ�-�!�jTI����2?j�<�%�)�GއhFISS�8��Q\�v�S3�u!�$hf�~��;�6����b�}h
ۿs�a�AT��ȤSj�"�|$�ь����F��^�Ak!0^�s�a�V=6�ؕ�q��������I	2\5���m9v@�5�,F�-����'��ŶlfB������xV�$����������*�5%���aB��ў^���U�
z���l#���"�8�*��ۅԓ��ܯ^G�w�|��5%��Ѡ3���Ƚv��NЉ�XF|�-M� y�(�rf�J�޹[^z	E9��K��>{��ͧ�Ry�-�%r'v5�m��a�#,$P�-=�]��ֹu�qX����$�:��^r[I	 �$��L�V	�'6�t�9P�� @��:�-�Q@4�t�ll�fH�L5�E�w��wM��X
b��G]ٸf����> m EvW&���j�K���rn�ʫj���/-�_/~������X�[�-49����^<����٨A����#���+5\�vC�$�ˠ!�A�(g�OK�*�[� ,O�;�R�2�k&���A�*��k�2��N}���ɮH�� v��A'QE>�c(�GF�������s,�����`�r
y����Za�#X;�g��b���%���P�SJ̌|�!�(¢��N��#�<�:tV�l�l�k櫳������"��x�Y��Ϊ��=#T�R/�[���HE�Q��X��%c$�k�C�6+ؘds�t��z��lW���6�������;��Xʯ������%8�H�7����g�^l݉�ﾇ'O�~K��v�f��������96R	 ����7G�YϯQ@�p�������3�S��}����>^���	���'?��F�?Ӄ�6�w(#���!�/���m�����?�������vo>�.�����s̻j7:�-/ᵟ���{L��}f�~l{_����7��Lv�D\ӐS�ې����<���@�o����5���?l��`�0�[����r4�a0�C�m�/X�H�LS5A�#��C1�;]�0S��(��8ײ SC�k��	0�{Ӷ�Ě���YmU�, I���YF�F�S%�z��LL $ů��@�����'�!��LMx�z���}��Il�F�Vɪ,��f&*�\���-l��p~l����������~	v2i��TM\O�I�sZ��0�+הc�#�U�굗��K4�0"NR'I�8X�Ҳ%�">Vje��Ɠ�b���|�W�/������s"�`-?��_-w+����`�s�-4�>h6q̘�n~�r9�5к�9��ޜ;�v��Ť�;u�4�{�}u��s��(1�@y9�ǎ���|	{�ߏ��'���*g���j�GC���ܜ�C{��Gѕ����F�h:A�u�P�*,�	��G�|Ks�ʁ�F��ĉ����]s²��{�R9�ĄsǤ�-/-+�
;�tI������{��E��,
?������{�ΜB��v�n����D�Ƣ�=���Ӿq�
ʱq���7��C�۠*v�J��r-�F��Qx_�#��,��.� �{�s�)G�?�>Z|�do?���}�k����_�e�fY�6��)Yy��́������n�2�h$2ۥbD�Q�7�A ]�Xѭ@�pޔ�� g~�Q��\Y�
��?I�O��T����C�P<!7�Uޗe��@V�r�b�-'�P	ڜ�B)fWT4�N�طX�n�*��wt�3Ymp`F� �SA���a��	��(y^��1^~�Nj�:({��㔞�JZyA�\�.*�Z:���(�m�J�"Ar݌�Ӓ(�s5&k��ϐ �x��_���1q��p�q�/_�������	��fzH��*���5���c��hX�X�h��[�-��YfL��`���"�b�*���Jo����y��*�m�ㆬ�G��صZ���� ��1�ǪFd8����ڲ��w&
ںbC[պ�U�	d���g�9��}��*��jNW����g�����E�� ��Mp�It���:1p����)*�F~f4i��	���<���Hh�mw���j�=y�m���P̣U.�?׃�ެ&&>���>���x��5�p������W_����u���?D&6�� �z��-��o�����r�z� ��u�~�8��c��<��Bm6 1P�`eZ�ѕ���~�#��V����P������͘�?Yz�~/��P,}�X`�}�~_�ַ��8��`��D�ki�>�5�p|3ϭ�����˱�l�v��"�����W�Ϳ�}��<FLD�ʃ ��e��Fښ%�1��뫰sJn����(蠵�3-s6*����J{ȶgFI^�,`R5�P�����k:�qt�N�<�/N�2�.���[E��Ԙ@�Rɠ�<o�.OL�_�/�������v�ۧv��Im��e mG �M��Iho����
��co�0zS�--�J��ӑÚ���#������ߏ��2��\�Sij^�܊�ю�޴8�Fzz�YҔ�V�~�Kg{F��0n\;0r7uʪt���]�HT�
.7u��V�v���ѣay���D�N.�Y�(G��[\��A%�RM��Ƒ�`��#���3ر}�nƂ����������|������]�$v��B�c��V`ёC�h���ҷ�٭,��X���fk�C�vYZ�̧�pRTۑ���׵A���֌
	�s3�gP�q�1D�r=�x3�/��Z=�� �J�e�nԴ~�����/aU4�^Ebd ��^���ڮi\��ns�
=��+@|�pvm��Œxzd� ȑ�����B���ڽ���k�%l��y!M�𐃌�gs��+ˇ~0F�4��x�����{2��[^�-��[���i����F��0��mޯѪ�� ��.g�i��d,MDs����h�"AV\M-#��r_�Zߴ�r0�Y��K�$K�@5�B��r��}�|��[��˽�eB�r�����Y�Z� E�K�DJ6ى���6�#��Ӄ����\B'��P_�8��8쨎Wc������s*�/��ָ�X�ՀR��7e	fY�ec�N�	KK�Ie���X��?SQ!�]Lpu=���ک%�{*�V�!�vT�Cy����8(Kw�����tn��`h8g)��s�٭J^��	 /�����9ێ��qu��iꪍ�g��r�,����{�Pl�$���<7��ӥ�8���Nxmr�)�*���AI�xҀ<6g�&�j�v����\+�59� C�������z�^���@+)kR�b��5���� ������|�2z���뾝��L�o+?�����X��\J�_�G��)yON>9Wp��`((��2y�c��ww��Y������{x�~��O�%�7��*��X�"�U�xr��2���ò|݇��y�]�ؿف^DY���|Yv_O^���s�4�:44���^\V�
�'���p2Q�͑r>Z䶏����wp?ܟ�{-xu͆W�POxg�im,jks��f��rH�hײ���W���T^K�V\�o*�w����O�nݵxD�F7�_�U,k���ي+P.�X�M�]Ƀd{��:�)�M D�����#��&���,d������+�1t��|�A���8~���a4Mn��b�y�,��W5e�t�k��g��������}<�F6mFJ"dK�>A,�r�g�x'�^����l��t{F��(��bIQ;�<�P9A�Uy1��[��Ѓ��_������;�FJ��Hi��QS�b�1#��Y��W�F���aF��'�讵����vmmSډ�L����[����0������uy_bVЮE��I�LRq>%�Z�a��e�	�tE�������R�i��صk��?:�N��_z�}��(fZ������R��ZU�$�ۚqv)�2-��CĬ�fki(#w��ݢ;;l`����z�b�"���hv�{�������bV����Q�{�Y<}��g�����7�q�,���}�Q������'��˘>r�3�N�O�t�j&�ӈO��x�5h9T�:�]a�㳰Ƨ$��'�<1����L���n��6����&�n8��۶�	� 1(̀s��`��{��1MP��ށS�)��D�Am1�M�`k��L���#��ý89?hb��%6�쎡"0��x�����6��d����&�I:	�t���%b�#g���w6_h61ۣsr۾��dI����w�@0,��0f�I�O4ʻ�YF-����(�Y�G[�R�y��ޝ�� r���TuT5�{���n�`�
G_��/�L��G�q���P��]�r�"���CHGS��UG��cXֱUo�P<�x-]g�s��
�Ժ&�n�����s(��3n�-.�͆�B��JL��J�c�Յ�1X��/"OΎ+`�4�ct���fP�ŷVA�mo��o��Lf�Ꝇ�){����n���l�d��lsĘ�d�y��re�G�P.h��۸������T4p,ō��N��:���6����7^@,�OҎ��R���^G�u\�6��s����b��M���� ٿ��X�̂��&��^�&?���10Ї���������_�.����~�(�j��e(9<#~a�,O���mf�%�?�����EQ��=C�vT~fZl舀����t� �ϗ *�L�p+�EQ�?%��s/?cE>�*��7��Ͻ��p�\ĩ���"$H�� Zw����"6=e�0P��ox6�Q@j��n�{UM�az�j�Z��P�]��F8r���X4��4֒����3�[t:1K)O	9<��9Ke�r�-%{+Y�6�t,�4ms,5��F�ʇ�udF��&�h����D�V��p
եg���/����q�o(/3��mDY��"�T`�|$��� �J����M�KT0��)���+x��[�o����z� �R���&�^ђ/#�݂Գr�#����#;:�:n�������_���-�.-_:�s�Ob��_6$�[�ܗ�A�N��O*����-y��j+3Y������h� ����X0/4�l$Ygx������'��%�Iűss���#9�r	����u���;w���䤖>��1�M3�s��0F�m���f��4�]�8�z�H;p\�e:a�^F��搐�J.��hq��	���D���sG,NU�B�C��ti˽e�݄�fxј�h�Dm�C��x�io����j;��8 {$�e���nA6هm�[0~�<�����q�Љ������F�o;f.�D���a�$�ı��\C�[1*�5��jԐ�.�Y�����3g��ufc����]�sӈ�S�r̎/y~������dќ�Cy}��)=I�h\-���S���|z�ƃʰF�]7�[�l���h:�H0�JƘ1�hG�M:A8�a�<�_��j�#��5;f�a��F�M�5}'�$E�l*K�7�r/��$Ktb�H��+pr��R���G5�v�}6)��eJ��fW_Ԍ^
��Ei68���V��v��Dk��؜��Љ ,�R6K����������*n
(4S���QY�*m(�t�i��d�)��� St�ER.�$��(�J0�H� \+qZ�f�S/�=ɜ��3|_����I�3��Q��{N���Ǧ%��S}8GlQ�=r���
p$3S�]ρFh &[�+�j =��˚Q�HW ���\����1�= v E�SM�:
d��CL�vK�|�x�4�Dͻ�^�庆����hv���VM+Ti9�QA�I����[Ac���D��� �q>��IY���R�R*!��QjLH+g׺fƱƞA୒:�׭����2'*����@��Q<(6���S�\��틏#/v}I�aarB�	^H7�M��:�s��f�(��i,^�	;w� ������v˞Z�zv�$jy���^L�>�������?����?���_�Zg���� �:��:��	��h��oi���ȴ?=�{zW� ��E�5f�]��,x ��k���K�#��I -k.k�2WB)��o�����!_ka��q��Q�j+(�$�jT�S����Q�J�M� �m'�2�PB�"��b#�
;k�9+j�X)mc<9xB&��n���H�+צ3�5� ���nܵ��Z�LSP�˱*ka�`���>��i�Zpp�QnT��<���v{��y��"�ǉ������6��o�si�Cj ��^P�2[��W�j'l�]C��}Z~? ��V2���g���
��#�:�ȓr�9y�1f#���3�p��Ω �L�Dq>�,>��h�x��wp�ãX,���_�
|�e�g1�ă�c#Fs�+p��y�T5à�N������O3V��]O�M�����P�����u����DܖF(W�o�w@@� �'�xTI�$G���FNG6d� ��|��I985Y�J���>�F�}���o�����N�J�+z��� �6�.]V�0P��-%���p�tG�`�2YM�V�gM�D'h.���xy�j��ghiS�<m����zc�N��rv�8j�o�Ǯ`+�C�hJ���,����>ԯ]A�����,%�G-�4�r�f�#�q�A��5N݌J�\��J"����R�L�A��L2��޼ey9Kb�ș�¸�Kv]Fj�us���mJ�t�I�>��*��N�1Rga��C��ʱ1Y����-3�Z%<o��T�o:�Z3�h���ݶ
�s���>3�������}�^]�.6�yL��M�2�S7t�k�KK�,ϰ���2��}Π�rP��A�蛮O�� p�@է0��������1X�N�a0�j M��w�Md��ܨ�Po-k�r�7^�lLY�#����^�zKf�K�&�|G3qq��e{�0�����If�"�Ȝ��K��P� ٦~w��6��47li�U�㘙��>6Q�C�H.�4ԒxD�z�ٖ.?�<؈,��L��x��y��3�s#��J��'�&��v� �inM|�Pt�m���s"�X9Z�z�����K�r�`�RA3J�ɱ�-��l��������9r��	�bTԟ��������g�9p?F7�`T��E���B�V=��@�{���j�~�+�@�QC� ���6ף�`�Y��q��?ơ��c��_�����7���1~��y��,M��l�U72ZQ	4bx�يԅH;�P	.3��{��b��,��-�:ǩ+����F�fN�	�����=����(�#��߿����
��Sh�=��%�>���_ cF�o�(��u	)y��s�+�1��x̢�Zq]>�~��+�,��@ՠ�q3��!/.nt���*�U^�pilu�<ĥs��O�Qs��M�o��G��h<�˭����<�>��C�p��'���L_�
��@V�n6!I�v��ɸD�54����$+?8E-"*twbʽ0�mʹ
���51�6�b�b�@P�,/�Sb����ƶ�x�;�Ƴ_��Ł���/1~�F6���y��G@��T�:���i�����L	nm��
ǭ�����`#ڎ�����	^�)��gِ�]�VowK�3�}���ܻ�=y��1�Z% �ΙL��l6�~>��M����h �=9ܚ����gږF{m;h�����u��&Z�����r���t>gލ|VZl�0�:�LH^��SHDV%=�N����+�Ҿ��M��Z;�^��w��.ʽm�%��� {��쬴8��[۳�cg�..a[����<�_ V��m�s��>��\w�W�u+�L�o��d�
ݨ��yȜC���&=��(߱�N'�M�Ȧ\G�?�߆�y��E{�� �o�6�ŀŚUy�F��uR�S6�G#H���L��T�v��n��.+�����{����*���KTkGBil¹�0"�6�s�x�f7���dM��`����teGb��-'�!$h3�D��+�6�BG�0�8εb5"b�1B25��L�'��ł:�5wTj!�<����AU�<é�=�pv�wd���p�^�'�nM<�KW�,�Z�,Z�L�S@�d@# FQ� ��ox���I�ۨ����!=�Y��� \�_�`r�Y[���;�
TV�V#�$6���$��Ć�[��
�%(l�M~,7�}NT3�QC�iȰ���}T�B��Z��I.}ƈ��$ �R�W �����	䔳{^��iw��S��˜E�0�Y-~-�+/LW��㭱�w�w�*�<57�sa�e%����Jq� <�$�<����2�;�Qr)%O_��&Ѹ��T�AʦF-OC��@
�׾�z�yn�$h���(����Z�̌�Wf��_�=F��s��}�	����1/�u���;�r�۞�o���-d7���+�
e(m�kL����:e�z���,���4��̦�������c��|�W���/?���1�7V�Ŗԛ�mt���]��1~�3�K*�rKJG�	��]�����&~�*l^�wN� Z���&"_6���T�����۱h/�-gx��	:�x�R�aj�R��D[�VZF$� ��~�������㹉	A��	�����Dg	���Oh�}y!qe^P
�%f���JSYTE�]�,�h�
$8��[� u.�M�.M�ilD�g�̋��#O<��8��܇GQkW��m�p}���f EO��و�0) ��AJ5��-�pb�=aF��O0����/�b���R�<�?�9ʼ�O  |�IDAT!���+���!f��!��;�I0��6:6�#�7��;%E%�qP���)�dսSdӌ�UFT����'�%�����[�#0�\��&G��[赕ۘH�5K��c�cV�:g2ʖ!��a�YN/,�9&Je�~]LЕ��̒���p�&���B��9����){��9�>fTmV��6J����-۰��/���&�x\��AE��)���5�:ؚ�m�yr�
"�#1_O��].b��ix�H�ۍs�yl��(���`���%�j$M8�c�`y�<�H�u�,(�Iȃ�ǴS��C�W��z�d�k��;�t��گ][��ҹ� @쿮�S��R$��(�A������n���zk������
��e��=Q�F��	���8V@���R�u�8Q����?�V`Wg��0ſ^�c2�!:���Ry�
���{�:F"�2r0�v�F�����o����V��rd5.Y"�w!�@�����-�d �8�OC+�� �Xw��uU ����[ۘ�?���N�l�6~�-4P[^�#6��X�>�Xʔ32$4�*P�#�Y	�����O?�w���t��f_�rg��HN� ל���:r���s�j'�\��̪g�#���Y6�D�,�그�8ns��X���D}�+��^;�e6
Xk7\6X*��E��^={�`�/�V�FO�����=�E����5�+�(���q$�V��I%𩯶Y���z�y�Wp�V���Qt��W1-��������mNq����L�<�A�����h�{d��Ɖp���(��i���>����FM�9�<���,�GF�����s��v�>��c���̎M�*����x���F{�=%����	܂BM���;�o�N�<WX�eЕͥ%(\3�� o5��n�i?� GV@gȰڝF�rkLs���G�A��6�`�B�c������g$�=���l���d�zͱq����x����'����7����71���~$忢8і_�C7�H�Иz�A�$��d�W�V#JI���(��a��e�V�Na�����,�88����o=��~�:
G�cjf����B	��b�DB9��닥7�uL"̸݊ۮ+�1�~8��]���������Ѡ����Y;6���J+�V�Vj7P�_۩�ѝ�|�X��'��w�G���9,�
�ƍՓ͠ Π�H�?5 �" ��K�Cm��b���}{5�et�ݨ%¾�
��j_�	�y\�@��y���"��}V��t����� �/d��+����H��L'�@��z�AYs֝�/��~���9?��ݿѥ�ﾁ��3^,c�_�$�ɶ� ���U�sR��Ȳ��Q,�S���(�m�j2AM���`O
'V0��/�����Ljem�=�IaH����s��ăx�����>�}�;����~�m$���H�$�����G|Y:��Ñ�f*;�u��dy�훃�u�"ؿ֪5�B�M��%��V�?��]�F��@��ay��Iq��вT8_��J��^���/m�dy0y��^weI�f�ym�F���1U<��c5�݇���t=�~�cu���do�QD]�����@��RQ��s��LS�[9Z1��A3�����*�M.n �"�V�(dN�t��̊�����D,���z֢f�4��YC�q<��]3)D�x/3��YP��S��y���x�~݃L�ذ��A}��ց�=G�u�t�`��������ϏI ժ�B��?G����Y��3�J�5%1˹y�Y�!rӶ�B����P��%���<I|���i}f�ʤ ��l����ޝ�!�T�``xC�1\y+��Z[������ۛ�����O�r#��`U��p����0]�?[F���nUқ"+\{�}�L��ʣ���"3�Oʹ|�i�y�4W�c�f#Qi��a9��r+$S���:�1����������/�&��<%@o��1�g�bsߐڬ^�錣����
Rј�y�|��۰dn�?�J<�o9?�\"��ƯNO��Kb����w��g���y ���/���_�+��I�A1�FϤ��-HɹhV%�w�)�ok��ڦ�Pe�;��7��P{)�����ɄQ����߆)ys��p���?��l�;�=��
^B�7˷�>[�M6%>\+�R���V>PF�m�8�B���ꊖ#�*>��aTQ����ķ���V�8����0+�iG����Qj��`����;n��7Ɨ�N� YӭJ����L`�4�
�Ir^b�Rcl�ބ��
/}�0�Ӈ�?�9���&fnܐ��G�����+`{<�L������j�B���c{C��m�Qbw�-������Q	]�PlZ��ሩ��{��n��	�fH�4m+���M*��6
����%��m��b�z6cwON5�,
:s �ĥ���]��ui��8>��R�m���g��GL�6^��1����t�.�WQZ[�9�LeS�ȿ�Ke��P��ֻV�C0�QIW	�m���$�5�$��mr�VJH��(K`Avyt�b�E�\G��qj1d�.ʅ	�Ɂ�Ȟ݆�s����X(�(�4��R�m4��4{� �{���_��r�sT%��:�s8��`�3�#9�	W?<���/ûxI@��eF"w��<' �뙑�=3U�<۵J�ث���q�kއ:u�o	�tB��5W%b�^�/Ze��I{�X���<l����Nu��zb�&�MR����Q,ĐN���k� @�<�5�y�S��)/	1 ÎY� R�8OM�����g���!�����ϝ���oխ{����������(lZH���U��,l�/Ny��
��O�6Q�3o�r�
�P<P�y�쎌�5�>��/R��<Ò`%��\��tv �4gT��zRBK��JV����D�o���!�=1�N	F<�+��h�l/�5ū���}��Iy�+�7y�E��e(�Z2$g���ѹ1�o��ѡ��	��+�m��8<�"�A�x�V��p8�� ���!��Lc��/M?֬t��%���j�w+E�x࿞:�ªϚY#d&ƐRR���&�[ZQPĈ�Id��)����x1�mqQQy�+�yC6F�}�����
%y�h�Ts=���;=�~����{y)�����T���рU�Ȇ�t�W��`S!�3�~/���#9��z�.��g��O�'���:�������߿������������~��N�e0Q��~�á���
������/�)�qce��|&��R�(�z�My�w~S~�?�{�������#)��/�����~_��<�j�7u�}|O��+;��6�_q��$��_Zs����.������7�������o��=��+�a|��x0@d:�!��)��
��D��U ����#�����[:��-�L�z5E�|x /�����!�yZ����P�4�������꿔�_�����?���d��Hn�	��U�@�9�u���M�)��q����	�"x`aա"-<\E���w��ɗ~����)�����?�c������hE}����W�\~mk,o���9��D?g��4�ؼ� ��v���R��O׺
ZD��"�̍?Rl�jыg�yۡ�d5Kȁ�Ux��xEbQU��{�"�(��/dy�3��,?���>���6ӵ�h�4ɝ[��(�EEV:��l�3.�I�<��\��cy��W؁d���#���ՅC� KK��W�U������rzb)���+��W`�!���zIf���>[�ŕq0�t�T&OPZ����H��I�����=9��ߒ�dWn�A6��
�'6��|);jd�0�P��U&E���R�[� �K?�X��*�H��ߗ��&`������N�|��,����+r��"��|)*%Kfr�x@
�d��2;!eh��R��p��L� ����l�[��C!k@ŖYg4�"w@��EG`j-M��7��,��	���M��.	��qd�8i���z���js�rhn�+�P9����"��Coj8���pA�82�?S�l��|5�eȍu�˓�q莉L	����f�  ���e>��4HspDЇ�v�|�~�����I{�����a��E�*D�mh7U��-���<�����v��8�B�������P��4���|�P;���DA �j��6�P����,�ĥ��@M�\G��8�a���z~�@w��F`c��:�l����[�w/v���9��솁����j�,�H]:�r���/x�Gj{z̆E�op��{���y�轣&t���߽�U��I�re�)aϷv\fI�W't3�k}�(��a��gU/T�2�!���$ĸa�Ѧ3@us�N)�s����Ͻ,���|Per0̥����������Y���ȗ���?��G��_~[��g�J�����CY*8|�H�节J���i�T�iY.)=�@��'���w�z�կ]~��~O~�k��uG���O�B���������.Y�b�(8:������Y>��Q�l��hc����~���q�	�.N߮9y>����|�� X/���� /��"��"Xyo���JXD�½�ڕ�<{%78���
��h`��z���yj0I>>�7vw��"��(_B�#����S��?��rp�����������L���;�o��ʟ��,����2r��,��42�Y��Ф���=k%�j ge�n��������ڿ�MY��������ߗ~�cyZ-d�h��VH3�[;�����	��"E���e���M]�.X�U�YR��E%p����	)3��F��9%�7mJ�F�+����"�����H����e<^�9��B�6ՃCI�@f��T��S��@7��w��ƺ��L|��H�ݾ���|p�ZY��/����t�r�s	�
j�:wH�l�����s����2���&lA��(�]�,�֎.�#¦���1�C���L�^�侄�)HU��Bԕ==���T��֠OLy��9�&2 i6��,��5k���ŭ��_�~g��?��~o �~����B^Fg��Y���8��/� ��̞*���͠]�����u����?��A�6W7�%��@EV���$���"���2�xmH�*�c����Dԣ@u@ �)x;���|��"�&�3p<��E�u)Q�P��Z����b%uzs� ���JS�tÃ��3�.�<y��Dэü�;X��@�
=o�֮�8�&�{r�� � v���A ���D�m�A^R�/c]��uY%rŪ
����w��m��vK{i�*6>�);۷��E���d~t"�dfQ6:�V��PJ)P����荢����E]��N[H��LmD7N�̣��6�$w��c_c@\:��g֎����<�7�ji|�Q��ɨZ��.���Gƌ���^�7[��)��*���B)��<p�
n�z�ڹ�{g��m@o�0���;g�A��U� ���=�E�:p�c���.�9Z��9JjW
^�\j�!l����D���Z��k��}���?��=��|�g��?�w~���7�)�?�R�������?���>���/��p>ӵ7��&�\'j??��w��/�#w�����Uy�so���ٟ~G>�����ޓ'�}&�b.�&F���T��}���}U^��/�����Z٭0^SMl0�"����{�8۝H�F��0q�a�c��Q���\h����[N���?�[,�>Zd�q��uX��P݄�A$�\
+�
'A�2����o��'J���+:��xWF��o=y$���z�����{��Å<�;ߐ_���%�����o~]������7ߗ�ѱ��J���br�x�9k/+FR��T�<+r�?�z?�������o��'���c)�����_�H��ʏ��T��,�����B�#_��t���_N�<��ð�vW��FL������u������ue�8�&�X���c�}�-�WU�U�z��_4w��O���F8P�5�u�P42���Ns�M;O���i�6"��9�GO�u�oء�Cԣ��n�x�tv�q���M�������6����vk�`��׎�W�۷��Ml�
uXE�Yl|�����a�׌�3���/���6R�;b�䘨W���t?�Ðb�gvFW����[JS9X��\������ñ���:�t ����D��*wk��0�������~Е	����j�������(cB��zm̈́�8Ec�'p�B�`��_�(��(��Y-�z�:>����Y�΃:F]�U��������7(��\��JvU�A�f��+�)O,hs�en���-����Yz�1"Z��%�K�05�@���.5:����ڑ� �'�߃�=	w�ҽ}������q��7"|����p��& �B�R]���Qp>0��I1T�>�L�P�I� ����'g1(�oʨOĵ�h��y�5s��Y�Fm��t�� �&�<���[h'W}�y$ �9����
� ~�)l(9Ί �֙��n#�mو�qp���=������:kR����xUj{ПV�?�(x�PVPd�ו��S�k#z�uZt|T�#���m=�r��/T��LLk�V��>T� ��c��� ������q�y�3�<����<t� 8��0��-&����ˉ�8fd�Y����o����u�h~�ű��B�u�?\J��pM��|�N����R��qK73'���j���u^3�QGoaz�T����g���8������Ӿߓs4$X1PO���M�u�T�u�@>�u|�`/��88�����$��]��3譯|IF_�
�q���~W�>R�|z*��T=}"G������no�p�-w^{Mvo�qP#��H��L��S9��/�ɧ��O>���;z G�ľ[ݣ���FwO~��o��'����	N�V���9b�y �]E;ַ�>a�o�{�G�s����L`~1��`�^��&�����L={�ƓE�����ۺ(M;�RmgE����24J~����Gs<9�f����c��Ww��{M7�����7���ى,��>y��ߓO����},_��ߔϿ�Ey�����Oߓ���_�������SἯ��,�誇��%�G���;==�Qi�r�䵯~U���G�������{��o[}�����@?�C=��H;�1�D���-}�]�DTO��X����2���6Pw��P-�?gE��]V
�r���o���F�a��O!�Y�����jd��a��~n(�:&GJi���#m�iYTvü���:`_Hv�,}:��3{tt�Q<<C�b�uF=3��V�!W�[����!�KkSZ^�� � �W�؝J�<���w5S1�������o]E5�9.��!��ɭ)0��60ٝ �D\X�Y?b��?t�!>����T.zF��l��ՃFjI�j���E\�ˮvOD�
HDT�����񤤕��l�j��f��� ���gZ�5e��3����U���*l}ʂ:����"t4 ��Gjd3����ۭ��F��ˮ���#a胋JB:-�&����0p�� �1��gxo��`��ᐹ,M�/ �:�T5��� SZ#�� sSD����Q��_a�hZ��.��X��AVm\�!ry�H�������lXK����4g��]���t��x��<Uk-��Y�ĥ�`������iQ;U�gKB�n��*��\g�̫]��iC���)@�B���
E4�&���l�w��'6ڗ& G�,-*ܡ��-��B\y����S�݃К��,�h3��~^	�l�4!��l��E��*��#���/�x_����Tf���!��+9|���b����o�ߺ+o���ŷe��W��o�%��2`_��M�����U���=9�Ƀ_�ß�/����G������R|�G/uur�>�]o_P��w����ά:��qA��Km���0'/0��C�3	��¢�n�n��Z�kQv������ /t^�/}���?UЕ���l��fR�M�+�z;�&ba���ާr�T�d(6�����i!�߷��W���D����H7Q���P���o����_��|��!�}����;�>�O>�@�u�F>O�<�_��=yx�3�tz,u�//������W��W_g�`�{K����7T����O�+����������<=>�e��բ��-�締����P��

���o���fCu�r"�A���F�7����Y+��yC����b���)=�ر�bJP�Ot�IGf z �Q����&Z�~/���bd���Zi����JW�
{\�r� ��E� qM�φ�or���X�Kg�ل`���<�Sb�n�5���6�C��ni�p�m[�$V��
@<8=�������Kv����qUD�M��"yX�'��(퀬�a�����*���z8z���Q�0����GϢ|�	�J������;�{&_uP�P6�AK�E����->ԍ��%�!���2%��
��������6�4 QX��}�/��9;{�����z���f�'B�^����F
�#��l��h�_�~��������:��[��Z0vm�&�O}�X�)${L�t����嗼S������.-#ubFI��$�:�G:/������gX�*�TrPW�-l
n`�����"}��s���mT��@E"�N5l�F*�S��um��I����y�MU�K~G�6��=e;�P:H�gؙҭc?���ݜR8!��D�`/p-�ݕ��*�[����!&UC�St���]�S&�h*��&r/;�i�K��%��Jr����=��"l�ȭ�^������������5t�J]�rzp(P��Me��P>�'O)�u�����;=I��ҽ��G��{��ŭ�la5>��Qm�f?5m�ĸ�z9���2pΛ5�t�)4�*�~7
�ky�0�9�o�<C�,o�B�#-Bj�+��
��(���M-!ln���W�P#Qٽ�UZ5n�
�'a�Q�" Y%�����|�ũ|�H</!.���|��Gr�����~"/�����;���o�K_{� %��t<��<z�P� ~zwnݕ�ݗ�}���>=�哧�ٿ����?����L��(�����T���F���vܑ�����u���;��f��
/g%�����Ϛk�ls�yd�N��EFR(�Y�~���ؿ�E���X�����y�I�:��e�G��pH�<�cC��0lZ*��������ͳ8���~�������1��ϟ�K�'�|,�f�Z	�Ӊ:���=�R��@�C���RQRo�{�2��U�=���F|�)��K���f���8�.P���$H``���#X؍F �H�0��6,�v�}���� Dd9�"�� rM�����-{~V���
�u�7�����u�~��Q��X[Wwn��*,�h+�>�}ˎ �T��4�r�5cuq����n>c��y�Xj�VBG�/]�,�
ov��&�����D�5U� y�
Q��UgS�$� Рc!Hd`�\7�)����1E[������=F켢��u��F��ʟ>�6h�?�d��֫w��{K���2�tʔf�:�@Ŧ-b7�y�<�7\KP�yhkr��jٛ�:V�nl�R��Bd�\yHG
:������2�z�����v����9�pD�i�o���7xF�5E��Z�����%��W��EL� K'������j6��5t�,��w%>~,�g�p"�=�sD��Bm�����q�GtrPDHe��Xd��\,glq�ui�E����H�
\�ө�W����;w^���/��Y�12W_ai��C~~S�$ af�Y���	fi�EY�������F�����p�z�1����aؓ�"�-�¶A@.� �f�H�� B�]5�7X�y����|0}�ְrvp��!r4��-T+���W�uE�?:=�NO������l����;-�~���p�{���e��-	���z��me|疼>~M�����GG���gr��=�t�������ާ��ၜLg$4l��F�PQ���������fW��KⰎ�:�l�<@S�&zѳ�L]\�W��j�dƺtAN�t�[��'[W5�_Q8/(4����qA7.�޸�ԽX7�.���DJ��G}yaw��hvh�"W7\Z�1hZ-؊��w���<<��ۅ��υhLxm�_�t��ߖ�n���Tz��E��܁�$�W ��Qr<��ڼ�:�0��BP}���<>����ق�#�s�N�6�������p�����u�N��mhsT������g/T�A�#	͋D�
���#�t����3�8\�y�i���,Ou�g$h���P_�}Ա�D^��(�*Z�Z�?�ds���wʞ��)�+3 �>ĉ3Wg�����;���t�� ��o�X�e�7^��/\g+X��C��X=�vK ��.����Q�3Ν����}�%���i�+D��1�����Bꍺ#�V�h��&�� �@�)O8n�ˉU�C�*l@�ؔ����v��8��E-�^�+�}u���z�B�
1R}���qs���~.2 ��h�L(���6���s�׃`��`���U��I�E"��>C��}y:誽��-�l}��.�r���`6��2�d�k{�8l��F��\�ěE������f+Q�X�{/;���3�ؐ�W@�T��s���ѡ�W±Fח%Ah�� �M����ځC���l��m$�	�� ya��08���|E�5�,�K:]�X�ZǛU��}�َs�Zꕎ�i�|��Ԋ3����S���w�\�H����<�����}���,c]��W{e �E.'8���"s>�Q%o�����zV��IH���[:.}���yug$��e�zF+����>�u��3c�8��ոz�z~4&7vVB�`�Z���`�l����<��5��K�z��@0Ce�.��.�%���Kم�&Q��j@������K����-�\��
� a�v�h�>t��t�\Aږ������z�.NH&�Ӯp�����{?�G?_�~"�/�-�C�>��IUʳ�����%Q����I1����fhB���H�0p
>_Q���h���{2�R�	�#��zfqri����E�8 .��"U��x�\K�9���@����֞)�߇��24I�d��+��s	O��O$������x�D,���V�ڦm �fy�(����XS�9����������l����oz�c�7��AX����Ž[��8���By?Tϕg�\SX#.��4���Хa���z��]7�9ST�e�>3�� (����	Eي���@�קE�ݽ_�U+ɳ�ĸ��� S�f>M{�Ū�ʧ��f��H��wɞ���֫�?�Zd���b����u<���%�.Įv.|��I��Ǐ��$E&:�H�H� sk�x��ΚO���lZM1:���F.@o���X��^@r����t���R�p��8��ʃu�������	�%�\e+Re�H��%�MWxq�' Kgdt�����ᑌNdK�q^/1��nw�B�8"x�tRk�!����:p�9A�.�A����R�,"�M��6gR�,�6���U-�w=1I-�L̕]�턁�g\�\b�������#I�Ʒ�mE�����3���T�胞al��|�`/ hu±�\����f��%������3V��ݑ��<?��P�+e.O˜���X����{�
��<��th���8����kg7N��Hn�Cys�����s=�� .Y4��qũ��Dҍ�S�N,�F"��k洮�Kk"���i��u������:���.��+9}a,黯���}y�<���-��V}Vz������+L][3�pVŅP�;�~��٩�_���T��!���L��,�xs8�ON�ror*O�0z("��u���;�����t��J=f^�#����P������P���~�L���.�׆]��p[^��sɤXZoD���&:�h�ԛ��Ft��$7�߮��g>�# {��om��o���#jYUfT������Ҥ���jF��,��}�wM��v ��cT�h��X%�n��H�{�p�O4��ޢ^�Y.iDЙ�F<�M%��\�0|~��q	7�v) $�g�&g�F9��rj��X7��`$s���R���
Z���&��߭��"E������Rvظ4'�+8�<g7;׎{yi��j��E� ����` �(Xs��@ܧ�C�h�ׇ���OX��up�Q�����#�]b4�yĠ��w�Ϯ�A���	]��}�9�j��D谓�����;������cZ�]�ĵ�c̢��#��H���%J��S�6���65=-���1���};�����mX�n���Ѳ4�1�ZCFa�
��Y�<�LM똑C$\��M�8`
��Vq#Q^�Ir-?XP��k���ߙ�6�Yp�߃ y�g�����E�.d��?�[W�I��ء@��2����Tg	"�=����ĸT�/��Y�9C ��J}M4���A%�or�s�Cg���֯�<��;A��#�?��ل�������#,*�������򫂼pا�c�/��k��D/�U�
�܂F:���@�n��/ޕ��	+���_N��S�?�qS��+PnB�Ǌ�EU����P���� ��ڧ}uj������,L��#V�����QA���rs��e�H���� `���{��0goe�dc��Ƌ|�y��+׫�����@��Y���6�޴��UE�_|[���<��������WSL���90C��o�Jz��ￃ�����+;�����/l6=�RTO�8�x��ݨ+�̏�j0I�1��5Pp
�Vƭ���m��r�s�ix0��t�+�e"{I(/v����/�)x�E������ԻA��>@�󴦦�nR �\m�}Ky ����"��j���0S�����������,n��Fo��R��b)S�4����3BT㞰�kI��4�\K���"�w� �&�x���s� ͣ���L�p��-� m�6�f�i��,
i��yCc���s�k�?����ݯ��|9L��_J4y`�֌��9��jN���搴��u0�Gw�
7��y�G�����B��8��&�߼\E�F�Hct�SRm�A۩i�Gk��ְ��ƾ�c窱�x�̕�7�E�fƍ�b׶�27~OxP��7z�j{��<{���j���| B+���K��E3"�B�xM����:�[�Du��AP�g�\�E5>m��Ȼ�,�Ύ6�`�a��
BJ�%�
��� [�9.\>/�E��۪QM�|��IGφ[G��>ԞS��38D���xO.�Pk�ݠ����F�gH�\�ň��X��G}���w0��&/z�Vu���������p:׭5W�2!zt<t�c֬��_>`Rg%�Ǿ(ʙ�e���18�
�"W'aaݡ,�C0@��/
i=���] y)��[W�w�2n�8��ų��k?�zW�)�;(5+�%q���|��u��o�S��k]N�baPИw5 ij�l�ӡ��A/�]g}�h�"�;3�`��dH��+�V�</���5�@E�e��|&��K}<w˜NEX�)��
���>c�i� �2�0����T��Vg�x�����-O�y���׍�0)�L���l"��B'�c*l�'2���|z,?��%C�c���Ŧ���'Ƞ] �E���lgM/<�MHZK8���B��<�̡�,��*T����P��M0�	��`$�u{��ž�����Y�` :N35\���`ӣA�Qvd�.���*�g�-��PFz_o��e_'��.�!#�Th�0� i�3��.�hz5V���%�^�d���& -q��K����*s����MX�_��¼?�,b-W�(����C�-}:<� �N�шU�hVr9�
%��cV���0u���X#&*+��H�l܇[~v�����՘m)�?�>��z�)��
�z�zc\'j[[�m�Sc�a�=���F��l������<��)Oȍ��X�s�.V:^��KĜS��K�T^l�u`��kY�1݄�*1�zQ��M~)�a�sd}8�3�8��@���a�Y��{LW���Cc4�`Ӣ.؏�P��y0�+������; ��ؾ�l)t1Ūx}e[' 5�#T�*��!��q�700�.R[p^X�mQ��]��qS��@`\{"3B���\5�$�a
J�`\�b�.���E)PП�`訓�$dM;:s]�����.�Tm_�����:S��+�B"��Ve��a��@��sj�~�!U`�vN��#���R�]&�.�Ut����7	���P�!�LQ�&{M� ��������l=Yю�K耝�U(E����B��A\���_�b�56"�+�=�݇�=]#��~�*|���պւ>�mi�t�g�C8�5��ƅC���Q��J�#lms�S�*0�Z����`����VU1���S���Mt^��I��0=�;�(������K������@^�YS�w��$	���MNe�g�Jm�@���.��p�+ݿ]�����-��JYL��5 ��BH�pq݌�q�g� 3e}�m�yJ@ΐF]F�4�w�ژ8���<�ReX�t�!c֝��'V�!H�&�ȗcr}��Y�{f}�U�گ���
rl�������;���S8�հ�8mC`�������	�6���B�J�H ^;V��8b� _�ψ�7��V7K�Py�|`�7E���O)��T��#)�P���> C�!��!ǡU1���bU7���Kn�Ɗh׺j�\1z����`3!U5̋]�Ǌ�y��m롛޾+���02sLT��54�fqf^���P����&Կ#�ZAE��\���B��FE
��~}sciU.buO,h�������(�?�����N�����CAm"������u ;�!PJ>�I��X"�s�cI���-D�o��)C�Mh�'\o�L|�ӓ����e]j��w���	
.7��zq�q�Cn<�=K��~�e*��������a ��C����ҙ`�76xtӶSU]�#�>y�D�Uos>�KW�-= ��t'�ܤ���}�;���9�ὕ�p\zknMsG.��ܜ���0��SR[�W���F٢)���*服q�g>�lzS��>͂>	un` `�u����S͡�$�*��n�V�G�^�Hg��^tq��.X4�q���e�P!"w��C13����m!d���z����B�?u�t��ˈCm�;#SJ5�g9�����T8�Q	�|>A�@�l��\�n`WM�W�� O,�M�)-V+��)(����@�@  �Θ!x���S�`�O���>�eh+
F�ح��^���E�qyN���IJ���HK	�=��Xk_7�a6a�."�Um�}x��C@u�-���5�ܫ�����v ���R7���Y0��du���_� E�����i2�҃pݘ�Y��(TxK��<���讲�W�h���$�3ك�� i���*�����&���Wi�*�5�n܋�t&b��R����+�,%ɜ�QIB�˄�� �1�6�V,Tm�46gX۞��C�ƫ�wN�?3����5M��~�:�x:Lu!��y���Mi.7.g��{k��-��O����Z�Ģ���t:���+�L^U�o0_1���a��䘷/]¦�+��T�r�,/t����q��IAtɧp0`�z�ꉌ�ؠ���TrW��.�X�F����y5Hi��5�� �Ba�D�'g��LQ����(�J'0cy#��'?�g��gB������Զ�)��/�3f�#1�RLTӆ�s���9���3`�����t{(�@5-<Ǐ�qA9�$�*�(�a"��H]P�1\]ı�Z	S�ƣ���⚪���E.zx�41@����|�Z&N�~��܉���7cRȣ��D�'�c���kԭ(Gl��ac���;�P=Wc��"�Ԍ
��3*���s�%�I�/�ֺΘ�6����a����^.��xy��X���0��vFM֓$�T������*���֔Xcuve�0�\�/m��t��m~�����Q�ڭ������N�������yW�sX3e;y�'m�7d$�����-�Ǡ3�҅��"C�W~�e��$����u�����ƥ��� V�m�5sEo�0l�y�(q�?,��7���7���E/e8y�h�	��P����S��� e9�!&�
Vt��Ř1w�dsf�L���k"������b��զ|N���K[��ډ:[3�SΡ������MK"�#�����}���C���N�B�g,��?���W�jK��CD+��
l���x=��;N�Tr�W�Y]{B�F'�s�^|���`�yYS���%�;#��<g��^�����g����3�T���S_�fb�t�7E��R��-g����~�υ�
�E�Q{��\_5mF+!Cȹ�@}�!!9�خ�޼Z<Ơu�y�t|�r5ҡQ)���t|���U4��eEoW-������d��ވ�-X�ڙS�K��
��]� Q)H�
rR�=\�q,�B��@o'�N��1^|^i���U��WT	y$`���b]�If� #��{f9yI�&Q���ja�	�UR�Z��x�j�s8 ����@��f���`_�����;�=#�F���i�Ĵ�)'�Ħב���On��B�.�����x>�bV��M�k�E�B� �j΢� XW��Z�M�C3R��U뾺�
�R�K+����g�����wB��djj�k�jV��G�/������d�W|S�x��t�[C)u͕	z�FM� �*��,a�����yfչ�i|^���^/�yټ�ܷ������E�I_�U��f���.
�#$���Q�����Ep7�V�.=�֧�����f���^[� h0�E����N�ξ��I�-�F��/�i,7��A�(kK;$�y���t���.jK���,���j��m�mp�.{����\��mr�+Rr_AMIT�ZDߡD0�l��Z�@�*M-�������C��UW][dr8���>$��^����ʀ Ҩ�ǌk�Z`Lӣ�s�V��=P8INumN+�}�Gc�r����5�(|i�z�&���j>��aN�u$��Kjz�֮HF\ڝ΍�����s�����tU7ZO��q�ʑ<;5�$Pm�$���j�k��72$����M�Bj &
 "�8��ܿ�1i��;Y `C�"A'#wg��������"�(pݗ�k����DrP�Ϸa�.zI��4r�ѱ)yP� SRe�mY�{U{�Ҡ�*U�h.�`]�����ϙ�od��	^m���c�!�C[�����9�=x��+>88h�R�X��Y�Й�W���HF�HV����N<�n �ɩ��:�94w���%��b_ܗ��۲��%��zJ(�7��0W��9#�^�H���h����� �����yx �Ib<�qx�)��⃉��C�$9B�3�\;lKU����Z���j��'+��Y�������%��*A����֮�^�Q�^[Y�&t!�|U:�tLNL�Ț��3��g�~�8�h��ߵZA�$���X���2�q�gO�D��Q����I��&��VP�,K��a�E_9�]�s��ߟ4�z�#	m�X��k��T�㢇8 ��/��P�+Z}��ل�u���U�1fb��YnQm�!�&����X>�M������#hm�ʭK�{>Vz��D��O������&�W[�U���6e�͏!X
c�b��V�ީ������%��!��g�gޅ\⥎g��
�kX.*�1���y�~����������V$.rip���z�کQ�m��]�"�����w$A%���ܳ���c��tz]~&��Ԃ���؁�SvU�>b��K�G`�^±�4E��+]�0u�$x���� �1dU��_��$�SqԵ0ǡ�O�-�
�J�mQ>Ղ R�%͍�ݰa����޴
�0o��A1$� �PMidU��
�����-�h�����g8�1�X� ��E��-Kc����v}>�Ɂ+�}Ud�Li����
:�H���3�)h�RX�M���k�8X��N���4r�XL�`3��K#�W��b<��@|"+p��B�Z%��@N�"�l=�7+�k���v��Fx��ϔ��EW�9�FFr:]���QǺ^L��`&X38#��)@��������tM�ø��ul\��q�u�\�P�"�I����q&�E -V���7ZUEg�SUB�6�]�q�ڧ�̦����������V��_��g;����Iqy�& ��
.ӵ,}��C+�ǳ22�\�9�w�T����!�s;�m�,,�"����wؗ���,�>��e�C��K	�3�^�Č]�M����ڒ��Wd;[���M�ˑ�U.4TX�s�Rf.�}Y�0$
!��1Z9�J]�w�Q|�v�pEk&Dv��K}���	���?D������*
)'!��n\_�r�$�|_�w�7�j��kW�`�Ov ��"H� |S,�{[�٤�i���\�{6ܿ�X�"}��WT��.L�����Z���JIFEJ�ٗ��1�R+�g9�KG�z}��,>9]H9p=9��j�sc�Y��Th\��m��N�tO�pK�����d�-���u���+�1���Q��W��y[�~
j9icedxS�`k [o�t��LO���W��'���S\wg�����9�mx���$��,��U�T��H�w=�l��z#@C ����]f٢e0�v����a�\��ǥ�nvU���g/��1G]=��fƻL�րxmnq�ގ��Qi5��� ��	�^�X��i.'�:'��T?�	88�h�L�Y-���,\�T��*ӡ�Y(�@��z�0�6V�$#��J�vzr��7��o�bk<q"ۡ����Mｏ.��� g��G6>�fob/&��(���Z����1������VV�2U������,CC2��S!?ׂ��Z9=�ȥ��
z��4������U`^un� �C�gQls	���0��Ђ��Тّm:1	�58hk�V�:x-&���nl��f��=_�(��{F��Ru���%�|y-�,�M^�rp���ߕ翐)���P�4jatG��}s{�$[��6* �>�(c�VX&F�W�,���6����a��Sm	,��=猟��U��]��_M��M�ZK���.[y��@Dz/Rٸ�ue2��E��s�t��R��G2�g2&���J���0J�_6���h"��#��»�ł���(�T��bK����L��*���wO�et�S$��xxR:�����$,+�Jҭ�n�L����,���B�	Q�y�K�h¶�[W����. �Ǎ_z���nL�١�F�7��T�h����W��΀�8��&��P�46D<�[%��}�^Ҹ���T��B�+K}Xcrk�l��wY����G�隫)SC��4G��'3y�>�R<l�Cն����1�ޓ���C5u�&�j,�8qqC���k�Ł�k����'�N-�G@���!1��C�\�ƾ�yc�ȥ	7���W��%~���r /v��G�n�G�!��Y�-�/����!��2��$(����Y[.���=��]�fG\�[;�0D��w#V�fs�H�͙��M���#qڗ.*�S��.�*н�HA�^�_�ڍː2!�Y�XA1`C^<+���H�=�jO���e+=�w�,��N'p* 4q`�K��b����e��r'��|i�3K��-��z�t��p�s1q^����!�W.�,�Q��6엸B�����&�O�4�n�%8	wK�oɨ��{#��4=��y�k�Х�@M�~\��T"����et�ڶ��놏.��<���!p�Ddu�M����(n�����d��t�@+���{E�� q����|������
�N$�Wn��۲���T[�64GO�*��֧���p����!\s�sfqϑ�����
��=zĮ���KhF�K��x¢o��L[�J���)Pծ��W�|�m�Y��v|7�C�Zl��]����[�O�E+y���rp��'� �뵓�>s�V1Y����ǽ�H��I�R�M�6��+�kA^W�y\�rz|(�����pK ���Ϥ��w<Ԫb�Z�m�t�\R2Z(Bv,-〶%�!��4`�FrVT����=����fɗ���Y�Unp���h�1�
�klx���IUE��E��e�����<�J�Aͣ��ۗEn\��G갅�}G��!�ډA[u��u��ܕ�Ea��at��e( ��`��d��n1�Mk��m�U�9�ku�����Q�2���B�Ij�^�l��6o(���.�#q��Z��g�����N�E�.h+���@����D��qhQqZ��KW����j���u��wg��p�t�c���g2����C���Q��2�*1)�Ll��M<v#։8jq� �󅁐�  @D��������ҸB��4�_�J:r�����hl\I�Z�@�M�у}��Ƽ �
<
�Ɲ�"�p$P���L���GHE��Og䋡�_X[��zn��������_5�Ot����*_�gYaT�O�I���]O�9��] �'�.�����}�zt�,� ���n��C����2RJub3^�D�ޚzЭ�R]tP���Tl�yjg"��{}�9��#����v�B�8 ���I�m�~^�������}e�@H_����(�����/�L��,ֳLiA:R�҉����ig�;"��?�԰~u70��+��N��;��'�J��M��a�@NR�C��PV�	�%DU����@����]�*7��d���uQ<�E�}����D_�q\�ٯ^O
�n�=��[��ٹ�`n���!��� 'г0]9�rë�zdK��-ʦ� ��� t�H���2q�����OXe��1E[Yj�	GY��B8RA�s@�P��ͱ3�<|f�8ʵk�����݇\�Q��Z�|J՜ev�⸦�IK�Ulh}ܥW��ڠ��=��xԅ��O���W�����<�IG=����Y-����_ك�凞_o-!�OA)\�w�b�~U���(؀L
<J>,TiY�.ۨ)�VV��HN��AM�O}T�~J� q��D�^p��x��Z��3WYH<2�c�)r�ؐ*��z=Q��V��"�ڕ�܅֌�R+he��#���h�4��JJ/[r6�1�@7[0?bD+J$�:F��[��ƽri,/:^4������	�P��$�e!��B���$;�QwKw67q��4��x0�AWyE�ɞ���}�`��ik��=����d$/��:kW2�>�ulR��ڒ�k���Χ��F������K+K�*xcn���*ɂ�Q�����u��w���;��r�ynk>r*���U�?n���|�'���*������Tz�^���15�*z�i��UV9v�7*S^���;�(�(����ۀW��1�ө�a��\D�PR�7����v.�����u�;�b[�5�
Mƪe�P":}�c�(r���ĕ��Ḇ�ee�K��v0�Y��c���ܒlyl����COG ��,�ؑ�U�t4;!��@�-A�-L�K��]u�5�l`;�W��c�-��0)�~�*��IP����1�=�_=�o�ݗ''S��q�:jumn�پ�~�7K�O&:!���a�:#��*F��K��FG��6#���[�c��Z\��޺%�p,��=%f��wR�K��?���s�޷%~,J�
���Z/]�:�:��K]��x�t�BH�ԟ!Z��@¥���'ؕl�dE��XY�ך37�v6�I�EM������wz���[�J8~8���R�:8�a�y�:��:3�>�v�8��!��z�[�V3?���nUm��`�v�/��[r4Y����y9Ե�6�t����ɩ�t��&Şu���\o�;�S�ؑ9�*(̀�M䪭�j����(��=��[������#H�>��Fq\뙓J���d޻-XTP� �z�������|WĀ�mz��o�@��F}����ZCOm=l)�J�o�N!<{9 v�ڳ"�,"CV՘LV�
f�˖Z2�k�V�. g �7���i��y���,�׻X�o����ì�}6�c�܂	<c��� TmI��].�-JZ�=���NG��reg�X��#�1�[���G#T__t5 �+�;�X�DG=$�!�i�U�e�> <邞o�&V��ώ)F����٘ ����Q�hb���E9Ya
Osbh|6�P��8���NH�YQY9��J Z�U��f�7��F�$�~�W�[�� '�J�']����S]d裈�B:��Y|>W�X�QM�B�~\��"[��yp�5�^e�,�3�V����S
'Q�;�w�|�kk�r�I�Y�F��N��d-t�������.ִ�� �����E��x#�@@oD�3���*��}5�76ҵB)P��� �@Z��Z	a�Q#���'ӊy`��	̿h :H޽aK�6W��t!'�����f����H���C�U�����:�+E�*AĂ��}E'V�A�.�<ׯ�}�/,L �(���� ��kDCW�f��5��`��ՁT�uu{����v���U\�.D�'�V�:lz ��#��<6�ەK��4ҙ�#1�:ū��ϋ
�|���fĎ�;0��KxZ�;_S�
j8]+x�F8�C�Q�{1K��ْ�ζ� x8�v�%�ߖro�ܪ��)�s�2[G�\,�U���X�B�p�T�ʐ�l��]p.�P�5��|$��l:����թ��h��AJ�}J�@���N�� =�A�����8��U;�ӳa�W�#���wNyy��(0���P�>��]U����θ/�>7A�dp�+�F^���"�������w)��)��B+@J(�3�P�O�ի]%i��sTѬ>�Q���:L�N�p�WG�1l3��Yz_�=���K�z��jG+;��c���*������.�:�MM��c��9����['1�)p��	R*(FLtn!ҟG���m�4�䆭��L���!sC�a݇�XI1��E�g_�*�ȸ��փ���xNS.	[/�]�r�"�>J�3(eK@+�نn�j8��I�����7���pT�S2C�h2�5
Z`y��X�d���6OX7�	�G�m�c���Q*�ڒ(U��v�2Ս=ߎ���C�$�����u�Z%<��3<t�2�z�c����Ri�c����.�"�0�#h�+:�SuuhDF�N�:J���5�\�p[�V�(]��^a�����)�O� 0��,#K-��En-�0��ͥU��u�u�C!E�8��D-���ha��z��� !|T"⹶�cWDD���u��7
���3<�3�%I�S���;��DG _��e\ѡX�1�eT�v4D�Ol�N��m_�h�����rkNBQ�v!3�'������*w|�d�DԖ��8T)���B1�
i4�&��4��t�1)-Z ~!����uL,��t�<��ɱ�D����S!ЌXU?��C�i4�g�d� ��"F>P��aD�&F:\�\�o����5�s�����{�8c�%�=�z029�Qb�VU��
Y�NI���\�'��3
/<�k����q�\Z���yq/����T�"���N,�h%������ԮX�W)����#�7�4+�c�`�6��w�k�@,�Y� �c*3b:���=�69�D�r�[�;r�N;�:����l�W_��wߕ�~$�Չ޻i>�u���49�j� N�]Z���L��4� ^�t�U�����tُ-��o��s:�Hi��	h��,�ʰH�������S�m0�xo[� �Y*7r)Y�d��4��Xe>��.�������>8��EX׋SH͸z�Qq~�8��%���H^�sWN�����Xv`�ف�lժbg�PA�
@@�9���tibŁ��ߍ{��:�?�#����w{,H��L�B͹���n�c�^�1�Kt�0�2��}�s��ŵ��S��=��A3H��C�)�s�b����+g3��Ɣ@$?(�\��Q2�*�'�h8V�t�@�� 
�
(R ��>w�����ِZ��i[ ��	���NB�uU��P!z\�6
�����=g��(p�x#��e��e��t�Y�U��e�6c�)E+��m׬����:�����i��l� ��뵬���C؍��Lf1��#ġ��)�jCO���е>Y.X�p��>�����\�ӄ@�<.�)F�-)�cI�}��Jd�:�sؚ�_���9���F=>׼�ܺ�E)�R�����ET�����Љ	�E0>��J�9�S�f�:y�5⎻���!����E���a���U��Vm	a���HX�$��w)c�	$V�4�ۖj�]�����PJ�� O\F�#��F?\[BK*���*2���a���������H�/�n��
2.�]��ȃ0���0��h�6gd8�;�<��8�W_,[/�����o��.�۷oK��'R�Nu�w��j6�'�c,X�_1�,��3�6��-�Pߤ,���Jm�� lE)�Q ��!v��O�>���uQʠ�aH�q�n��C�(�N���.L�RT��C ё@=h4$'@�FW��ѳ]�I�z�,K�T���ZE�bָ*�T9W^[k���S�u0���f��@�`㲋�>0�v�1�Q'��lwui�!�ޕ�OZ���yP2��hUV�l�f�S.#&���վ��,.�s3�Kv<�\���"��?�P��{N����!��n5H��ήt��HӀ��lɭ�ߔ���猈�s]�ǔ�8(�(�R�w���Z��G���)Q ���v�n´:��=�i�%�M)��)�Aw����k�GjwK��9)��S�l\`K �Ї1���C����Ai��V�&�Nj� ��%�5��Ljs ��"�S�)z�/!��NT7�uE�G�w���(�QG:C��Xb���J�ct�gYHP��t0��F{W��%"� ��rMF��!���%&��ӇR�,�)-6A_a��!JF]�7d+�E�����������:�����d
Z@�#��;�2?<V�ܓ��ʠE�� S�"�I�JY��S�ywk[��m��<��$T' xA>}�P6/S�(t-�չ�u�*�Ś�C��e�֯��@=�S�iW���rj~�XQ�5a�5@�[lO��y�Pbl`Ǘ˥,��{N�m�{<陈7����s�H�r������Y����<�/dx0,�����\�C-�ɂ�k+	Gm!ֲ�@ >�vtd� r�.F��@�8*���`D��ˮ�sŷ��̦:�C�u��@�ڬ4�6��nd�@�@��:�2au�k#Reٙ��<�X�ҵ1�M�a#��<!��R(&^&�|�4��ŅU�!��τ�]��P!��ӛ���I��^�ڥi ��>gGe�H2����Ɓ���!k�+��Հ-��dgF[��� �G�t
[�E�%�������"��� p)��{���!w|r��eXR������Чi��,_�d����=]0�?��&������ڨ�)*�tcuK�������Tⴌ�9�ʸ�mq^���P�\��NXͷS�ƚ,%��-o}���/�#c��!x��uU�z��0<��Q�o�U�L���P�:�aJO��X�v �z�
�O��/�&��g�{2F��7^���/%�N��$�'�:����h���N��X?��vdV.)����9=YbH�/ƍ�@[X�ZX5�5��1�"q,�g^o�t5�j�f��͊���� ?���N�h1�8l��l}��ͼ&n�yAx�T3@�vܓ�^*��
�=��3I�C�8q��#23�",��tΒ-��1Ӕ(D*��ԗ��O S,t�N�&F��� ���j��CE4iR
�����!�s��D�\v��.י<<8�|ԗ�J���emU�=0Ý��}��DzEʔx�0���|D�;����	�����s��8��:�=�ϴ,��[:mKo�'��g17��@f����ZU|{�+ꙮ&o�� �W�{��Q�*�'vI'�v!.���<E�`{X��e� ����j;�Q�ALh�aܣ�#�.�S�6f���`(�����ń���Bm�{K�fqgG
u���&g�J�N�v�hW��:�:�'GG�<��C]cIs2Z��f�7�_�=��K<�ȉ��,<�UR�ޞ:�
×_�L��T�X�c�#�	�2��@�Z�-[Z�<������:*�a��8�P��L��ҳ�@�O$�;}JǼ��m+<a�$��b[&u$�C���x��kR�_�U� vq$�P�oo�v���|Ѽl��~yO>��|�@
�����kDDu]�E"��ا)�#Dy-��FI�/�H׵�40-\#��X0 (s
��=ѯ>q]Yp���� �{_�yۜ�[Ũ�!��hҐ/dv�T@/��zB���dN�8�}�{��OH5�(����=�
�Y���L�����J`5��
x.ᐞ?U��
�+�f�Y]�����0��Ahƹ��2�کG��c�5�{a®��/�j=u��q�4�x;m� ��A��r!;S���0�@�84V�E�nQ���f�}�p�p�ӹE6j�S=*<]���r�L��W^���C]�K�U��=�$,���ԅ�$�pkLɍ8���X��� �0�8�Y����&�{�e����҉��"���~�n��""���7���؄v���]}��#��j�{O�d��+H��Օ�Xt��z�u�Ѐ���F��A`��+0�+������P����Q�H���y�~�K�3���ގ���Q/��c�K�%Hw�RR�gX)H�X���j#"�5��m����vm��x!���K��$_���壟�P�����v��0��Ģ!�3(U �����׃�^M)���Ͳ@準���|�j�ˇ���O�U\����]T���d'�Y�*�0g �i�e�gX@�:x0��!�pû��W0�ֶ���c/p)$����j�;�nc� �0�u^QG�U�B^����ܢ��� ��X��2��T��ړhw�=�כ��*���n�(P0����C�KJFu#���5�.��W��z�߻%G$x"��ݓb{W�ޖ��S9)2�~�s���}���_����~&��'R(h�Q�)CZv���'׳�?��Ll�Ѹ�J���5Z��%�D�H����P|���蝻��xy�& ����9��
�7�a˨U�S�
s��\A�i�⬝>�@�5-�n��ՑdoK"����}�ת�oV���P�3�s5ڕ�ޖ���\�d!YTڹ�s=�q��;�{W�:g�L���	�P���saБ���MԞ��V��Rqk��Ց*�n'
�iQ{ܾ-���r�� ~!�Sp��:FTewwe�;2އ[���c)'S'{
x��� �'|����]�����aM.z��Bz>�[�����<3�쩳8<�yGA"ׁ�8W��2]]�a��R���x̬ӳ88�P��:w���.9����S�`�� �������u�
�Ȕ�jl^l�j�v(�@�T2���/,Lb=��k��ս���En:c��-s�송Yv�qk���!�N!��C��j���_|�?�{aem`���ղICa}�)�R8��(l �&oc�/��<O�ۘ����{a�>��EqJ�ӛ��|t:��JS�.����6��ڲ� �Q%i�Bz�,�_�4�T:_�z6#%E�<�T<�},�)�!iQ���W��`P�_ؗ��		���$��R]+"�5DJ��0�A8�s��&�O�o����K�=Ku�b	U�cV������I뿍�aD�Q?.C��9�ż���� c�~�b)̏e�r����l�K~�j����om���C��F6E��PA�j���������cJ�Xw�5VG�L�������dR|�W�Vg�4�7��_�{��$e��qp{��׏��|4Y��0#b�� \ܴ�L����F
j�ޖ`{� ��-�� �h��4bJ�Ǯb_i�@ 3���4W`�m������!�HZ����P��-{�{QNer8ױ��,ޓ=5��S|q,/��y���ޮ~��Ux�Tm���;R5��Έ-�V�W�rd�55��{w$H{4�K�-�s��eH[Wf8J�0�Ў��(�xK�v��v�����z�6��%)Q"�z�x�c�M��h�h8?��}l�C�A�pǉg4��h�DJ⦞s?R��V23E~��ν��sK��K}���F��E�y�Lp}���\��ئ���Nz᫸i�9S#d���SmӐ�_�9�'ʑm�*��ٗ���NL�V�8ü���c�K�L�u����'�&L � U��)�����W��-��쎜1BD M���/u� ��p
�� �\b������5&im%�g+���dTe��\��� �U �& PA8õ|�}Q���g�plTs�t*����,�	�.4�p7S ��٩����gS�5[ꉩzL���ͅ�Aa�9�q��QJ^F�v�E!	vs��0ܔ�mt�~=������x`���̣T�粲� ��r�j99px���t�y2��h�vI�2:Xg�b���|6�v�-���.�w,4�w@�e/�	΀��D?��	>��$_?�E2��OT׳����^� ���s��|,�JM,�A�T�T9zLn������~jZ��S�4o;��\���G2;?�x�yX*�9��r��]8�@'Q��z[���3���42�Y�2<ɓ�
��}��]���h*Z
��� =���lb?��ŵ� �5@hE9j�f�X���Gѭ�<VRQ�H�R8����6<yb�m�=Ξ� �eY�QV�钒���I�M�0�ږ]1	���������V)�<U��,UZ���NW9��ڴ��3���03-R����1�Fp�jf��t6�4���
e������n�Վ���]��i���-��0Q�S���\�"X�����in��}_S{�އ��(��<�l�I��n����B*��ݭ��h�e�gL�H�憩��e�2l6�$پ�i �6�� R;��x�GvR�d���0 Uz�E~��j������?��ѷ+�NL̔CV6���i|��ӭ��ɟY�\���
�:F�][����*~������â_�x�=�"� h���vB�9~ *���)s����R��9��[����<�1U@S����H�(O`��0x�]<��ʣ�Wn���2/ ���f60�O?�L.p��G�����꼰����r3���1�����6f��~�Va�v�x����e��-�˴��|1�_�9��q$V�ɕFW�'sM�j�b�����5�hǘ�Bm35�Ɯ�"sX���d$���UI2�O��L�)��.���� �	��ta�y�����8�y0���
�G
�k���{�tes:��` ��o��s�=�B���`�)���@܊k"��y�8�u}q$�X+�R���q���q�	����-!�;��[�l��n��e�T�����򥜮#��x����h�bC���MApF�iKz�\�2]���ّܻ�wo�^ȓ3�ˎ�1`�z�F,��0��珥��+��X#�jy�ve�^=��l�c��ڄi*�߃��r�mje��4Q @X �º)&����]=�˕]%J����X�/ڨ�b.�q$�{@>�_��%���I�iG���mc_,e@-U\�[C7�i
.#� S�M^���y^�0�H�y�9韞�n��.A^�X�<ƽ{˞\�Iw@c��� ;p��á$K��0v#�/��>�F�u�/�u�:תG���P����g�m���'}��w����ͷ%�>&S���$�@�f�B{����L� ���Ʒ�!{�
��G��D�Q���L� ����%��w��~*>;b�0~g��Y�"[��L#��<��NH�Uȉ�0Vo�V�����-q�jK��%_�Z��کEǇ �u��ئ"��2��X�F�Z�����-:��ߋց*FRPw8>�"T���:؆��:�E�lO:�� �xHgx�Ƣ��Dǋ�@4�E>��x����܈f�#��g�?f��&ݬ>&�.5M�ط���t�\8��ZGm,�����"�#�����r���R���6�<��o�[i�fZ���^��"l�����gU=ݘY�̌�Ik�'*0a��BL`�=��Ya5��B�\:S�lX:@�$���G��U�
.�Yf�X��&3�.K��|ۀ���2M�8��%ILK��fsX�p��a�K�횉$1�G�VA�ci�j &�����}�V71[;����d9L�|-G�<��B�Eլ*= ����9�f�,�!�v��ް��<X0j�'�b�j4��\#U�E �?Q�#�j���oTOoA��͢h�e�A��� �Ӫ,��9%){��<iW�b6��:٫������y�!���|��'�y�>1 ��*s��u͒W���s�:�Fu#V�
�� ֮���<�R�H�h�cҿf��K�&�GyB"�Rn?�'G v�?���rYh�T�IJ����q�=���>�)$����h:��:'�~%�VMZ�I���3�./��r5R���S:)S�����I�ni�aSDPeD����:X��a�j\,2�^"��I��e]NΟh��G�L�Nd[������Is���iwt��g���e�E��A�JJD4���r�3�:%��(F3�O��7媏=n�n+5�����WF��#�a9R��  ^�P��\;KY`�)3ñP�& &jF�#��0oss�Oe
{���vdr2�� ��1}��l���T]32 �)���s	�r���x}a�Lp�1��j�r�2�N�R�� ?�����`9����W�޺%ؠ	�ѣ����Ӟ��f�qM��0Z\E4��q�s���r݆y(M�����}IV�#�03
��`=�Qۗ�xG�o�g��:ݪ�Q[�P��z�/�(/A	Jw���)y���P!�q(iI���_'�n%Q�Tg��d�`��8�҉<;�Z~������-�bOx>O���t.K�q8�1�5E�YϔX^�����mS�r���L�@���=�/K�_<+,�\X�\�yU޹{M�ә���%�������m����%]����}����s�\���������GL�G� @cj�/�0�ˏ�ߕ�r��u9�$��oE��\�x�ݿ�NNqE~G����b_� �T��e�Ksk�sj��t���ܿ�{���c<w���2<��f�	�%��(]s߁/�o���F��5)�W�_�s7국^��P��� h_�RV����w��!��W���ϱ�EؓU�=��ȕ�ܴq���ҨKh�68 ����h��)8O^lz�$ ���9�    IEND�B`�PK   �X�XW���Y�   /   images/a615f73c-88fd-4a5c-a08d-6962f48a0070.png��y\S��>����(M�2�P��@��5B(ȠTQ@��AfK�(S�*aP�a1Ȍ��H� "2q C�����{�����ǫ�}�Y{�g=�Y���Km,7|��+�6������bؗ�uR�'�$�¿��������'bݯ4��K���R0L��-���a{�C��#T{�SԐ�'����3�����'��=3&[1�;�gҿ��G�¯����V��Z���?D�&�^�i)��S��]ڸY�0u����~�?��c|{"��z��ʇ'�5)�ʂ���o�7��p��N}��ƞ��L�/z����j_c�����U���O�;_�.T��p����(�������C�=,l>�&\�\��ѳfa�T��pW���ao���ܩ�wĕI��G�`W����������!��x����]�d~L����Ҟd%��ѓ�T��^ZI����>�����i����]�	d;[ZZFWR�5�lt=��}t{O_9�߈��>�±|��T�G]��h�w���1+�%���'��
���Q��ߴ��tz�T�G�F׿� [j����wZ'�8��ĉ��ྷ]*h�������G�<��nr��Kn�J�#�~K�q����h5�KՈ:����%7d�����Z��$�g��h�?�>y�d9����q��.�����RRE	��}k��C�MMM\'��>�U��
d�ytq��S�J��m7��s����+���=�=�8p����z ^��!��u�3tt�>�9Nܾ};J��*@�c�'�r*�������u�M��׮]�}F���0F#r�#�������m5�^ҫ�_r3��3h�f�mN�x�����[�����GQ��x�1C'�ACm���*����ue����Ʉ%v�T����w��yZ?��6�W��e�� **+/=���Tc���(6�RSޢ�Ydh�K;�hS#���m&�0@�޽���*%�����)�T�[�u����ˢi�C���3�˟����tʟ��1�Vç�#f6�ۅ��*���S�b��OB04��s{Eд��"��gu��S�Y����o?`c��J���M�_�����gv�<?ک2��?��_ll��i���+a�.����KOPT�%���m�h�6��z������s��b��F��6d[6���"�������o�eJ�.]
�H_�/x@��)!�����\�_���gϞ�h����	SOJJ�la5�32����ND�&n�{�EC����lٲ�۔��F\ǥ6���p��w�'�w��{��6�!�2H���nZ�)10f�ӹ���3����6����Wed�)ง*E2<�r2"b�&�Ґ���FQ�g֜=�&fc��������R�5�{y}K��(�9� �?�Hw���ٶ�8�&^�qc>�&�-^��W��ߤ�����D�W����(<od�QĜ��O�f�����~�"�guƒ$#Ng� ��:I��c_XfCMk��@�%����;b�Ƥ^�{ws_���P���,%��{���M���~]3��p�Z���[ �F�F_��:�(�-����|���z�l��-�Gmp��3�dk��顡!op>6\���؊��^u�#��z�n������{^466�0R������΅��t�F��m�o3m0X<hŏ�]�{\z��r�3�HC��)#�<�2��i�*,�5��P=Rv�%N5jL��W�1I��<Gr��!^L[@T ����rjMlx2��1U\v�OS�-�����B!����8&��l�(L{ݨ���Ą��r{���t��ɂʇ �w�õ7��Y�7�%�|�OF�ǝ����k=�l{��2'f8D/��Z�@YP���������A���|;+ՍD�'Ʂ�c��YXXHY�Q7���^�v�0�!�e3n�Z�>@��'=��i~��	�1\�[�R��Uv"�3M���}칳`h�[e��|ox�ޮce�]��w�ksW]��^	�q��������i]�Lbip?raFU[�×��~~H�Y�|��arg�l��-ζ���Q9Pc�[�mrYN�]�*��3u#���P��&�������dG���y)�$��^�C�{P��C��&�&q9��3>����!E���h��:���Q�U6�Z�(g>��_T%��HKK���[]�|�9^Z����]�`���h�Eb�d�B��֖ԯb���h��4��t�݉=��2:������ؚ����oq+����q$w�P.��Q�e��-d|����V�Z1�&Q wA�oW�5~���w|�Cv?i�x�_�+�*~-��^c�0k u�[~���ȓ�*8:�6�k�"#P���̞+õwq�Vq��[������a��xQ�̛ ȥ˴����UW�-f[XZr]+=�����g��ۧ�H�S���(��*=��!G=3�H�w�+6W��hT�)ꪨO�t+Bh��oi�}e����ƠNoO?����-̐@����,%k����a>>#?3�9�h�)Q��xK�e��Rc�7�߽{�A�_�+�[��'
JT���,�-��߶����z��H��%���+���=�d����f�ĭUW䏘B!��3:�]���(�p�u�ۻ�PqE�Ycgŗ?�|��d}Sӥ��d����4[����y6�ŷ�n����U/I�zո��̌�d���r���
�����I��&��R,�8�?Bdj0VTp�bƌ^h&+ϔ*���ە�ya����ϠCV��8Y�(7~҇��9Ð�F+�����]����R�uȮ8�����*1-��W�BH0�l�"?�$B
$���f�`!n.F�Wտ�^uc��h�Ad�˹��5%ԧ�vW���8�O���
�p�������ga��x��=����� m\��� M��?�����a~�L��!
�Fa��������*������)�@���12\R���f�*��I�*R�3o���䠓$j�Ĳ�X�AYK�~��K���x��n�?M��\�����Ye���䦁Z�"Z�S��6i)��M�.��T�ז�x�_�G��ϊ���`�*�dk����@ �i�nb�c6E?�|~ӓ'Y���g(�ڶ!2`�'��\�̗c�_���"#P�.&�9�G�_�֫!
t_���� �h��.�Dx�!���w��K�v*O�DxW.܄[Rc�j�o���K `�OZ���9!:����nbKb��@��©Y�vkov=p�ZF�lN�l�I�����$P����&��(�aN(�\za'!%l�q���w��Ug)����ߐ!Æ�{{�w O�fQ���G�^�ov����X>p;/��'e��*n������R��`o�!��2����k]-��w}����묾ٰttC�wW��"�r,M�1���
zW�_�f�9���;��7��*�X��e����?�of2+!e�jF�֪�����>&nb6O&�f���ɺ���!t�����e��U�n��3�&��B箂����o���"���R���s{�_E��U�e�?�A�$�'Sq���f";̛�5�~���ձ�1)�wqM�LaѸ~5�K桡�Jp�'��vk/�](H&5�8h�>A�Nm�>�A ���&V>9��S���]v�t��6m�����`���� ����$�O?0�?I�,�㤀,{rg*J�;�5[eP=�_�w�?����O+����MO�>���t�.L�#y��Q�1�����S#Q��]f�i��Y�U_�C�L�u�"���}��%��V�}N~uyn���ށ,����E�UTڀ�	�3�kgHu%<)�;w��D1���x�-tXx	��65k�(�[p��U7���E�f��u9��	Tm5��'���Y�UQ�9�$�wS�Pd3��O;�Z��R)f&�w�=<�K�)ϿR@Ȩ���{z���֨��S�\L+��'��Ea�?��p�A���	x�T!�o�H�M�2��d9�o6�FL�Y=�b.�WX�r��Ǐ�E�����JY�c�-�f�ݓ����G�S��Y�1����|tϑCï
��K��gb<p�xt
{��x�����D���n�5"<s�k����d��Ϊ8�c��'�3-�C���Zɩ�Z��D�p#Cz)��=�w�{�GT�Y �a�֓�T�/O���"|��,�S'F�Hʚ|��v^��L&?.�hJԼeL�-]uf��LN��h��x��-��v+��V�o8��_�d������鋪NU�����㏡P'�L�ˎ$�<��f="QH٥��j#j�O��Pf�����:ɎKcI���]�왒�M|�h�j<񋭭en��L���{u��9�i����n��=���K��|��S�N%��Xz]�)�-rr֞%<������Ǹ�2��{3���YZy����~F�W��U6��=p�F���k��6\0P�� ��+����{n1��]���{� �^�eZ��z���a�"�.��P��������F�b��9e�
[[ۺݼ2�@���g�ف�R�֬���&�
s����u�/R8DR���Ĥ��LWO�]���ۿxO�e2啔ve>�y蚚3R�y���A�Eh=U� ��|K���_"�D7�ثm8ۊ������;�P2KZ^����R�E.��b�B&��v:��
��A�
�cqq�$ MM���)�LR1u2�G�kYw(&�=fP���B]9��֐:tp�
���[\�0���>mv�����CzqBnt�� B����3�!`G0��%�o�̺̕�y��sjq��҂�8^�^�N"�28&I��$�p<�ND^Z�0U��Wb�~ ^�T�r��966�a��o��í��ޮ����	;��Y� ���{�����d��"�Xw��a8�0Y{����_�xj�M^p��~C/T&_���$*����V���� ��N��ǳ�Y�=z����d�^��%{�Q>傦��e��/��4���k;}�3���;��Ͼvm6�6[�Y!�齲�0>а�!�\�V��`��>J]��%�=���ɾHa_ /3D<��
,qw��nw]�o��{���x�!���\�Uh:Q�b2��|J�������p�#�j'�Wu�FY�)����O Kj�cb(�� �nP��sm�qH&~ۋZ?]6���^//"��t5����FE�;��n���H�6��<��I�1�RZRrP<w������ߘU�n�p�g���}]'A=o��Ӄ|��k����n�'Ԗ�Y�]�������N���H$/�599)��)���3;��_9�%JJoL���.���d�e�Xc�@�Xb�H})�$�!��G���[�Mm�5^y� ���� L���;dң���2�qd�g����O�7��:h"xNm�5n����*rq�Kt���3g��Z�"� !_��eOFG]����c	"����7�KQU	�:��V���f�qrڙ����pk#��n��Q��̞�Ii����A�5.	�nb?9��k�W�!M�9�ހ&��د�B������<�8V���d^������-Q��Rj]�@i���p����9�^WDƶ�Ĺ�>i�!��M�O���=q���-[��׿�W}�s 3:\�M5�P���x7��j�F(+��TG�
a	��X���ʥ�rO	M����d#�7�z�ߒ�| >@Ų�φ�1��n�qp�}�=�����uO-��ꅝ^�˺we��L��*�_��a/�H�UQq����r�L�Փ�S��h@ˀb�^�ņˑ�A�.�2���n�.d=9/)-�L�)��4�Lf�e5�4�����BVv�MHR6�B�q4�[��D�7����Psd�T����S�k��F�U-���p �[Eeh/�h9��/b�2�޽_��2RB��0# VL^X�,[,�Rl��3BS�K�	_�"1Ӷ�`*T��C;����Sbh�Ӏ��(szŻ$���1�L�o�7lM�@��U�ﭪ&v�^��/"c��#f����⼬� $�r�[O�1w
�I��Mo�TC}�U�� P���<�� 'r�V��cr�cåQE���F+��L�>U��ʭj���.S?��).==.������<bi'A|9:��'�Ǿ�_q��i� ʀ~
���kY�q���������f2�9W(ڙww����J�ǠnH��v[dM�E.H/2$M�k�၈-4��m@~#��Px��*�jS���?lYp�D:$4���?�+`6�LO������JoTZ�A�*C��l�L� ���t�t
?����[Ҫ?Ό��:9tʞ��Y[!���������B���'�׭(�M�b>uˉ_�� �Y
p�f�cg#6�7�?�I�n����y���bŔ�.p8v���0sZ��}q�+�^��mﴤ(�:>�_=S�K=���k6*~�`��ū�$�J=����䀙SŎrE��JH	�oddĻT�����2,F�lh5 \����������Ǐߤ>	Ы`������舩��R�+M��T9�s˩2M9�
����f���S!G!�y�V&�/���@3̕M���E�6��@ԟ*��+�fzV!?��d�5�<wwE����ݯ�B����s�F��w��F(^MٛE)Ԗ�6��֠E�����kik�:x�m�[��mM\����QX�5�jn d�����2II9�9�{��9�A������um��, ��,�!d���i����]@�Y��Xi����4�	}�F�F�3������ߟL.��:�w&}�'���楜R]�aA"Y�������Io23�AQSSkZ��=��Y�=\驖)va����Ns��Gj���������-��;�l�����Ǔ�h�<R�E���ەޯ�&(C���T˝����U�s�h��U���M����"�49B����'ϧp$q����P��A7'�0ww�����3��.��o�����Rµ��h����h��h7��Ij,����+%k3�V�y=fn &�F-��tg�L�#&�J�>fGYr�u3NhѨ�'�΍�DE����o$!�V��+۟��ݽ{7�͙<S5����)o1�>�v�(��E#����Γ��ո&�ڬ�I>$�[ɿ}���v�@�}� gRo�]�/=W�©�LV��۽;p䒶�Q��^�X�w�2�V���Q\���;|���,i��ʠ�˽=�; �aaF[�$-�m��M�V�6�\8�����=T�5f����z ���7;����iN�_�;Ğێ�����mL}����W��O½�W�7wtt�8�c����B,�4}� k�9V��s&�`HK�Zi��»ޠD%U���6�R6a�������� ��L.��؆P���z�CI,��)<����j�P��#e��r�֌Er����
_5�Y�$'��\*�0Q~7�L��{w=`��,�
���P��z�3���o�O�d�	z��)����q�c{��@����,Z�~0�1u�>��?�zs6�e�[�٧�yfo��rI�_���z��4I�g���2��V��O���޷��0�a)'���.��ګ6%���w�i���"��32����uS�y�'�M�:n�*NNq��6�$V��E"�E��JŰ��Z�l)b�,zj�]1qx*�ʕ+�yYa���nva.�jm|ֱ��XN� śroG*ul�!��W۷z�H<��򍧵2Rj�;W���M�2bs:F^��.Љ�{L&��㣾�-�[���[���C@=F�^�U���6yS��
c��WֽR��禥��oh0^�,����@wSt_��`d ?�������']�:�cÁ���uW��-�F9;�l�r��P��ҕ+8[���*�n�g�>���dŷT|�9�a}>`4ǯg�g>���mr[b���}ؕL���fG/�ɦn�-�:�X.�����ڃ�:l�%�3\��҆x�R��+�
{)�P�b|u�p+��9��VVV�kg�n���u�p�R��8�tx]$R!U3ϳ�x�x˵�5v�l��9��ᢪ��=���jmϘ�
]��&����@�(\�ȍy�:ٜ����S�f�}�?`16���}�A���y�.�*�֡��,�p����PzN�����3��?��8�Ϳ�=_D�Lf�,�q%�Z2P��p�Өi��}H�F.�m#�f����@�j6`Q5�D\��s\�䣕걷y��ݼŏ��}����6	(qJ���^:�ih�)LgE?��285Eݥ���ɎљN��J�*��w9tJ��렗%�~��h�}����R8�5�o��};/|
��C}�I5�-�0_>G/1!���C���p�ڱ5���۱�;F�q�b������}����7�{���#� M6qe��JZ��$ȵi xsq3�N��x�6;�P�F��P;�����lH5eiY�]�%����nY��qc�{��	��hN�*�Icɋ=���x�1���t/�_��~��9�������J���i~���(���/z[��?7��)�hlE�ؐVV��8�X[Է�!-�iP;�X'����2�����������8f�n�(�Bm��O*R�u[qD�V&z���<n�uQ/�v�@�l�uh���/���9��1+�gP6���])��V�שO�Y���ɠ����$�6��0SvHonx�����,�����N�QgI�������\1z���e��p��پ �%������@���bؽG���e�
3���������ke�%0�1s+��r���@�U�T��g�

w2�k�v�-�o�e��$�]Mb��|I,�����X_`��R8r�A�闚l���2���޽�|˲��.���z�*�t��ͦ%z�J/�-�?ԡ6�ލXN����MP�_��h+K��Y˿#�ޠ��l��>�>P������ |f䒤�Ƃ'��J��?�ۢ{*<ra^U�׷���;���@�p�`1�����k8y��H�ׯni�b�m�8�����������ɏ-UVMu�m�$ַ��-*�2�������څ��H�s뱘��T<.=\𠅣�e~�]����Ycɂdr�*�տ��*x���3E����fJ�!�&����iv�P��6�ʺ��=g�c��/ȹV�t-^���(HbԒ����V� Aಷ����q�A�����f�9,��V��P�Z��5O��S��h�к-���&a^�؍�HhL!�=��j�ҥ�#E��_)ˁ�$
S�$��:��9����JZ$��+>ǰ����: �a�~R����A�2�/d��+9ƲhtS1�.<}���P#�箇����c��
ǰZ�pn��� ������/0�3R��	�����V�*r�tW�3����i-�	�CzQZ��W�V����A�V�-��(eCx��>�Q���Ƽ��۵kW���L㡳���Vwʤ�U�JMߪ���Ǿ��	f�e���Z�:�&�����G7�=#�"U�@��ꌂ���K�9�^�S�PО�@���VL\�l�LJ�!�2y�Ϸ�����0N%l�o��ǿ��dSol���XE�z�8���J4���۳U��T��ق5��vv<-J�m�F	�9�1��k�o�\<r$#�T�o*��)�K�trt�/վ|�P/��;n0H�p�������f/q������X�AK���&<D�$����1-�S�����s�B���mB�ƒhV@5�jRB�H����}�,qG�h�W�\UC��l�7������q�K��}K�e��p���x7�)�^M�������7+���&�-��ێjW�?���&&���J���%��	�S�X�Bo�NY��6ot�լ,�E(taP�p�b�}��333|+5���-�Z�zk�"5�N������ �\�B;z��'����c��NQ�с@�,��H��~U訽k�b-4�dR�k�����޲�K
��M$j_��X�����۷D�c�"�[��&���f1��#Ԕ�=�`�lȍL���i��KY����ݓ͚�Τ7�,�R�i� T�����٫v7؄�|��~/��b\\h��4Cu��N�������G�%�U���$����4�s˓�++Y�3ݮ_I�3ø�� 4��G����R�A���hO��Y[R�lt�����S!��XZ���IǾ���Gԋ�U��a��0�����W�W��
HZgf.��f;�/����o��oK(�H�|��LX�hϵt;�#��A��	�=�n�*wU­B���l�����kTc�D������R�< �!�%b�MxF�x�ST ��Y�e����-D���ʗh ��&��R�E]�:ɴ	�V��{azQ�8�|سv����3W]IZ�����;�Ϫ�?_I�����Z���_���w��6�f _;'��ڢC*ʹY����� z��6t��'��	E0a �C,��+�{����+	tx/�ż�~�gwW�KV�:	L��K�k�Q�e,�F�͇hm-�H���x�گؐ4�@�-%��@G5��_spV�Gy�ǈ�c��[2��p�L��_�jdX=�a*GXhh�K�Ql����?;� �#%	��G����-��7�UlȪ6���sd��}�Z�Y�1V�I"5� ��|�G񠐚�)���2����\����C���`�������ҩw���`��&>��l	R!���S8�<x�U;�9V]N����`�����h\z�nC��ΧOJj0|���-,,� ���cՓ�TC�P��LP%�֣����ȡ�q6~� ���q�B��±��*�����H͏FkV�F����,G���y
���H�������.�[�6�U�;m�'����f�>,��,�-�-�E�U2�{��q\?�!5H���o������*��ã� �!"~��Cr(ôPR/:}4� ~ ��Ye���E��B"����ҟ��6�F(4�]!���f���1�P��(���� =U�h����k{Ȧ �B����o���ج'��9�f��|&�\=t
{n/�Ӑ	D���t��������\�3�~i��]%�Q�ZU+�z���q�cl y���#�+�5�������[4��	hH��G�~l���_.�J�f�y����Sn)i��x�v����7�*�m�����`����k�e|w����jW�s���c����-�Z���:���6�4�[
z{��LA�͠S�MLM�<�"�� M�#����c�>}2 TXL�	H��i֖/C(c(��R��
1j1WZ��ѠJ5/z�޽��h�$��/_�Z�Eg_s��S�^!�j_0)Y�n����ހ�x��d��ayp,����>�����E���=������oqYMk0Sw ���1�w'�n��^���"�g�HO�"�G(/�����ڪj��M`Km�>m|Z�|
��v���]��Ě����Pɘm��.��EZ(Z��&,+�������#�;�:6c�bN�B#I&�\��+�I�iD Adr&����[�1�W�Nds��_:wծ2Vr#��$�4�ݓ�D�w=����V��`��2oܨ�I����,�rjRJP*��8��
���5����Sesʸ�K��e�L~��o��G���rV��]ƌ슻��h�U
��E�L���+%���M�`H
Et�Rf7�Y�4�n�޽A>t!+gA�����p�´��)��o�xs�h&��x�.��h���,�p�98)����4虚F�q��x�{ _���L���`��?�Jɧ���JcT���y�!�#�}�ɴ캗��?���Q4Gs|���F�1���;�A2 �Q����f����J�&TP���B��k�Rh屪�7ގM�N��ɣש�#�%��x\��[����$��=zz��)Y�߽����(2%�6�<��MH���3�py"sj0�'Cl�����
mE�6|:�<��$s;���p�xLH�ƓO��GX�	~Q̻}�WGYK�b2�&''��i+�C��D�T��/��uu�/�+�L'�h���-�cH���n"��T�d����&�h��5�maHrt�$xBHj�K��ґ��Z�'�ޱȝ��GQ�?�$i6�\d�,o��t��0���j?(�
����C�(^�Y@����H	��`ԡ�n\䠍 �:mg�~ C_�ӫ|,�����-xi�ضz�hC�l�j1�i�7ǿ&c���;"��7��:��FD�W�@B��#w�`F�`LmTW�����9��\H� �qի�4_�+�s�W��������?)�
�y�ܯ�=��'2:������� ��h��N/.���>T��8��Ss�syb�mw@vL9uqvBh�h	�5�A�Cݍ������!ʣ������{^�Z\W16g�^�N�K)Bs�����x�� ���X�/�O�4+v��g��Kq�,dB�aa7�}�%���Ev
2��W��c�5��L�r;�.x]X�E�C��?�܌��7rU��>j,2*�rq������;��@�=��]� yj���a;N�:ujo��a�nLF��A���V��f��g�p�R 
忂=*V��PtDKƞ*#l�- ��t!c#ŝ^c��6ߊ���N�k
6�Y�����fYF�A�ע���$�,:�8d	�z�v}�%�.�c}�#���!V�oM��O�I�p.X���7�=�+��E��#����'E�\�oĉ_!�\p�>��ŋ���$06:߭���>G�~m3�R~p'V��aE�[G!Zڿ�W+s;���+vϑǥ�=IT;�Y�8��Am�s��vcݿ�@7�l,E��¬%3i΅�­,1L%�#�D���GC|G�|
M�������Y��N/:%/O������!E�=�C�=��{ڹ�\ :n��<b�U�r��-&Ӂ=�=�=��ΊҲ����P,W���\`����WO��5%�8�&�'���^mt�T ��@.?���v��I�٢��j�Yu���% ��&�y�.�rL�'�"�F��D�|��J\~K�ߙ(���=@�tY#�Tm�덾��+n=�J��K�����7�>T������ׄtLG�%\Fǒ��������u�K�]cZ�V[��N�୿~XSXPq�*����Z�v9��9[=�s��Ӭ�v�hd`��s�>O��JEq���/��訆_nH�r�} dP���r�~��>������ͮm	<�
�k�S�4�؏�Oyz�h��h����06"i��?s�6��,�ٹ���7��������*�af�6�K��۴k�)0n���=���_l�C���Y�#U�D�:��U��E�ˮ���*�k����󝸉���#��u�S�n��#e�2}�gv�}G����>�4�}_;Ѝ���o�H@�N
d{*�BO6�1�o������ѻ񮁷��oz�Ć�М�����*�}Y���-X̡R�s��z����t׭5���)�'<%�Tp����[r����)M�-EXi�6����r��Ŭ㑝�c2M8��4��}oP�K�G�т��ʇ廱�/7�X�a_Gַ���>	L~sKj�0�'g�U�l���*��f�)�y��'�]^�97h�-��*�=z�݃��fMIsU$M(J^`�;��Lf��BXWۙ=L�k�������D�(��Ѽ072���;�i�\�4�˛�������,�']��޴4�7�)������ۿlx�h��cc����[1��f�@�o�~�Wξ>��@�
��.��M��}�^1�IL|d=^�N�X���G�:a�ž��cj�^uԛu�'N�_:��~��]e'���� 㻴��i�����-0g�����ȭ���Y�'B��L�@����w`�ܫ[�k}M�閍U:3A0$���HlǨz�#���/'��[���`�7�-)�������26�
c`�+x�l*��}�Y�L~�q�`��ӹ�W���kY.X
"��!���\�N<MX�a�L&�j�OT�k��sC�O�vZKԟC�p�gԷz䉖��Wy��=Ȩ˲�����k0��`�l�)��?'��M6�_^UMbX�)__��+�U��-~)r�{��kE۳��`�T}t�媄�|O������xѷz�a�@�`���*%�N1��Ж���GE(�Uɂ�3�P���nY��9��mk!+��n��J��,�Yp���]Upc��}^���Nb�m�1S�(B.VϠ`�?}F�sb�&Њ��c�	���h���w���9��)�l$�^�Kn,蒽 �B�����i����g�o���	�j���ň�~P���(:���E]��IS�$��B��y�-JG��'�A�hB���=5�ܣ�+����~�.���ڧåD��z��I�\�`�l�����Z4�����c��Y�����o�F�`S"C���[�{S�~%,�Y�x�^��ix���mh�?�ß��ʭ>7Y�S�J^=�*wk�������n]�SCM����6'A��B����%[>��N@Z��b�v��,Z��Q�j��^����ƛ)��$����/�"��&&&@0�0y�����胏:T��ش��ʽ�6?h�>=�*�s'����C�`*&E�-7�W��/ �㊄���}���٩�Z��}l��Z3�I�e-Q7���P��>����F��MH��5%�uX��ץM�x����wT�
�6ML�=���z�	>*d�Ua��Zl�<�ДZN_�S�u��@��M��׷��aJ����$�ؐ�.�\Z�]j������Vw�R�*Y��AAeK��J<�Ξ/}W��f�z��7Άr����ׁ+��_�=�DzN@ _>�a�}���?hib���m��� �N�����:���|�Coעo��?�(�&�(�Nj���U׭87�Y�L��`��N?ȨN'9���k[�V~+�+ך���*��2M�����g^zE+��S|	�P��0y	o����+r��*E}[�moF�I�:��H�!Ѫ�g�|�Ϭ,B����9�w��q¸Ľ[�Ϝ&?N�����Hw_tcjf?7G��k���B�Q�p�&�z��0{�AW���.%X.��'�'���3I�l%��~�x�n����q,���A���%xfTc��a�mq�v���"3�I���F���~�sd����5��V!�Zd֘��YI�?U�Q�����p2�x�U&�Aw��Ect"��V�0T:�?_<�(�OZE����Q����Y~D�}D�����_:�'�!�v�$����lF�g����|5F$G���H9�0
�h��E�u%w�DF6|.5� ��i��⧕�yG�p�\1�+6��V)[�@���fG�9�oY]A�60��e�j�G����ÆE���4��[�l�x,i�G��O���X������>�#����~�Bz�W�M�5��� =�m���u����VJ�P�^������fQ3��ٍHk�H��g��}����fn��鄇�U�R$rЎ�S�6� �\@+����Hτ��U�Љ���n©3��;�c��ؙŅ�&��]h�1@.���u$w����¼lc7�aj�E�f�s�/��/r�F�aE 7�P�s��{(B:FK<ť��j�=�O�|�l8����.=ٜ},BbqM�қTke���i�Q�B|���у+=|����4��I	0߳/�g-�Zk��I+����;eSD[~�I�]��1[},�)���L=Ѳ1�ɬ��?���ǭ���:�kW�p�����y��bRN���dF=`��c�1722���̼LS���ؾ��]��r@�S�չ�;Eۨ��I�E���4���XS�y�F��Dx��U�Q�"����`ن����d =U��^�����/�0��WȀn��_���;tGR�gzr]�4-���u��"�b��C*($�|� �P}���4�'��n酲`͎�s���i������O�#���VlpP�K9�KE�^��<=*��Pȭ�r'x����B�rHo�9/�A��<��{z&��z��zok��Ec���/��̐��&ֱq\�ʓ�y�/�l=�J�g��t8��#��j�F��Ce@�cf�/�|�/�*�#'�4va��-�L�JIs?���r3�p�O��&J�Յ���Jm0	�9����;�d���kb��16�o:�6�c͒٩�(��]��{ ?���-@�L��Z܄�q�������؅��Β���DGC��=�i����R�\*=�
Q���&�^�����R��*�������b���4-ԒL6�^S��ԃ��z�p~�}�w	��_s;�#S���Ce��B��p��9`�]����x3�~���G�ko#�Cn�W~C��8T�.29�����L�mQa��e��B(s�^Vײ��V�hBZ>�&��䥙��D�y���ѻ�������Pw���c`%T�Rm̼��teI����E�HF2`����Ɍ�QWWm 6�l�z�)�[t��ш�q&�́<=�v�my�;�A}�Sa�n�fccP'� *kAr��b�����Ԙ�<Һ<��P�D�g&��wE��3a����1V3o�������;�:��gh�ٲ�Z.�����Ͳ��
1��	��$
{��������O�c"q~0��hVy���S��JR��˂��$��l������L�%�n�/1:ǬI�\�}_���s �H�z����{��(��|8����x�mik1�m�_�:�gB���ُ.y����%�ywz-?8gS%�c�kLg���覤	�z�O�a�/����3 z��;&�:ˣ��ųU�Yh����4:B��p,2y��z��������GB[�]�#&ӹr�ak�x�v�_@0Ӑ�����EF�u��3��Ǌ�����h��2�B��=G&}r�?�������@o	��ּ�5|Q"mԂs�)����gx�!��5wݢ>_-��mimM6�Iw��V��%F~p��Ʀ���UPT��xY���2�%��eQ%�A�u����n�6Gˤʶ�b[��߃c���tT8�r����_l����0����J���g�O�X��m֘3��98:&�bS�:=Y,/���\!���V9�k�X6��O�0SrU\'�����=V���P~�~����� �"�opcP+ �2q�}�x��V+��9gk�T�2����N=P�R)��m0���3bj���<��vww��'�^&-Ģ��Was���=�����/I�a�1�m�B�v�ȫ�sn?`��j�sO�o�zu�F�nF��?� I�.�B_Ԩ=�^]�t����$1�6K�-�<��"� ����I̙ve�ڕ?���.����X0�]��wj^.��mLԹD�E��*zc^�.d#�U�v�x��>�M��E��{����b�z等��r
2��BU�!�8L�f1b�� ��a�������L��M���_��螭�G���lx�A���dr�i�`�=Y�T��@��N_TH�l)����?fDU����>{���������{��.�&T�L�cFR1���5��8������%�W�P�48~�6������ �'�=�L��6��i���E��G*�o�b�O�<��#|(K	�]��B�~�c�D� �6ꢯ�ی��s��<�}0�DQ��$10H�}�N��X'�p;B[P�A#�z���m�l�ސ�#�zL�^rQ�P�()-�,�YF X��e��Gj,$�G��%����M�q���J�����(u�?H�l<���|E��&�.��*$΢��-�k|v���	�Q&G!�%���?�'j��
�2�C��ī���4q�3_�����wC�o9
�m�d�s�6�^�����S�$��"���f4�Ԙ̣=�NŭL�m-�;wB���wКA��wd�D͑��:U�?h��I�	NQ�Iџ�oh�<�!��}+�`����#Hj��י3oΆ���>h�_5!�|b�������Q���ԑ|�����&{�$�(�8�T�U�mt�� Qk��K�8`�L?��F-�njZ	��:U��N_ֻ���w猱)�I��Зu_�$u�fkh�s@�.FR�_����ߌF+��?��;*���ވY1��HTPrP$JP�$HΡ�c h�$�$H�Jh�� 9�s������}���{��q�t�U�֚kΪڅ�\Ŭ�b�&5�$�;�W̪Z���������-��餥e������$1���x��{X��`����>D�ei����]0/�0/��ջO֥뙎R/�p��J�h����8u9��.q������E/I?L=D+��Pi�Q������v�Xg�lv�i\���Jœ	�4B�5�(�6Lmd���$*��G���@��T�Np����{��#[�2qg�Q4b�ĢЖ؊yŷV��!�G;��PՕy����^�iη�Г�������Q����6��2����Sn�lV����D��% )$$魲�UG�*,���8�y�Bk�z�m�}u#���;���nJ���6,��	{�puu�l!�F�b޸��i>�����T����ov�rGP`(����t#���d~��Hk����I��ۓ��f[|]n�,q�+��������ځf�N���ŏ`�l'�p�II̴��1�!������"{�[��>�!�t@��)�@�x�wBC�*�AN�	���y�u���	�ѝt��MDbj�sBp7m�Q�%�=$�E#|eG2��|��7X�s(��������u�H<�{h��4W�v� �w��@\��T.�l�PJl��X�>~���O���D}�m:�!��4�Yx�_�A�JJ�[P�7tz��y���sHd8[�I�|���	�m Wg7�I��>���E V��Z�^���,�&�����E��\9(d����z)��F�cs����CUt���7ۆ`�:9���;9,��9�N�3:� {�|��h�3�L�-���)�u݂p�DF�Hg��		i��)�|��JuE�vY99�-�v���1�;����&�����'%T튄�|�\�:y��s��;��L�!������r{?$v����)��0m#���ȩ��4L���5�B�E���g�T�ֈ�h�7�7\,��ؘ�ߟ�ߟv���������Q�O��L�����/����|��2���Ǝ�����A��p�����d��i��s��,G�ÜB��V�tmY�g��%��H�t�׍'�t\];�� � �t�8a;��V��{���OTUp�LIJ�S����g����I>�Ϛ�j+C��������]g��l+�k��kߠ&����6��h(�]�Q�9��8�RWwT���.Aq ��B3���RI�N6�����	��B���0:&��g$B��љ�; Ir�Y3�"�y��Y]}P9��Q�D�h��̌�lm:>5�J;��|�?����M�<a>�M��S!�"B�w<r�ֺ�+�ˇ�<�1�(>�XB~��+��`��W���5
��|k��+�,����F[�'�������k;F�k��>�#��(z{L".���~O��s���CJ�����lھك�>�X�N�)�	��B��[���ʱj���[d�s�M�e	������t�x84ܨL��Go���3c�okL�S��9�6/�<�!���u͚�uÉ�bNE⎢��iӟGҷ��TFx�DHy��UCc�8���.ZOqP8>v�|��m.��
���ɧ�>솭��6H?~��Tng��W���3l�li�i���K��l{{?�xLv#�|F�1 y�hZ����o*!`:
���3+�A��tY��6$�W�s�4���9=��X�����^%�|��q˻�f�Aee尃h��7�'#-͕�����V�܎qBR�O��P'nu���� �2g���������Ţv(�w�Lv$��q.���i\��P��O�0_"n�������WVu��r��Dq˃�^W%�CDH|
��!�V_�x_�7TN�؁��dv�>�MJ`�����iL��!�e(�'zE��JŃ���Ѿm��Ԁ�5���s��L���F[�s���E�fE^͆d�WF�ە���U9B;��w�~�Λ���͍6�/��$��=�H�����D��U��I�+
#KO�X�s2'7ߛ�1�uQW��L*�(�d�X���_�W"̈́7(��.����}�����u9N��$g���+���<қm�^^c��SЊ�܋]��F�e��ˇ6%Yh��V�a�]��J��Yմ�M���z������Z
t�!�� è��� 	�j
���s~�����Y�7__%�l��Y���+
���|�����E�3}�U~U�&l�Z������?�[왔ކ]�Q�0٫1���1��6���t�6�Q���%�63��J߄Ex^��Q�k�%LV!a��tC���Q4;\�p����<�3�C�� q�j��E ����8J�vӵk�d�䠋���>�Kk7�#w��Fgx�q���_��be�:�z�����^�������h���F�[|��1o����Z.�1J�{�8�Lwg�K����w0��/�a�$&��ρ3��t�x/#+�s6�?�0�ú=�=�1X5�Vn̕t+STޓ|��w2�d�YII�9�k�;�]�/^֡��a�6*�����.��Q�.%���@�,z�$��6c�`�Ё6��)J�
�	�죖��3B��{�w�|2�o����b+�h9������Ü(x�Z̧���K�wvP�ɣsNQvQb�����(\�qm�J��>�mE�
�X�|[��/��e�~�]G0��d5�N�3��ള.h���)�J�s�1��>��:������K�[{J~���<��oI7��+	�������$��	�	�y*� ����z�������<!��-}/[��C��q_@^/AG( ���k�� T�/}e�q@� Ŋ102>��Ȁ��v���.+��C$w�I S�34d5����_�}r��H�sbu���2���[1j��IjA�I����Q��R�E�:=�Ĵ��r����ej������@UP[U"�u�g��=Hz����Ns��5�e�)�Ki����C�=Y����s��Ñ��۷ёߦ{�Z�Vz���LR8q��b1t�ʟϿ6��k��<���<������ދQ�wT�n��b��ţ�����^��K�� ��(��ᩤ��8<�T��:��:�������O�ُQ!mC%����s`Jw�[�f�@�����5quA��[��v/:7*C�o���\��+��ТM�������]�9T�\z�}�R$bM�l��/�g�d;׾\Ꜭu´�Q�]���$���gJ	j�;�'���b}��o�`��i�E�Y<��A1~�>�J�x�s��
ƾ%D>�s��HC&V��^��9�ҕű�h�򜕿~�m�Wr�3��]<]Q≦������L�@����h�~z(��"]+��X��	X�LV6�])�0���-/(�0��y%����knnǢ��|�g��f��hhh��DH�Ǝ�Y<����07����mmZ������
.���G�|�a@w�AO/Š�,�Z�;x�AF��'Dŗ�e ȡc��$�t��h�c�8ǩ�h��@9�R�w��=�+ lgw�իWﻬBk)0��"H�
$��/�H���
[�*�ϼM������*
at^3�ώ.A��TE��7���SP�^�FGȄ�] )���9����q�_�c����� ���c��h���
[�1��$&��I�:�1XS�����ҽ���.	�O�x�����
�(�ڶ�TXJ���ˢ�W�~������v`V]��0�_�ї�a�7��X�� Ǥ�3<���|?��艮	߅^R�?�UT�ޔ�Y�1@ ,^�;�Q�O��uH,� ?N{M�N%@�(Y_E��C����)�?���������<���^9��	IJn�����${д�����6��,��]����~��r;����)�u�EÌ��'�\� gB���?0�������'~0���`U?<�����q��gv�_��|{�C���BU4(�W���Z@�[:��@?'&���}UU��z3�q�:�$H?�Hq������c�:���vf�;}7
N!�4��y�H35�C�� ʡ�f1!d�������l�Cy�EO�eѺ\(ה�dA��؁yZ�p�NR.2()ɡ�^o&���܌����Bђam@�q5�[�����ǩS���?�`�C���qD�'��Y�#�iךk�{���[`u���4���e 94��.��-�殁Yh�Q9�I���J	j����j[C���6�O�����beYh�)ӷ2���P����."���ZZZ�
,*���/�N�m���$��F���6$�q�jч�"��_S�P�9(�����I��>'���.��� �V�]��e��EA�G vH4���~��o�]�R5��n��m@.D�<���E���$�<
����)��
䒭��r�<�V���O�V���.�<�8��]���'!�U����n�-d*�$��A+;��}��Cu�%�`�n�'`��?�V��F������n7U.b��}�!�тGٞ'��}��va
���)j��T�[�۽���(�v^�h�+1b_S�'�$�{��f?���(�sd��ЗHI L��l$���~��qq�.�7 �|Q��t��l����i:V�ͱ)�)��4&Z��o$� �
�#��my�,[�h�P�mtgDH�vsf(� �
B>�X� R ]��8�Gb����N��˒��Gۦ2������n�U���W1JcW�ȟh 	U޳��@��/�X�\4��t�β�?r�a�9����wB�������F��Uѐ�K0/ر��:�y7���n��ѭS�'�M�Y/L���J�M)*0��l����8Fky�
����h���s����x6�@�}��ްm<?ܜ�;�qi���|^�����6�1u��ʪj��]���ϓy;���Vc2 9��mW�P��[e�S�X=8S�J�-���<7O]䔛�;е�80��y����2��e�BBw�9躔����z�_k��%
'�gQb��`hS?�XY���	������vY���+*`8:������~�*n�z�"ļѮ����mg�����Ja1�E�Xo�!���������2add��� Uç��,Oh����������ޟз_�/I^o��k�����U��D�SbS�{`��^{N��~Ĩt�r��v��V���{N�6��[}J������	?���
J:wc�=��ƑU��n�ǩ��ihh�g�t���G+/�݅-]�b��BXKk��Y��n	�#Z����.%'��	�ӓ��US���l�ײ�0f��~���X�WW�V5ӂU���	�o��ƣ���Y^�uu<��l���)�S�U�����2��'w[�0���L,8���G+�H���`��V�{��M8z�����ky�6,-b⢑߉	�A�x�IF�Q�����Uq;�-��X55FwK��%�B0lI5%���Y�
�meeM�!|-�˟��żMЧ�%���X{��������&���������U؛uL��g�R�R׾%`�+��7��$hT`X�.��A��ջ;j�X��ݨ�[�Z�''	��w�<3�ih|Jb-2��X<Y�:1=���Vϻ���xz����U'.�0*~��u�˅�+����&�Wߘfg���z��.N8�/���&F[�v�zyIYMNHn_��|x�CA�B;4���H���diڻi  ���l��,��zP��_8h���Y�RG��k��7�l0�de�n��A���aS�vCx)�lj�J�|s#�o��l�������4������C$���յ��![�������П��Jo��(��;BC���\�/W��8��m6�xi����yt~Ŗ�u	��>�e�{j��%7��߶�z7`�DP۽���U���GktAK�]��p������˖ь��#����T#���L���9�n�����zhF�c(��gS@���U�_w)�io��lp���Q���'!��������L��0ja}��V��k�+�8U�L`:.zCqm���ke9Ԡ�[���$yݺ|�g�ֵ��������/�ݚ��K�����u�����n�۾}������5�@<���gS���?ŝ]mxCK�L����7����dٿ������o��u��\�򦣝���|~�����慪���=PR�z�'~�N�n������M�\ݍ����ѷͻ6��^�Fk����h�H.c��Ug��������������j �tww������|>��M�ה|y�j�2W��/�"�
9��������������G>�s��l�7Orʇ�T.x�JDٱ|�T�M�aE�+����+�ژ�[ļC��L�6����X��Iee����PdKn����a�?Ӏ���dmi2/qo��]��K;n{p������9|�@\�����Y�ǂ���3��U�_ysw�������8���媈��Շ�~c��p�D���l]��vR���u��?w�H�mu	V��e�p��??b2�����߯��uL�7[������	Ϟ=3��1(rQ�|��١ϧB��~��f|�����խroIF)�����5�'i�X��hwl�x\~g?��
����\��jo�o�MH���R����q���=J�6���}�}����ttuee��xW~��N��e�����v�ؑC��fan^�3�4�.�^�́*��ӽ�)=gk�d�׌���*p�!�������uB���Ǉ�vٽ�=��{���n����ݼ��H%Y3��׷��e������z᠗/��9t��Ǐ7�u5%��s!�0��.��_��'�ol��$W�䘙��'�Kh�2\���>����C�����J2��BBB�=S`@k�R�;�S�@ݕo/'!!�΂���댹�=3cw���:��������juUUC���bwY���A�Ă������_�<�P짦�<�̲q��cS�i]c1�(�իO��.x���#G�p
	i�Vk�W�jh���̼�����{�����j�=)`��8Y�y�Cj��1�l�00�*؞��C���@���0�����UT!p3�>O�4��'�zu4�ӧ��\�b��iz���$5+�4;{��%"|����<�z��UR��l�4���SP�յ��W@�&&&�ȹUڙ�-M3H�L~��kħane~��m>ɪ3��|��Z��O��MMf���pq�2��­������r��c##cs[���O���cS�P�5������ҷ��'>>���i--6���=��v���O��?8����e_�;z30&�@�:miI����т'4._~ȫWP��l��c�y��k`�6�ϨSr��r���c߯�UǉN�)/}JJ�9Jl���U��"~EA�ٙ3gX$�=\�ψ���_�R��0��a�+�Z��<>�_���=�}=�^4o8Q��;����O�bQQQK���"�t}���s������߫���\���������{Q�(nj�����\P����^�4�Fkњf;+�۠D���<�P&���ظ�<{޺��цh|l����Ϸ�9��+s���ֿS  ؓj��D����y��FUT�w*rxuSӄ����
���K��P�h��Ĝ����s�ށ!�L�K 7�δ��z��y6nݍG7�F��bx�{�#u5��#\�������ϟ+�Y�������)�%� ��QHPP�����Gy��IkK����,�v����۳a�tq0��/��j�Խx�A�+�����Vn5U�֭��`�����{�gBBC;X*O�v�.!��ؚ����cZ�[=�����	"�C�c?�D�~��ܵ�>��i���֐��;�T~��C4Ru���,;b*�T�'�K��Ԃ&{�a���ǝ,��_��d(΂�e
z�6i�:�	d\C�	�}A��j���4%�ڦ�94-�/��a�'���l��)x����|�{�Ѹ�!$Q�M}�4��uSb������߾o��;����x��1t������H�o�a6����emy�Wvvv{�s:9�����A�u�P�Z�p�je����4��K�H�O��#FJ �N>��48�.5=�-=j��V�Ј�*t�:���ev0�c"o�+W��g??ʧϝ�i�d�1�r��ds�������h��|�A���N��k���KrdD=}v��AS�d�����އ4�QQ��1y����YޱCN��w���]�F���b`z85�����. ����I�����o޼i/r��	3u~��.��a���v�|��ӫ���+�^QMNX�2�x�����y��ɓ9r��m�uu
�xr=�]]�%�z)�;��r�/q�T�l�d���77h�[��z<�fI�\	���x��	o�2t�`�_ޓ�䆲�I<n6����]�AT��x3�!�O��P��	�=�[�|xc�%�c{�Ϻ����YX��o��<%G�m1!��M1˔�#��%pN�w��Nܕ��S�=f�/�2
z�8���;�h`a�8ڒ���}�-��Bn���#S�5?@���-njj��^��r屾׺��yE^{�N�܀]�b�23U���5TKZ g������߇�/o�D��P
�Hv�~���%~�U�[7R��V4��PmD��h+�1�e5��\���.F�ҁ y�^�P@��������K^���Cy����a�l%T����⯇��]�����Z�S�f���*?z�,��E&?�����=
np=���Xj�@���g�k-�P����!\}���J�5.0�#��SAA�UW�k^ww���Ƙ]4,�;xzz�ݾm�O9��L��e,|?��*..����r~~��o�T��#���7�DZ����0"X�o��f���Y��E��#4�2����]�/c�Z�!����}���&�n�k��<��X2���b� &�C)�H�V�J����3$�N����V;^���R�y^����҉�*�n������ss�KK7�5?~4A�T��M��a�_������'���[舡	��g�1��b�JLb~���U����:0.(T�zz�Ϟ��)���mL�o�4Ў����ɘÿwyyr(�i���=8�߶_en�D8�P�O��3�@_��WI���gv���&Cw555�RW�������j4?5:�������]��g��
u�����f���{��\E�	71�"��n�1��/��) /�"F������UK�n�r�32�۩��dZ䭒���no��kPb��H`�)C�u���C@NQ�s#�3��&���#?��������]A�(TO�����4Hf�>��M��3���d�h�J<�9��o���d�CSϏ��n�S|{���Q�ؗ/�*g������apm܋�D|_��1�����FZ} f��GD4�t�.I�(��oך�ڵ(�ϖ۱TJ�]�5�	Y���݊�^Ug�y�����Z�۔*f�	��ą�{33���NW�Y�Cp?u6��>�J��%(�����3� �+xL?�f�=����t�{8��ߐ�Vε]�L_��%��c�f q����s�au�>�{��e�L��$� ��zZ�-���kvx�\LR�����`�h���=�][��oqC�U�h5"y�%s����]ڨW�⛓5-:r���]N��k1/Q��H������T�a����b����*M/�Ғ��IO.���v\�V����@�e�Z��v$��J��cu�OP�x���kS���ꈃV��hg1��B���<��MQm�j�ӇU�����ݽfޕju��!��P�>�%?��.ͪ_a�Kq/\��(N����� S<�	��9��1�������v��.�:����R�(M=�`�Lգ����bM--CZC�۷QxNW�Yw˺8nn΁����.�<�[���iY-�;�i��W���21)=��Y�������<�M��:��� '�
���Xl7�l�gs��V%G��S���|�`X�����l/.���Y�X�>=�������Y�TXؑ�4�f�tȤ���5ix�m.Gm�/ϒ�<�����T�Ot�J� �
y��������������ũ0�s�=�� 300�q�-((���cf`ʧ�Y1��[?�;9]ta��4��q�}�\��)ţ�BR��.�7������jQk�c��MK��@S�s����tԹt5"^)��q 1w�̗��]ɓ�����@�d;�j����wB�"f`"{
+Tq�o���9�;��E�w{����u�t}�D�����'�aw��_	�[rm�2Dj�o&�����A��7����U�7��y���&��K�%����{�#]�~5(x��[1�K��"o��uyC�!y���.�cƫ��o�Gym�	u��O�X;���nu��O��3ۢ�7��7P@�R	a� ��`p$�A)9>�*0���������W�h=�t;,��:V'%)�P����w��D�KU�{:�{����9쮈�0b�
[��"�W��Ἰ��I)	���#���G�ﭯ̋[^(^��貒r�z@=&�j��Lȋ �7��4de����@���d��ߟ�9��E�|q@;�o8�(i��b�m
F�B&jҝh�"!
w/�����FW9}��&�X=�����H� �ۜ���N��[���uvH��8$��<��.*"�;�Q��e�Jm�㖍��)�NO���ǃ_�;r�IQ\L�b���\�kӀ����hEEK��cL�w/9;�R3	��Р�R���Y��}jP+�c$�C��FJX�8#""Vf���I�U@�U�cǻ����B�뫋��/%��s�g��" �=�h��$�Z9DG��oo�;шcQ*��V�@��eFVB��.�~`�֪��X�F���ӐǌD��EnKZ����+p�6�	���w���͛�x����}�ߧO��iBBM�C�OtV���X���5�ӝ� ��M=V�s��
D�C��O?��Ɲ;��T��39p�p�qk�Ҙ7,x9�&U0+���מ Uː�~�J`euu~}����T�|��O'	��'��B�4�����߿���3i;L�s��O�jl��i1_�?}B<#]5��G�0d�����Ո�&L�/�Y��t>q�T_y��DO��W�i�~H���j�����r��v��	��)I�AW�!1Q�ͭ ��O�V]oL�j������\�S�:	M��
[4�^�r��)�2 �����)��}�Y�3@o�У�B���� ���G�pց"}�k駶a�:��c ��{��Z��-��jL�Y� 46�6QP�$K\�^�/)��f�k@�c���h߿8Ҙ�u�d�YTg�HVE����}cI���������r9r$`�'�U�p�b���l�Pț7��LtwlXYX.�l�ug}�X��q��$�,qqu� ��O��w'Hf#ұÇ?��V�-c�[��)EI��,j�0\OLL�)��ߘK��Ӱ ��-%ճ��/ѕIS����b�E?�v!�^1�Х��3�#�B��#�~���z���X����`�b��r�E@�C\�LnnX�h}�f����|b CB���a�5#��i?DE�3��\�x4U_��]?|�ӳ�~699٨�H����r����<���A$�2�O)G� �B�g�$M���<f�Nt[ W5Y�9WV��s_�]_���R�4=�o�'��~6,,���rU� ��'YYY�J�-��2��'�*�Qyг��J��ں���-]����
4�%�t�5MO��<k�n܃1��;�����y�Ї�\på���k�~�I�o��j��������վw��O���}4^7@a����!�W:z6�'&�:bNU�������
�.�V�8�������`RR�_$������c�3Ҁ�s���tR�(ûާAk��OS�=�I�k�;#��%�5,9h��ٙB��ԅ�!�U�H�NM�q���蘝1���L�}�	�=Y���� �[�ѕ��9&�WnB�>{�\�f&u�y�u]]��P|� ;������'|�x�Nᵣ�}6ZrLH)2u�G�]��y����@��ꢿ��Am�N�ᦆ��`Lb������!\�Q�nhk_�����p0�����\���h�C�@�'���?���صs��HB������qj.^�n%Aě��J�'��ͫ"+�μ�q:���p�q4,���9�Wh+���ss��u��`�R8W^H#���ˏ���(���d����srr�`C&}�6�b' ���DU-�['���Y���������y�w�
�
��!����*..��`����:����;�E��$9}�9�Ц0���JXxCQe����ry����̓Z0'F�O��R��
Rv�-�@�k'�.(���73�@��I�mg:��Џ�L�f���>�MY�A�u1�������tڰ�����XO���puu����+�hƭf���"�o�c<��/i��5w��������i������扃T;AV��:n�����)�W?Yvl�fw����orbo���5N��n8���ʻ*�"#Y�SQѹ��Q�lj)`'�U���O���}i��������5��tAaa0O��������?-�`)}`5:z�k�C�� �9�3�ȉ�["��������Z�+
�?DTŜ�оϸ�@WWW��r�έ[���1�~�h(�o��".�p1�JA����3��'9���5�L��3JG&:m6� ނ8�dOq����~�-K�zն6@�LF�W ��8�f��<|�!⃏�٧O���X�/9"1g��`)�e��շQ{y�Ͷ�ttrjg�A��y��e���|]^c�3�YYYP}��o�ڰF@�b$�ܫl�C���(������l��')��f#~�^:sKĨ����ٻ��]��#���[�=��~HOW��F�O�6E$�ϊ>��;v�(�D�\��A�X���� }�in�X�]/��?��s`n���?��~��%T���|۝�� �kQQH�V���uwuݟ[simn6�d�g͗�/�ӂ�k�s=6���5@B8"���V�Q�~����ۂ�N���]�N���R�o6J,WQah�Z������M��q���yee4�qv�:j������� ���_�};���n�'1���ˣ=�D�ͭU������6�7wub::��}hF�<�7f������myX3myt��V	�u��Jok��ن�7AN�wv�2���o�����p��b���=�Z<�ʵ0����ՠ�5��wVF'��!���ͨ��sZ��"dBMc���9~���!�P�;Xvɟ��] 2����j����ATK?\��/���z�ͽ\K���][����mT�����l�F����_���XjE�{*���h4ח��B��[Kv�-*����J@�h��mln@�Y�`��*95�|d��j��^�/����(�/n!�^��[��Np��|���C�_�^E`�%��D��*v.���r�L��	gKZ��##h��ppD�n�2|��#��8zܭ\�����i��Q����~�G`��a�4q)���j(������.�$�\t���,%�GS�99��O�Q%��k�E���ޱ�.���L"����/��Y���1*�!~���zP����o)��g������DȌ���m�����낰tCRb�mlp��d���y�k��l�����N6x��&��9��`/��e�A}P333L����{&�O��"���\����8!�'Ā�{�<c,g����^~����Ǘd>>d�w���E^���ggoOt�gggW���+�hg�����fj�S�#��0N��Kp�u�L��gX{x���Hw��l��}$���%�n��OZ\��{lr3Nq�罹f�*?��^>���������Z\{_���ʉ{����H\(S�~��rv,�������=�ż����R���/�A[ۄ�"��H�G7�.0E�����Sr��$�b��x)���V����\�i7����
��|�8���|�����ٵ�A�^A���_����i+�b�>R�'� �|��zql��3Z�d�ġ�pb��e��ā�tR��q�y}���lAx8ܼ�-���EH���k�4ZyO�H��NOL��+��(�R�z5��~�t��===�Y7��6��i���kF/�"Hѫz�%���? >�pW�)W����U���#i����=ƃ�C���8

0Q'��t� �V���@B0U�3qX�e��X^+�W��ځ��
��gG�P��olp��^z�¥)����㯯����G��9zp߷?�ީ|v䭔WI�Xc��o;��z��sx8�"�ZW+∶�K���t����*Τ�� �&�ͻe;��Լ>[���Uw��IF�5�B�Խ��1W3215���0W�3��z̗)��8��W�˻�!Y�<��$�Z"�N��#�k�����}���dSs��F|o�eA 4fCAK�1$�K�xx������X {��v� ZѮ�˓�Lz�)����{���^�_P�y�lyf0�$';{d�gV����ȗ�sF�n>��~p0bǏNw!Vo�����ⅷͷ�i��.�v T�<�s����+����@�W4-�j|,���P��Տy{y�<"CP�@�C@������oajݩ���#'�#�i�ց�$fe5��0�P���?��&�Z�B�;zk�{mmˏ7�a~A����m�S�ig����Y����mooG�AN@�|�|�h�
���0�[�p6��;�O��[���A���?�U���x�Ç_�;!m��T�]M?���v� ʡ/`�� {�c��|҇򕕕gxy5�^�z��Wxm�3��:���{PU7��G\Bp�@G�r��
}�N�0<��um?pPj� �!!q ���wvv�P����E+/ڠ��|��hIQ�~��'��	�y ?�x%�-���pJQ�.|1C��޾�߲.��J��G+Q��R�u���>�Ĕ#S�PY�p���6q{-;!�A�GSc�d���qϡSf@=�) ��]�]�/�? ����Z�~��i�y�b[9L��$�Se�����N;bk_��JS�n�t������U�	Vy},��.��d́�WB;h�4����6q��\��+?[��N@O���\��8�A7Lyjj�9(�q����}����4��dddt�(��I����q�M-Fޜ���%��y|Go8�z���Ȝ�̏Aˏ3u�f}O��l�i��'����{�6B,!FO�D��ģ<:wO�	l/pL�Y35.��'�>>�N/�_���B빺�ҏ���>��dZ���ߑ�XZڣ�1˿^��gD�0���yVN)\8@5�ҥb��`��y�W!k��?�w�&Ô³��׃�O����V��mz�����o;����777k�\�~�1��52T�1���Ăp��c���=Q�ݭ?ޞ��kՕ)�כ�v�������7���b�\���_r����=�3wޱN��ǻ
5����Q�1�ɼ�TȫW:��2l��Q)���u�Y�ڔ	�����µx�*��x��C�1� @��0��
S�F�jA;��o�)j�1^�:��wݙ��&kK�n�<� ��?A8]�L�?�t"�ߞf�ZܜۃKF;uO�<�����1�Ʀ�b��]�NɞϷ놗!���C?��}�ŭ��1B=�(X�,�{HFe�C��O����p��sv��Gz\8�.��Oe��}ٔ�6���C�8P�0F=YC���s��/f	�&�����e��'�m"�o�lPJ��Yn��Zϩ��JraSH]��S��[���	��oHZS��!��$�V�fB{���MM��=;�)|)���5�}|E��?�4]_]D%��J�_�ȭ�&��`��ؾ�;�؁�Kj{P!L.�V�3��b���x�b�MM7�}���lD��T���p%�2������_�}��E+""d��n�)Ak?F�j���nP��"��'P$���[Ll^B@\`u`Lw	���U�K���l�4wu�T;:8|�\���B#��4/o��dQ0p�G��B�����ս�����!���c}�̥�$V����_�=R�'ڧ\Y]m!�J�LI�So�/�╣�G[���K�;�-���Դ�|�<��9��d���q�_/o�Ë�ŋO����T×:Zj�#����P���|8v����Z�4<�yC�۩�����a �Skn??t�EAa��U�׼��:��	9��!� ۀ�c{��"������D�@rI��	�g�"ʏr|�\��U𴱩�/�A�!!��x��.�jPJm}ss���(y��o��t��7^ww���a/n@<$\���5j�̬�[[Rom�Q�t��a��I0�d�n� v��[��xn:8�,�N20�9�y�6߽�����dKOA��<�����W����on�}� t��9_�a�Q9nz::~���Ó�@��8)��a�)�L�/�:Yz�����g�JK�)['��I|F�!�W������𘆎���m�ff��e�h��m������s�I��xZ572F��^t�q�-r���Z��٦D@)��W󋋌Q�1�i?)�������xۄ��k ��h�ȓ'O>y�:u8V�fʨ�'�_���<�������t�w�}��b�~3�J�<����Ҁ\��$"eӟ��俼�dpz�̳���f��w��Kb9�(��)G��8�{����� %fH�u�������0��L�g�'��VdS��Q����qЩ����Љm�G�b'��ЇI_����{���a�@�B޺>����r����8�s����_ߍ1��?�q���-5�
m�A}�vp9��qSkk(b#��Q}2�3������������bNc7 ��E�#z&�t�H���PVۖ������'{��$�
�\����|�١����L��Ņ��x�xK���+)#l"*~�B���]]]h�FU
�@��l�_��2q��d3mIM��{p�Z�����^4r�bLB��,K�{P���jP�N�y�����S7�k�3��:ΈD)-�n+��H T��D�55;X�$(E4��*��=���ʐ���t�u@)o�D�Ė+�����Q�*(*B� �o�4�̷� �߄�����7 +a�����D�h?�2c?��>���̜�X���������O�(����>�8��<B�+y�̏��	"_R�������J9��;T�#ʡ���%Uɳ��3�J�T��p�7�*t�d�`��)�\����Y�f�nE�|�g��ܵ+�6�[TT�/2
*�ܚ��JO���?�>��}�:��b��X�W���}?��cH�,p��ݻtb^w�>�:r���O)��	���i�
���fn %�R�"z��e��.e�/�N:���Z����5c��RF����g�RB�?߾Q�4��2�����a�a??���!1��7��?{�1�?V�i��$�M#��(<צ	h�8��8$%=ZSǛ�8#
���8���?[���%�Pz-��q�s�r���s/P�nؘ���sg9r�(C������L�s��VNBl�VXtj�uH�Ʋ2�l�)����Db(�����[��p�y��]AA��=�4�Q��Ӄ�x.G�`���eC��է���]��8R�ɩ$��Õ\��~7�R��w��D�՟,F�h뱵���y�?��o�jl��J��.^�(TPV�}�J�̍�=��"�aR֘���D���_����4'u��\�����*A��ihJ��Z�Ѭ랴�7�e:�F`g�]� �+�)����4�C��=��Ô[1:���Ԟ�B[���D2!6�C�;��3"��hl[��MJ�>�e���v�h�<Nu���ѱÆU�e�:tN�#���7Bۛ�A�������d�O/�ٞmA^��RI�/�C�\0᩿�G oS���߻w�mcn��?��f�}!���ch�b`��g��"��<އN�s�_Y��L�ϵ��$d�}��~'ܕ+W�Cވ�Ǔ�-���g�ǃDK�n�!�)wJqz�K)Aaa���D:�� �U�΅]-ݻ��������9�< �?8��4��uyC~��ɹϘk1>�}��h���Y#mu��s���E�R�lnk3Cs��g��.{���jj�D+K˦4���{3e��ԁ/U��>��C3f�~�3OskCC&�=J�?V�e5'krII�Lw>y�l�M۴�L�����$�������{�E��o�:��q��9P�4F� Z�[����T9؊?|��a���|�k����v�tX_qD�����|�T�����f�dJP��K@�-��B��p)�<<�e� VV�,r�x���hk:$���"�T�����{}�l����KJ:6�@�R��T�lbYA�ǊL�z�#ǎ����ݝz�>�����VF��Ơ4g\�e,�@oNw����f�	@�ʶ���˥�h����ޗ�S���*J�&�h�RT(�J������iKdh2/ɸLi�P�ʔyGR��q�)�$SX�+k�����K�{~��u�s����;�����s?��?�3��;�Y�ԖT�5:���J����"E��'5D�m>1>���6��ۅ�F�^y=�T���".�p�D;]�0�f��޾��>�ɚ����ND�vu����?�Ā'���`�V�鳲@�#�?�[�y�I�=�?�13�t�٭'��&�@3AϩW�3�B��F�|:�U2pk؝��U��b�CP�Y)���k 5]RB�,�(��ݸ;)D�dA��k��HA�"]˷����j�stl�j8ooco���{�dlp��߮��xb�5���<��Y��{��G(&��+U��'C�ss������ڽ�#_mڶ�:��4..$�'�],�[-�}De;+��B����e�l4	,Wp����3XB��B�3�����]ZQQQ^���������^��� � ��H��.	�I��k�V�ʄ�TQ�]�a��ʵj�-���<l��jhp9�����ԓ��-�}�r�P��(�]ØSfi�8l&�|˳�:V��2�>555�d�H{@F��Y"����g[�ZZ�-���B.����,\w~I�c�/;M��o����积!�(j"�kVk煄��U�����J�?Q�0�Nv��UA*d��8�#�~y�M�L����GQq�b�@WȾ�]G�~D&I�)�fq��=?-u�2x�֭B.�� .R��P���!3�P5�\ﭮ�^lMXy��A�
�*�;:44	�	��e͠���-�4fû��LŜ������<)<�����[+�o��+Yd�C1��S<�O�P��9A���ކ�=Ε(r�x�r��KU�]G�J6& �!�p�~+)���wf~��>)aV��ɑ�^��,ύ�b0s\������2�)[i��5��T��x�#�
i��79H�ƿ����!2��h�:�q��i]�t���ƿ!��8��~V6�������s��Po#�,�=q ?�SdG�X��cj����-Dbj�����#�������\�\��zt�����=��x��&#�qN�m{�:��ff�_��1���BJ��.�ԣR����o�"3�$�o�N6J�������.rV��˧�a�ѩP�c\??�-|��V�e�%p��,���7d���"�,��=qB����w�R�q;;dw�=R���'koB��4<��_˦>4?9xƝ;~t�C
�cn�;�(��|�;PqZ78ىa��aͽ}��bN�9���`u���lWB���	��;����&�z9��s��QZ��R
����1�k�湱���q>�������;v�R�։' �&�	�R�A)�P0�q�����s�,k�JI��[eQ\d%�DϹ�=�����8�
��8�W$_�������Ƶ��mGDz,��d��ߧo#s�AN�n�}�{�3�<�"����fR�C�� ��=-)�<�K�ƞ�Ϗl�IPθ��{x��.'��Z��/��ں^J�d��W���q�t��!�������{>��y�`^����r�릍�if�H�y5�8*�w�������u[^��+`�@s�􂭝�o �َ|IF&y{�U����+�,��o'�����Ь���A�����z�M�-ȁ2]�?q�����Tq� �o�|/�v��+�u�qdm�2�b�����/�eГr����"�6k	"ff	��?�,��}���8f��og��_Ή�%f�tv��V�3�ir 1�<��*BU=�H'E,���fLVVV�|��8u�/�����\�]�]�UA^��wo� ����\�5�s���}���`��5C�y��\����6p�k�V�b���Q���'ۋ?~��/�	��0����O������mr��)Ǟ��G�Y�l�W~_���*�_U��u���޹Zy�q�+��Ԇ���e�!�+u��A���+/����7����ʾ� ��c�I5v������G��U<�N�c�)4�F�CJì.SV�����V�UV(���C��7I"x����{u1k���)��"*���J-�ɰ(4��V�k��t�l���_M�������Jk;���$ծ�0Vk�rOO28���@�w*�u������f��T��ɘj��!�����{��պ��3ioh���X+���{]M�{����?k`a�����:���Å.�__��e�Ϗ6s��G�w����{k��o�[� �~~t��Ϗk�s��g,Gu���u%�"'�k��V��ڷ�#_ӊnu���6O���rꞛ\>Z�:�z�4�F���㽚K h��Ī$+6�<W��T�&O�)r���Q�� \�l�A�,ɤ9�I_�71��9R9R!x|���%�f>%KU~��XV��e�[�ǚ�q�������Z��Π�7��i	���Ϻ���nf��M/��_a����O���R�f��߷:BT9aIH�����t����D~GG�T�;_W���ZV������K�[�v�i
��[�w��\�j}(5��[A�Ǉ0c�;�#���:/]�6�M�d�|Ƙ�4�� V���r懵i3 Q���7v��y�k!��I-~W�r�|�����^�9ֲ~�S��T�0B�0B7��Un�����2���3^�`�Y�$-������������Yw4ǩ��Mj*��k?��H�o���)�nґ��hQ��Z*�/	�tRZk��~�u�ׯv+~��x��6�+�{�4AY��u(�	����T,�+)-��s
d�)��J���Eg��C�u��v�Z����$����a0Ye��gXl���C�

?�٩�U8���ɘ��K��y{Z}��o������[Q�ݲ��c�tT�"�:�"<�eh�M�l�Z�z4~����v��ߍ�C��n�⢋EXj����N��p�Ch�o�3�O�����j�Tj�㢫���Z��⇾DPg�;X���z��}�{��^�l|����}�fTQ�ϊ2��V���E�
*a��`���82��Ꮌ�y�Q�c��߳ �`q2���.����x����>�s[芭�m)����~���p7U�@	�ʖ�H-,U?��{d2�r���t{o&_w�ӫ�V_�HC�.���a///o�i�C4"��wO�����˾"Z�3J;ּ(�fC��<�ޡ�)�ڧ��_k��mc^��ن:���ޚ�����������y!]��	�I���=���2��\�د7��H��oEn���;�P(���N2����@Z���2�	��<8����=���z����lci���Ǒ�)�&�H,.IM]�<�����x&���l+�����i���2�~H�^�w?9�|C�E������ 2ܭ��ִD����Cs��V�Ls?��[{K�G�Q��t��t��� �>��>#����ݥ���v1"�խ��{a���q��&Mh!�rA��VD�	�c���(��$}毈	ߠN�I=��:���ۢ���������{
=ZGf&��S��N�r,�j�=��)���.|��h]�"��KZ����e��n58�q��7&�r�ˇ��B�9����$�3�7@���X�*����'����n�P�[I�s���N�Px�L���M����� ���=!b欑��S����y�/�v��F �P�Y�Qvt��"��Z@k��Ph����|�3o[X�<�z�<J�0WNЈ�]C:��V_�f�u��)EB�y�1}�q�w:]K��Zr�ooȹ&�[7��!���c&����=��V�H�w (�tY-�P����}�{;�ƒ�{�w����_�&�oe�ŝH�o5��ZO�n�� �܄~w{�BS'A�ڇ�!<WD�1�\C�
�V������8G�"�ڌ�f�,���OT��J�����Y{�w����T"�Y���`��W��OÓ���'_����贸�P�d�($,B��(���-�Q��l�<�&�0�j7�KX���G]��LA4�]h���0$�������:�q�~!ݡ{~f䊜V+S�Ϫl��ű�u��� �*�da<���z�4�[������{e�4O�y�J4@���x
0{�G<�B�X��R��2A�9�:�c�✵7��T����a���mcn��2��*.p�'����O�p�gǿͤ�����5��f�r�˚�'�:t���hEeVq��?����ª��z�d4�}��r�v}:���e��\�����qsā6�އ��;�ѫ_�`\Ɍ�}��xdd�4�\� �Q,��*�Mo)'tS�|΅��?�������/��Y���#=}�l��E��9l��D��Ћ뷀f8�p�L���
%_ Ό�Q�}���6�e��"z��Á-x��L��Ma@ֆ�.���8=���ߦ���j�.q$�����Dɱd@k�cƊ�;ޭ�}\o֫���p�������ݡ�T}��v�JPFTxEР!���9�:�l.+6�TZ��?��0��,yG�H"�X�x�=����F�v!)��iޕ%�7�4T��<�6�"f�)X���C@�*Pu�	��=� 9R�$"��^
����$��G�X��XC�Z�w������U!�]%��N�H�����	�tqw���:!��EL�����hٻ���Xy�:�	>45�}I�Eqi��ʠ!O���ZĔ����@�^�|ajjbj*|
憼!�<8!F�-b���ڴ����TC��!R,��P�����,�a�V�&�G�+�n���j]�
��@>�v��[j�%��e����Ԕ(���&Q�T�K��)=�3�GQ��[�'}<�'�M⑄�ȴUi����
���F��˿i<nҐG�:e� RN �<p�X�G�P��)�ܨ<�U�oA����<��9R��8m\<"�_"�����dw"C�������|��+�k��:"6��@��e��+Gak��q��:������Vv�L+2	H�+{ơ{e�*�yS��0nWP��O0Fd��~��)�*�kn�,�^��Q�����np9�C`GҥaIqt?�х����oz��A������n�2���S���mbJ5�ݦ���΁�FX����l^�H+2[aV�OvGl�Dث��z�?�����q��Fi������|T�0g�x+��ǥ�"��wpUyǥ9��?����{$�3#�9�ecMg.�F�Ǣ�[$�{���K����",eʶ�s�G,E����k���(k698�����J�_�V�柳ϟS�-ٸ��P���^@�Ƒ9|�Kd��ƛxܟ���oW���[�O/Fd�P=�C��n�މ�t�a�X��e�_b����O���*��[����T��l�p�֝�w�2l`��:���G13 �k�[��z�T�N��.3�^�4K��V�����F����D5��j�
9���
���ݎ��]B�^�H:�׭���.�P����*�D�Y̋*"�+�$t�ɉ|���n��a(�-��A�����W�O��yF4X~id
 ##��(��=�k9
�o�J�VMu�<T?l���5v ��jô"����$��		R���:���	��q�҄^��b+��D	�E;<���X��O-���<����R�m�{�Tns\H�����ꮲuk=F	%��(L�}��,��/ٓ�oI�H���4�)@}u��pC�lBs����ȗ��.=YY��m��P���̜����z_��t�E�x�����9q��nD�/�����@&c�Y��:F�D���A���	���Y�DH��5�&4�<��F�*�H�*�.I�\�p>�
��۱~�p×��M�������е&u)ٸcQU�������{��� PZ�N���")#����%.n�Y�7O��v��d7����=�{
�|b�l�K��Nӝj�$$�#IƶaH�F�>�����0<4�숼]�t��=ܢ����G-�5�������k)�����9�q���2u&�(�F}��KQaa!~�����k�Z�w�P�U|��!�N�~��$��>\є���{q�M�@�(��8_���[�=��Lw�;��p�#	(t���X�o��H%�� ��2�8�w�h�I��]@�Ӥ��&H��4�*�%�Ȭ�*G6��+Z����2�C����a���`�Dp"C�x�cR"P \L��ve��F��	̉�J�DC<��ޱ���U�	�&��֊<{Qy(@A$���=�{jic��؇0e�p&4'֙\���L�@i����h�%|M:Ҡ��2�5�rҺWJ���D������gѼ�WBɽ4i��.�f~����tRZA>�̹��T����-1�V�פ2��RSe�q㦁h^-���c��ޅ(����j}��{���y%�NY��N��T��]����
oZ�/��C2�������� �����[�/S��l������G/�F�3��c۞n��g�Љ���xx�)RS$��C��~~+���Oƈ����0^6�^�%���~�D�ei5�/�}P��Ok;�z'�u,=2T�J����iO@v����^��V9�p�^��m��Å�é���@��&�B���8$�����}^淪��=/��"�2����@��w����r����h�L��m�ϲ+�B~ߩ��8���a[��:�a2�u��Bײ:Nb�$���L��&+w�Th�{�Hh݁vZ^#'�8�5��ɘ���Z܊��,@��^c��S��	�}M]��y�z_l��� ����ሏ����<������s:mp��K������f}Ct��tm�n�%��V�W	3Q���\���7*����f�ŧEƽ�%k	��3��l���uz�C_�D��3������̤��Y/��p�4�s,ꑗ�'&2E �r�X�fW��fȪri�zL�!�p���P�kz���_�ͯYڨ�U�2:�Q�9d;S��Y.��u(D�'����X���4͏��$�(�C��"~U@ �p��@����Vh�3�]|��� ���D	�!y�����:ɋ�E�UI����-���V�U���(<WA�n{�{�Z�]��Vl�@�jF@�׸�qd��a��+t�S�gOOO�n��@��U�l�B����ܠ�.�wx�9�D(�?���,��ry��@�<`{��*��m#RKM���@@���5�����Ce���^��Ѡ�&�0��o�q�qk��,�>��ɾ�
[��������$����Rd���
L�����J�tw��g�Jd�O�5Z��#��<2|bk �#�v�o�/&�D���,w@2���j�����:L�ܭ ���֑��^�C]l���G�b�Xñ���r����..�,��b�-�,m>q��3�he�E�0Žg��Xz+_�X�2����)� �B�^1t73VV�֪��b���{.��?��\��/����t���:F-�uLB*�y���M��ڐ��I!��Y��r)}ާ��0B�=��V*�?U*�b�6�\�ϵ%�Lf�Տ��KO{Y�S��1
��G_�H50B����Q߻)��Β��[�-��j������PAɹ���D����i86Z������S�&y�E� ֮�饣9��{ҟ#-��D�]��qn%�N�`��̺��H��=2����^4�e(F��v,rH�����h�C����A���{�JFN�m.%�R��-�����z-��'K]��0�+��:�uPj�9�B�.�F�#�V�m�Q��k�>�4Y����yNj7��
����>���{��"b�W�:F�t�;YM�0��%������P��n����ߊ>�Xiq_�׾�e�'YE�:�'f�N���7lk(���p�V�LBs��m�hy��Ϭ_B ����|�i�O�_����w�j�g�o7Βj�Ș*��<_��5�Qҷ�n�+�Zb��ͩ�"biii��m�"/ϸ�N�|8H|�z�Is]Jf�z�~��uM�ZY!y��]�T��E��G˛��x|�	9���mtgo�1��O#�Ͼٟ�x\�l�E$nog�JE2^.(8���ה��V��u�fv����	O�Re�rjC鏚	���#L��D�
���R��K��2�so������W����B�_L�x�-�� m��%$������=�W�J��>�6�t��8�ř�7S�U�Mj�N��}(p`�w��]+�dr�X�-��4���=��=N�7�G�5����q8X48q~h����1����d�2	?��so�y��v�"6dnbb{�x��oy<���N�nMb䥫�'�6N�LkK]�=�͗�Ɔ���?��'Xv���ձ�~�xs4���FyUGL�����k��0ํ�԰�3��#S��t�8�v���R��O<nk���Y��u�њ~�2ie(0s'g����=o�����EY*PW�fK]�J����5s����ȍ���.�ąN�1�zEgH�B�tKܕ	��ܚ(]]�?�����V��4�b	��ŷc86���6�D����D8�. �T�P���X��g�bK�Tl$ �a��u%���n��#��"*�񆖸�={^A�4+�ʤ-b\�?�L5�IGH2��\��:]��O�@Qs7��Z�e�Ș�U!fk����V���ҡ{~i�e��n�� �h��"ʮܵ���K_�:R�Lqdmz]MW5�Y�I��s�g~�,Y\\��7��D����<k�89��,8y��q;QT	�B�i �`]A����� j�(��D�`���8�y���L���쐱�u
]yl�w��B��v��R�1��坜�X��v>3f��̕]�A��F�֪��m��Q^�Y�]�L�۱��ݝ��r]�Hw�3˨]��ĉ.�@�6[FQ��!g)6'e�	�>	�k�~�z��{a�:m���2P��5��6L�=�[��ȔU
�2��n"�q�1&�X\쒊�
��ǻeъ����C��OƬ��?�~ZȰ���{=�ͫ�I����b��$�=&\v1��n�����C�܌�O܁}M���f�:�P�a�֋��4I=�� ��j��A� ����B_ n�D��
��&3s�Q�U�~��t�H�'tQ�,�dpc�qr�B֚����k����)�Z���R�F��r
$�QdCM�xm���IG�i��ū��4g)�N�Iec�Z��|�� Y&��ɉ7l�}f�(q�J`�~�b�ݳ�t!��6�J\w>OӜ*�*�ƈ�t����hI��^��-�C�idIB)�QG*�U�g���Sl|��mp%��F��t�j� �8�8�4��.��Ά� U :�*�D��ӳ���^,<�i��I��Pt�=W;��37�X[�b��\zKmQ�V�u4�Ϯ����9��ǆ��3Jh�ؗ�1#E�ѯ��f�"O3i�������t��(
�aI�7��;]�Ö��ƃ���5�W�	}�ɐ�����$��S��␐w}��<r[^tY5�׎�D�T��SV/bI7L:������6�ˢe��}��,���J?��P�\>RQjmҡ��0�ġ&�@d�3�SU�a��݃�������:������J��FS�ʽ|h��LZ�Tͨ`�by���{u@�3V���6�z,ݽ����0�'X��0x ���1/*���ؒ��V6�_���`
���e�NW��R�:Qˌ���L�=��W^(�&:d��=!:�5:�OY�,����T�X�����,�>V��6�!�A�=)��X �G��n"�j�xտ��M:��ч�?��N�,�عt���'`�U�������W���6�*�}��p�/A}�2����t(�Ԫ�@���V�몬����8b���Ŗ�H�[�Z������z�;:��<��{�>�\cc?�²��D%��"�����.�������U'Ɗ߁l�	I帝�f7Ǩ��A�//��.ٜ='���PO��F�FV�󤲵�uIYh�vۡ��&�B��Ğ`�ÚهOI�-l�{��k�}��<��e{d�vM�	+}�s�e��d֧&e�_��lk�ش�t�O�~����_���{��O��Cl��o�=�{?�?M���?M������O����dJ&
d�}	�V
e�IKSv���^��Ә��V��R@�ltG�𷅅������8E����40��fy�3L#���lV���j%��Rv�¾�6Jln�-�fTU�fyn/'��Vs34��'���M:!�e�Zo�W!~�q��H=�@�jձ���o�
��ꞡq�������g4�O�4�O��&>kˈ*�zq�_��I^
lW��J��K�'o����n�j��?�=�}�5E�pr�N>3��M/S��S�ͮ����݈�?�^^�M�l~��%I��k����b�+o��`�7�(^�Ԏ��)�q�b_�n����+˯,�W���Q���-�lJ��XzTws���Ǐ�^�\M���8$D���]�Uڜ��s���uV�6c�����g/�w㱏�8сa������1���u�N+��*������$�jU�z��)������M�b/;"�2	x�.h�7��v�����g�,�J����
�ן�+�J���܏?W, qF}
۽p�C��U[��ikS�v#N�ɩv���SAxJZ^&��{�m^ܭ�b������1|�T��;w�"M	[��.���t�o�*(M�����])�3��U-�V�J�AдoRˏ6��|����Uf2��M��{��|M}�\�t:�l,�׌�x/�d��Yō�g�m"�W�)�PK[G�ڌ�@៯J��j�-���^�\����U__�Jx����k�/�5�$fnl��|C֣dV0?!�5+: �aC���(Y�/���b��a������ZƘ囬���S���V�R�k�`�9rD���� kZhJ�$9F Q|܎�zx�{qj[�mF�кN�y#�Q�_8�;^�z���ȝ�v#�z��cC�z�,�"�����/_���s��H���ub�Wܛ��(=�z�}L���0�~G��{'�
�8�`o189ߕ���"�l`�69M
�'���10<�G��qN��]��T`�^~�GO�Ì2Y	vpop��r���b��U���o�ň�ty��$��x_z����O�s���W�:R�$J��'���v9%��(�{7�ݢ���HL�7���79ѩ���E��%���>��Vr����S���%v{�L܋��U]"QH�YA�����/��GD�w�ޏ%���c���^.�Mʀ*}%��敥�ݾyޖv��	xe�j�>��l3���( �{:E������X�،LgԖ3]f~�,��k��)�^z~��+������4�����l�fR��@\�6��i�;��ӑ����)��4�Sc㲺��@��D��� (��1NJ�����!Xi ��o�te�ř����$G���ZWSS3����q{��y���m���f���}U��hJ�Z���!x�bwF�{s�R�u��;O���&'��p>��S��o۽һǟ�J��	��"F�����'�j|g��l�������n�݁�i�?�!��]��F�(��<iʹ*�=?����t,��s�)�����nXZZ✣�*�(m�Vp���3�ʓV�Rq*�2\wk���RSp�����+x�~|~��&�T��)#O9m�b?P�D��U����h$�'/}ԭ�鑸��i�裏���IF4Y�%_�Ql���o|Y����� ��е;o`�S�=����'XF�e��/C�c�y�...��w�.k��~�n¥��敥�b:k� �ud�~���^i���-�坹��>�%�wrVz���P����YIK������~/��߀zX�{X�~:��]i�Q�s(�:���t{�0��aDx�=6�
��K�㣳^~߼��v(L�N�|VW�&��n�q��[Z%�i[;e�:�*����4��2	�7"ܵq����$��_*<"�Bx�aWx���m����V���Ny������!9Ԥ������� ��Bm����ט˒�F��F��6�_*t�1tO�C)g>?�~���#�����N!���_��~��@�^}��R;2�F�kff*9~�+� ��ا8�^�]��%M�s9 @J���l`�*.9dٗ��R�BX^plOh��_�ړ��#�i�h����^8�l�Z�,Z��Z���HJ..+S652Z<Z�S�a؅��Y��\�-_'���Ӫ���k�s.va�리 �s:��<ԭ}�v&Na-g�h�����!�X2���Vv�:c�wЍ14���� bh���.MiB.]���ϙHa��
��zO7�;u�����������ad��:	��� $����;'J6_�-)YJԫ�$١V5�q�H6�e�ݼM���Y	}�Q!��<���6#��ep����D��@t/��M���d�ЈvЫ��=9,�?���٢$BS���@*�� �����ZU���N>%ēpKi�<���:f�Jr��� ""Bh�Do���T�Di�M/yj������6�p�����tkWr��d���c<�ݨ�l������@��v/Ւ���t��j-:�nDÁ�� �Jl?֣%Ӥx�3P�&!Od͌�B��Ǌ�!n�@���
����;m�o��+f�9�q{�笣���`� [����vP V�sj���*2�\��ǥB�'c�RY	7�X��aNs�?��x�b���� ����[	�^�
l3 W�&	���5�6<��_�%�n�/�.�J}���p;#3s�\��~��G�m��5�s����������#�<�Wa�3�1��"�+5�$D�]#w�?f� �7��1��DQ��K��Z�B��Z2����2���Y��5
��,�G����6[gF��ʦ�EE^������V4%{\BF&�������%iZ\;�xXt��@N;�s�?ab� ��`��ƹ�U�fgt8n�r�z��%9����( ɭ�%���gh�w~��ߘ�'�P�Cyl�x�u,��&���`S����Ц)ifђ �&�]�P D5�f�F�_��=�<�Xɡ����*�U_hc��yV����ϕ�c�U!^Ĉ�W�N���3�26��o�F�D������n��gV �;y!�?p�͝��7?)Rg�R��R��'&�/Z^��jI�,�dr� ����ÈW�i���:��*v���y���f�y��2ߛ�+����:�쑛�=�#wx�JI��.c9��[n͌�;!�����cE �����6��~V��[��J���� �s��۾�(Fr{����S�z�q4m��
M�
�ΈuTѵ�s*}���^�������-��+���m��f�?D��m��0>巵���e����_͘%�����f�ߓ7jFj�6��T�r�g"ʈv�:�F�ҁ|���Bʺv����U�;�YQ�Si�b��6�R��W���\��O�4�O�4�O��XH��nqp�#��ᢚ�j��PK   �X�X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   ���Xo�Z��  �% /   images/bf12b6e8-34f4-4879-8616-fd29946f5bfe.png��eP[�%����{pww���nNp���n�!�k �	�&����������lY{�OM���<����2��������[�￀��%�����~ I�
�z��̂�j*����z�[�<�`��% �*-�������`����>DWOEKB�#�����1ߦ����_����C&ͬ��������|��^m�f��y
}� D6 �)p��ht����j��"
�	��,5� Lc����:���H�.ِ�>�h �z�����=�g��` x8D|����)�v��w�	����JC�-����cP���wq��{'�oe�1�ˊl ��,M�\���{��Ē���ò��O�d���FR���2�o�	��"	�>��7�����,K=Μ��^�}�7]���a?;�ǟ��v��b`. �������.����Ӫ& %{w~��������c�3 `�OqU�q��<��^�g<�<���7xѵ<ڬ�-6� 7�hۨr�7A$u|��x�=����ot��_Zb��3O���*t����2�L@�Y<]Zm���%���А+���,�7:�;N��0vP�%���J�u��S��Y�B��^��݂yh3�����S$��p�Ƽ3ߍm w�O m��`K�A��%p�ֱ�/g���#S����x���yo��D��俖d���wyr���x�$M,�),s<�;,Pa����ף�U�?kr޽�$9��0݀�?���[�[���_���*�?�ۑg��%Q�v?�㈜	��M:臩���ت.����q꩘lZ�b�O��f���fף� ��� �]��h�쵲+�L���G�\�f�S�=Co$���B���E��<Cx��@����E���%�2A����#y�g�-w�8��w �x���9�=?<�3�?���1nRp�ϐ�Z�ݙ��B�����qz�N�N�M��k&L��t����[XK2w�ʑ8=:�$R�nU?x����/���� �9��e�@'~�B���j7�t�?���������$�L���v�!�;��.����E$�ꛭБ�����u�<�Q2����"���颰&ʸ�~�'ޅx��	�[gS:�/��ȷNONL	�Ͽ�K�*���n���#�����7�*��6kI���ZȻ9<�c���6�ܝ���;�7�����c�9k�$���w��^<4��%.����� ��	��|$��y�ז3X
��{ԍ��w+������n�ͧ�M@�����|j����fS�u�_����/`ٶ?`�h�w���*�#��-��^�M��Q�?����r�u� �G��ې�;���������<Gd��n�������+(�Rڼ�����!`��V�f�fy������8��\����7��ˣ?{��Cx�<�a�#l���yޱ:v����]����TD�@���������}'�4�j7��M|�e�U@=z��Ǯ�� ޟ�q�ߴ�����@�>V�t����2�?��@���M5�?�K�o��>�=�~�f��)9�H�����~�����O�����k[��A$��
/z�`�;D���~��#%�ǂ-���C������,��GB_����V;����{����p�������/
fx����xhl{�H��}�c	����Z�zD�q+,
K��(?� hj�v��OFF ӊ3�
m?��Qi3
��=�9�O��2��/�"��w�[ �'C���~������ w�{A�g����t染_�h�? ���3:��7�\���-�DN��6����ve�ľ�]4�ou�]�{�K�~CC��Z"���_��Τ;n�3h���I{3��������?��z�1%�	����C�k0�w��v�~tb й��I����(�Ǖ�Y�������o����`.���?J9@创�l������M���J �Om�ۨ.���S`Y.����T����KH
���^�.3���6��ۧ��?�c�Ӯ$4b�/^�(剐7]<�>�y<���ӕ�_K?u?fI��V�_8?#��?J������E��C��I�C���|����EHVfC��S|6�������cQ+�&2�����=�6��il� >r�Vh�\�����s�iČ���&�ͺ�MB�����iY�=��8��E06�oڇaCI�:ɩ��]כc�ZR�F�����|��T5�@��e�iUv��kC��ȭy�x�sSHE������ �ave��'=��!*p(uoV��4X���}(/������}f�A����K&�y��lCn����� ���˽��������Z@�������w�D���Tُ��*��W�8ރ;�|���8�!^� -�4� �P�Q�ݻ�-x�g���j��e�ņ������{���#A���#���}�?w�=���!y����m)��~Cu�����>7�7
.�m���t�cg��ֵ�{�>������?)NHR� �����I���*$W�Ob��1�#~9)<sk:�(���,�քF��#�=dg)�G�l�su?�-}*qymO+��EP��tc�g�嚫�>�H�,g�#*��#�8)�G'��t�����/�۲o��kEk��*���v\r3������ã���[KPFP#�.i�D�B,!-��aX"I,��C)2(�V�+�O?ï(�.K�4ް�84X���۩����m��,�����p'0�8Z�j�Y�:��D�Z\���;�@[ZTc 	�3��k*�8�灗 �k�]r�C�u�6�s��[�,<GR�w ��'[&�3�:�1X����IJ>z��`Y �!�ך$���g�\/X���B�=TK�(7.@�Xq��E�ѣ2��jF�C%��cE�L��Ԣ�Yԋ�E�i!����_
�6;��e��7���J�LY�3Q �9�Zme9��MXO�cr&�u2�-#�3N<�X��u"�������2B/,�\OĄ���=.O���&Z*�BUz-��M��'�<����JЈv��X8/,0w�R��}F�rLU�X"&�;\9��P�zOJNDq+�X��{�jT���B�0q@���I�w�&Nd�_����[��M j8��"b�y�A�X�A&��'���rJ6�
$*�8)��MdJV� �ԇ&8d3m��zҤ�"1W}�+�mJ�X�����v��9U(����Kn�t--
%L�c26l��b���n$5�y��izhyf�u����7��х��uIń#R��O�$�,{&Ϫ���q^�Zv.�$E�7L6XJx�������ߜ����c���(+P��,�&����nFבFx����1M����̍��_��$��9j����צ8Md�A�����6���I]G����%�����ӗ,�e{%�8�*�yV�b����V]e��	sW/P�������Q�e%eO�U���#r���:����\=�t�0ը�.k�}��	���ƙ�<���뙛w}�]����6��G�!�?�����p�����l?P|�}y?D��Ф�$�8�l@�G�FE2&\5P,#��"g!Y�<\9.7�Cy�>N�u0�X�L���2��L7t!�S܆B*��h�lL9�l1�/����M��R�Ą�M΢�p�5aB"���Tb���d<VD4x�� N��hK�<DbqI;��-�]8�M�f����yg����B��*37�-=�n��R�O&�&���zE:V
�� KL �.iZV@¨�c�4�4*r�3FR-�D�L�����,	�s�|E�$Ѥ�Lp�R(,�e�C�@� 'ђqsS�,(��#��qA���W��p/r���Y2�V�����sob	�d�7��8#�V$*��1��wy��$Rʷ;�r�`�vX �D��9U3�t������Hu�g�?��13�6	�e9��<X������(J(�V�i!�'��)�H\�0�-�P�(2!aN��'�4�������q\��R�!��YgC$C��#��%$Vp��,�i��%��Z�a$DE"Kr��о0�3�H�d���fD�7�d^A���sw�&x���s��z5KȢ����@zi$�1%cc��eb� ��0>iؠ���i��K��#�����Cͅsq^�{��1�a?�i7���U��L]�����~G�ز�W��{�3}{��S��@�-����������ĢH0��
�2�S:/���u!�H�LِT�x&
~_;
5�,ނ�,�A�$�w�ZD(2���h�n"�x�b k�~��DǛJ�;Ht�D���y�i��:Ŷ���rz��n�\yM�l�H"�ey�u!��L���W|;-��5� ���8��[<2_(ax<����4�%=���nvXX�- �"��`�8^>=w{̒��A�bY
�HJ��-�u/ZG��rG,�v�m�a�+-G"M�({���Yc���Q�B7ʒ0j���	��"FCy�%��u���PL*�;赪��!�5��!��-)LjH*�?c1�fn��	�^1�_�C��gI7�]YF�%W/�ۺ�dѨG��y�\>��0
%���rdп��B��t�O�3�E�����F��g�j�r�S��ر?a�L�2��p�	Y`�*�**G�~�Obr� &���"�X�?�$q55҅d#&[�61K&�	����5<��qΰ�:&�Ce�G����&��x��p-�߀��&:"�b��`ΐǨA�p,��!I̸t=���+�M��M"=B'��Q�āY��ß��^mh�8R��!�Z�1c��׀mH
��NM���|
ۛ��fr���(���_��䷹T���qn����&�c~.�|���1��w�5�qI�gs����L���	C
�efŨ�p_K�5 Ry0e��9Q(�@E�*��������A�H$�Oq�ǎ�Zp�E���J���B\�D�u��Z���$qf�4%6��8oj�vq�W�
e`����f
s�E�)�ZR�QbK���K�{ĥ�KݓE��_��ZO�Q�f�h�ʔ��VUJ���#�ψT�ʪ����d�� BYR"�$#k&J��C��db�=r5�Ij���6�1+s/���MN�i�GXV���fB��"7i���ʌ�n�Xf !G�Vb�* ��6'��/ 
���!YՈsBHsH��� S_�Q#b����>w��1�%��-�H�3�W�wP��eۉۀ���-�,Y�kd�>G����[���	�)�Ϭ���D$�_F���R�F|I�zU�4V_¯9*%*,��)	�*�M��&MAA�^E�7K
P�)�AHe28�!�X��Ccϧ����π�j��,��C0�5y�s���Ȍ@sۤ�� I�$�z;���}*d}�c��Q�ȗ�X����?"��E��(��I���C^F���C@�;OJ�	�܈l�u#ǘ�!�Y0����ǬH�����x�G�sH|mG�	d��S�b\�kb�䷸la�z�=� �O���;�')`9"�o3�{�Y����֬/��c8������b�5��r{6��z���dco����5)B���6��������5Aְ��JF���2~���e���ʰj��@�=�j������y���Ѿ#�a�p��R!��-��T���,���`H�����(6���r���E��Ѵ��&i��x�������2�,�rG��F�-gA�8���[5	�_;���8�-�pB�h��N@�B�D��/�<�Ga�M�aF�J&P�`��\���l�M�~������m�\L}<Vc J��(s~0x\�ۥ����$.4�k�����Z��u��pD֜��6���~�w�t�Jӊ��-ۭ}}UJ9�}j_���dv��2�z��uV�q|Y���Hj���n3v�����!�hB�� Q�-�^���Cw��Hh9gd��G|���k�"��b�3�q�6�3aD��lV��mY����	��6M����)��{
ck�8V���DО���DEr ��N-8z��ҁa�/<P�^׵4&H��E�p��D@mCr��?Y��tE���v�+f/v���n��E5}�bc���[�')*��<����kQ���ǽq��f᠟���ꄻa�F1��V�H��?[��uZ���j���	o�t����"5Z�/�y�6�Y��l�9���]R4J?�s�1a�)�ydx_0~�/=&M���4�0�5�<��u�ĺ�+IZ��d�G�S�|�|��+?&XZO-bh7��s��mͰ>��,�WF\�b�Y����̩k�Q��в�'�Y�3��߆=T�Jc$y[�+�!A���+u[�Џ�_�7��h�h<U�����$YM篊k�x��ԷHR���\p�	��2 @ f3 �yzv���4�:YS�J���
�)I���A�zs3��d�Ǉ�3Qtv�G�>�q��13�$��sa�D�([�p�i��ؙG0��Ì��"�C+G�������{�E.��㗥�䡂�5�"Ed��3-Z&�U�2�D��X �b���}�%�]]Gb�P�,j�K���l�|���+A����������q���G�T�pE�WGQ���+���T�⫫YaU�&^+��=xl�h �)+l|<nT��)X����:��"�'2�X�S�+�"]د*v�2������5`���cԤIs�C�����iJ�u,��ﱊ'��s�*�Os�Ϊ&�8|.�G�*(�� 
躡A?�qm֒��GP�j�,����b�p��!���H-=h��f��rr�hY�,CT��F[&;�w~�������0�
غo}nxX��J�K�;�[>S�/�.�����(on��]����F�������^����Ic�r��}Z������6���I�}.Ö^}���q#6�zl��xb�#�j&�#QgYJ�-UP�X�"A �pTT�zM� ���|�KI�V�ȫXd�w��8��1���rǨn�t���J��K U�j���ˍV��K�w���60�����p�_/g�0Ƅ�U�Lw�SG�dq@AӘ�0,`qs�,�KLbq��.��18�P��� -z��g���Ps0Bn�V�M���s�V	�:#pq��@�X~^n.Q��e�����.dr�CVȊ8eJ���Z�!V���tYD(T��Ʉ���E�,]��<HJt<�,!�A�9�0l��a�g���j$�C{%�"�	:	3�m���q�E������H���nr�����Mc2�������`�F��OT��=��=iy�~8QNCߖPw��w0��0�Z�s�)~~�F[��*�DW�sQ1�V�p9"�˨���U|+$��5����T�����˩wٟ���T�̠�xj�	��2����a���Dd������1h�O8*x��"��MX}Hu����,|���X�U���uB�갼��qW+_K�� �,+�s0���PZšy��G��R$�f��I_$���h��#	0����&x�L�q
���e-�b�YC�h���̈��l{�wJ�2�ϘEJ.�/c�;���{{;�8�?݃IEv,�e�{��B0�O0p�����9r[�9�FL���Ƒ�"X���:���ڋe�zR��ء��KK��Į��/����.྇�C����=�w	�/��^K	T��
ۄz�4�|>�s��zؖ�y���@v����ϩgkm%"�z�mM/W \�wf�8C�`�ih�>J�:����.3���1g�j��)j�J�(�xo>��8l����ZoC��v}��k8;Q,�s�������/�S��Si1��x�@��w�_\�������1Ъ�V���{e�L� ��V=�!!�n�<�A©1�#�$(��W�u���/�%�z-�ԁ�N:ʨ�/\��Gw�������̖+���W�U�����*ᎉH�x5�����\�]М����<L�ȡ���fA�2ﲶ�*�0��՞�{G�A��P����mX�d��gA=e�E��s�=?6�9��|��ec��ĸ��U�+�4fN��Qb���Dz3L�O�޷��m�ͅ���A����=�m�$'�)�u�\n��T_��v��~�Υ��c�_3m��)�"P�
ARqf�5Kgއ�}�
��J�D�3bU�\����5��esƂ �@]7��@���Տ��ˍ�|�}1�_p��(��Z_��Ҙ���1�Y:�n︮]����p��ې�f� �FA��2}�4^քdx��1q�nN$Fu1���u)��iF0��pX+�����m��ں��$��Tc�1��S���[����
��'�F�]o[�D���>"�}�W�7�����W��b��^ĭ6��]�/�K����[��ȡ�z����w_�s��?�5ezO+�Z�����_�Nď�Y|��z��2�����[��8�Brg^��w��lu�`�Z$z�y���E�`�P��5��$3�ĕh��6>�?�\N��ӌ�4��;q�h&Qʄ@9n{x`9b>}�Ҩ�������L��Q���t[�%�|�zGJ^_+�����c��?2��Xʕ6�+��^AY�P=;i8x8�}׶O+E�p[�H�Tvh��э����p�'~� ���/���j�
��b���4�(]�I��M�nA��e�ZT��[Hm78�he<�ѝ�,<�DS8�b8#0��J�
5��KDc���K�p-�rPo�R�����Y��®x詂)��2"��'X8--��?�ҰD�����Ui��Jr+t1,U�Ƽ�����{E����$�B��Z���D2\ �e���u�qHg#��6$ʐ{���|n]�j�����O��}�x��g�6�6�%��
r�t�v�a�x�hr-�n[��a�3��ty�An'{`:����syQ��<J�����wC��:���@:�ب�-���B���<�L���ݡ����5E`wpq$��t�?⥤�
��h��$m�Bv;�$'\�уZʆ�?Y�	\��53	�gN�/��a��40/�
�c�[��Qk��2�������2}:�݈zϭ��H^z�|��33^S#�F���p��Kt�g�Q�RRBF={�gNѵNO�96<2����,	�O�ɑW�>=��}�ϭ{u�xK[n��
�L���r!B�#�T��UGy�e�Ĉ���ƚVך�"�E�l��۔K��ٔ���	�g?��M�rP�&�>��j�T� ��e9�￢PS�9�Y��z{�#'�3�[GS��`U=�s�� �o���͝4�Q)9.���al�w��؂yٛ��\kJAI��+����_�0�H�˻�KW)B:���DM9c�(�*��J�˨�P����һ��Bd��@ �U�UMb�y��
���Hó'�VW��)8̋��qG��Cx�G���c��ڦe��宆�G�)��й�����>]̐�.��1q(Td�N.=��Bv4oLc��F�tX�s
Z�}�:���=���#>����瀂h/pN��͝r;V�^�� ?��tRu��B��SYP- ���:&"��yN�ѧ:�ybD�CǼ�fږ��n��Q�c5���+2���RO�6�o�9a�����|�������ڬ}b����E���̎bp������U�{5���g'vPuqyn��זk�����ג�17D ���|G����j�b��ۖ����㒼�Ü܄�&���>h�1f�ܽR�ڙf0"�2���W��<$�pU�ֽ)�:�E�c��@h���T�p��o6z�xG9��;��$栨�X�~�{�n����O�}��>ȏ��ჽ�-5}�~޴���[ 	d��t7I�6/l{��t�7��
���̊��0�G�\���v`�ߵ������GwFR��`�s8lj'��a"�\H��nd1����#�~R���\���f[�d:\�V����w��ATw04���VE���:/@l4�~�_%�������A�*5�Tgj��y�W����a��e�󭍲+ܗ[�b����2�1���������Z��<�
�Ϛ�'�5Ae|�6V�X
�-X�Y~M	.,��D�m*��zŵP[e('�;�vuǙ0�j�b�A��v=T`�P��v����1�Lal��Q��yq��TL�A�w��hk��?�X2~��\�˾͜��@B5&GkЬ|���`x�T_�<�۝��섋�)c���
��.����q��WZa�?�9�I{^X�|�F��$!�2�>��:�Ya��^�iV1H��kh��f�5%Q�{{$����S�V��M��������)�[5�#d�~_��0���U� �f�ϰ͆�h�0B��8�aC��8)�'"��?11�Vk[0�^�/"�&e氃��+d�������~�'h��|7���
�WQ��g�f��sA��
-�T����m|7���@m�Wi8�" ��K�r?���ܜ���1)�:J�6�Z�3kQ��������m�=�����%�Xb�ƘHɟ�.�d�d�z{d~����l�U8��dc����C�Ӥ�P"�����)���%�+զ߃U31�����F�u;�7	6p���
ǽ.\�+Ց�G�n$��΃�Oz}�w�6����t?�F������k�/�dlm�nŎ6*V-�.~��#&չ��p��	;�l�8��Ύ�T�UL����P���E^S���oJ��Nw�+�������vAE�ʬ���\@��l5m�M��0�=r��Z׽BZz�����?��"L����6�z�K3���7��
O��O8���2-W�LU�v
F����y�@n��b���N[w�%=/����0�@?>[	J����@�8M}{l/�a��-��y�̎�\)��.�l۾F	�xŹ�V���	.�R�e�[>?M>+����n=<>9�@D�l�5"y�;����j@Qk�
�s��n��=��V�?Cpŀ�ժXMH�b��úI�R��Js�}i+r����GT���=��RU�{=���P\"��M�������U�ܴn  !�Gum\+G��J�����5a�2��\m\��U�V�F��c������$'�I�fY��D�W|ί*����ڽ�~���ƒrq��-X��p�;��(��	�V��F��D�]�FE��keԟ`� sl=�נ�;3��A�n�]�mB�Y͒�Egu��2<!��(��� �h����K��>��~�q1aּ��� �����y�g����=����iOa��0QS�!�/L�MtP>��T��U4P��6�����hv���~����~�c� ����;S�IЗ�NF�k#��Iu|uɿ�Zܺ�ĥ�����؞���]'���zY�徱�>&�SvK�R�A!��}h������ 9og5<ga��D����Kv���*@��qQr^OZ.R�T�^��o�df�A����{��{~�yA�1GW�����T�^0��ٌ5p�Za?q��=�Gm�:9�I���%�"V-�{���1��]�����eN��f��a��*N�h�j��wq��*dr�v�r��
`ͮ�x���?0Q�ی�RF��L��_S \.}pN��G�P�*�$=j�]?��
<�<����:��M]lq͑��i����:�D0�?���L7
���~�U���R�b2��,UM�\����=�%��_�f�K�uϸ(�q��˝�����<c� ����,u�	f50^�0��ZK������Q�k>�dQs�] ϒA�a�������Ӭ���2[�Wp��0'G������R1 �ݫ1N���@f���]�O��k́�U�A�Ͷ�볮=0�hT��V+�4��2)tJ���oSI��_��
̲aA����u u���:g8��ہ��q�����v�w�ϊ��^�����1��u��!���W�oO���y�|v���U�sZ��������h鸝�vs�2A ���UmJ�6�2?S xF��gQ�2w�ŵ�Ɏ��;�r���h�9%�'��h�cEYo/�RebU$��2��_�m�x>��p�d��%�a���C/_l�WV��e��Q�
�`9����h��TJ�pL���4E[H��*�LR=*X~��Ҭ7L�+��e|�'��QF�s�u����:���n))�	
n��G��:������;VqȨر�mj����ˑ�aX��n�[]�[郜M|�����T�kzŤLX�;6�1�5�L�!C��0xTW�W&8����م,�x�.��������r�U���6/�/�y�z��8w.&�x۬�Ŧ��1�4��׀����\�������JE��qe�J���e�F�����3��|�vR�Y�d����O�j�uG��W/~ry���3��I�޿���eoA��
j�^�gM&7�U�
X^f�/��m5t ��th=Q�N+ފ$���������EE(�3��o�WB�_����{2*�u�g������L�:�qw�s�գ���#���`��
騖X�Y�8h4�OQ(�s��+K����`@�BT����l� eCL��۰�A�M�]�ǐ�bޏNp�,�@̣̓�;/%���h����J�mº�w���PxxN1���5�����G'+�[�x�����@��,�ʤ���1o�M�ᳮ�&��m~?5Y�jiX�UO�	��x�f�'���^�����F���J����a7-H��&BG�nƞ��+A��D����(+xK�J�E��&VN�b�*w�&4A��^��"Ǐ���g�m�	���c�Z$>ߗ�g-:��*�3���9���ptT��x�.F9�N�����c��"����'�hI��_�3���4Ye]�������%=���g[�A��xE�Gu@�(�\<W��^56�䭯��7�c^,�����&�O�����^l��2S�{�f�^�4�,j��-�[�W_0O�w�B �.�3�������-�����[=>��|�ᕶy=��
]O���`E�[�%���O$k��=0d���Cr��H��C��\���CR3�`�j�>�X�6���ѕ{|��Q,�k
C�>7�~!�����;�.�:�_��")��\��98D�I/�Q�G>#�>r�����=�k?zj�ƻקv^SZ�������v�4iDiT	#LTxO�ت�*n�-��6Xd��'��^�:-�`���s7͸�Ag�ܮsM��`���|p 9�.�@.��DG+���/<B��F�u�Ml�P��C����#��9A����#�����/���g��9/�5���g���"��\�p�޷���\˳d'RWI�tz�`��:���B��d~����B3���2�b췺�:��RE��P�aܾ��&���>�ᐟY�S�%�Io�"�t�E�x�Vȗ.)U�y�&|��dքٖ�M�ͭ��:@�6�YQ��?������k$���^.�$uB��k˾��7��h&rPc�G�+�G5�6X��vKo�}�e����[`i9�w��j-��S�O�"q`�8mu���^�&�30oK��w��ԲW�k��� _���,���[�1����%9ṋ��������~���*>'"�}����X|ׇ.���A�Ŗ��{�1����ط.IY���u���
�F��Lʠ���4˭�2)���ᓧ�K�L����Xn�%���9�t�u��P�Eri ��A#J�ZT��:����2ᤁ��w'Y~S��e.nePۗ��f苇�g��������8�WG?W]I/˸���1KAY�ʮ�0��O٥Đ;fiY; ������YDM~���ٵ�J+�<��v�0�idi/dc�sk��k.b�1����i��<�Q��1�u�k�n#?L8�M��eO�Ό"W��b�)����O��5�_r�.(5���H����d��:;@��W�Kf7��v�cY/F6�~%���#۽����%]�-Ok|�W����@.+ɪ�����	�X��3ƣ���)ZцR���5*U��8�K�W8^�0<7N��m	�ˊ̳�Cdĵa��F��p�0�>���6��-R`�D\��:�I�rL��_'���xu��Q���֖�9>?��*4ϘOi����{n'�x=4-��R�Π&��\�GmE�� jbϣ����.��޺U�:�Џs����jVs/LR9j�6۬�k7��r�'AB@*Y-�(�X�O���H����>�n_�aW�y;
z��у��I��p1��i�T����n��˞�x2��w�8���TM�j$��<')��.�R�kjLʣ�1T씡��a	1w)=��RF�F�R��N�]h�e����B��"'y�K�Z�~��}���?T�s/�E5f��eۻ�&!��|�t\xS�:�|�h�T����%gfi	��	����5�)��\P���r'zF�:���e(���h�0�N���~��:�5��'�~'�$���`�P;ɟ�R��)��5�gI�vJ��,�����O-5;������18.. J�V��Ke�̩c咏c��w�˭��-�"��N�åf��l�*���j��w�!�Ry�(��$���vb�0���3m��qE���xZA��u&~�NŪ�pԶt�M������O�Z�x#:�:C����$YQ�h�ˉI�����T]8.�v�:��)w��ߔ	TcB�}�痹9����O�:_:�6 W��O�����?'sq@��v��d�	W����S�ճ�Z�G��f}v'R�Cw������~�~�q����R�ؓ���<�S�V7�q�Rl=�9�e��K�?,�8�T@�b�
ʯʣ%�m$>f�G*8��F@�1�-hv�h�sZ)� 2W�ɔ�Dx���6.�p�b�_�N-���(���~�K����r-�Fih�fYb�*���ʙۈ��9e��~]���HJ�Dpx��F������p`���8��>
Sߤ��8���]�Z�k�'�L���ͳ��/�Z�~�ŋx��P��>�!+Hw��ԨV�LM���%{<$Qlڊk����w�mF��$wd���Ǒ��CH{!�V(M�2��ϻ$MdV�ﶾ`�c~�a�҄ݟ��Gx���%T4�x���o0ԏ�3.�ZQ��4^�b�&%3,f���!o�`�2-a��rEƪ{VLs<W��]��9i���HɠJ`z�V�EH�?�'e�5���<��[����$�c7�cs'lR������có�oWl��`;�r��s>�ߊ�"K�������\Q�~ h�~��Q��l����V���\m���H<hs�Pt�שSE���ߘD�V��0��bP�S*��D�j�����=�T��SLa$i�����<��O�C��L�������4��>���ŭr������J�R�j�&E
�+�P����g�;8�RQ�O1�"�=JrBIFrW 4(�����s�+BW`�qo�^�1Ԝ"��i�Ј��E�^Yi5JYh�f#�i��Aw?/��vЬ��S��ѹ%jX�dzu�T�GrGD�b�L���OK�"�y�%���g�t������J���k��d�o;M�?��f�(�#��@��(�Z�%C�k��q�(��Ynx�
��M���e
�o�
�7�VAO��t)��5������Xq�0�3Z���Yt�Z�_T�/�[����^�^W^�8�?��M�v=-���|V����Zj4�_��4r*ū�à�K�*s/�!֞�A^�d���7~8I����arDf�}J�ˮ�gL.�RS�+E58FL~���j�29R�l1��;�?���'��X���i�'��P�\�� �QV��e*�e~!V��*���}IO%HS��0�%��5Y�D�4����[I�fњ��&vfm�,�NS+�L�����g���p��@�</GE�|��]�>2+0X!?�Z�H���FӪ�R����+�~'"��c*qf�y������Y�e���'��ڭ���#�v0��p�(��
��5�0�{���z�fD[����*3g�N���}��#K%b�5���R8"c�I���x/Hh/4H*u�e.^���2=���]ʥ�&\����[[_&��Ի�����[���E���S:�G��A9�n�����H�V��k�����~���E�<�����H�G��m�y2ޡ�vh���b�9�7��e��Y݈�η$ű�sߌ�rE���f)�*H@��Ga���]f�s3ٵ�b�u��,�B��=��Z�����^`�t��LK���su��â�R^��eq斂0�F�
0��>�
U~u�Y1�o����`�v�H�]���j�94�H����\1(ڂ�4t��n�!���/��ʋ�%��Fu�P���h�-���[�x��b��GȠ"�uE�<��I��;��|��A"���Su���R������U<����_Ğ�F�(	A2y����ᛴ��Gs+���|����zGz~�%��eP��l: �s]	66A��H��/rl*KS'����11�c�َN�2���t?t�m��=�70Ec��C�3w�!:��
�'�Z��g�ay'�x�\���F���>o�'?O����׌��Y���f�O̜�و�A~se����\�ɹ��f���
�qs�@R�:�f�E���U����\�j3����	0����f�d���%6ͱ�������Y|�^�ov�M��pJv���4�&](�Nٶm۶N�>e۶m۶��m۶��A���=ٱ2rE��j��@�M�c婲V0�}�~X��`]�����St�,��k�,�
*X��Q��4%��kK������C�,M����ʵ^����˯'o�)*�DU<�c�y6��D��r�h+]#��I��^����|��y��co���&A�<L3�7y�9�;��{Z\~� �X�2���񤱶JQ	���w=�L����!����K�^M��`C&��ٹ�
∫�1 �a���5b��Z�2�Z�bg�p��v��<��綻���U߮��σ��Ӽ�}έ/���s��ѯơ��;���� (
&^]AUW<�}��;��OJYAݢ��2�1J�m�Kzv9��q�)��ZH,{%����Jzh儒�_����`e���8�bj)�h ��L������;Fq��4���~�`�9Fn5����͚	��ڨݒ�M������/N|<J��=��Xzg�����`���9*����BVE��B���r�'w�(tz���xǾ���0�鹂��5mu̳���-���������J0��P�6嚏N�Ԃ�Pv��G��X����z'X��y��sv�'���\G��|%5�P\�_7���*��Bar�uh꓿�oT�Uv�h��?��0\�?�M���s�RN	�{ +��ܿ���6Cm~?4_�����e�yce��>�8�J�L\�_/
�w)v���6�K(Ϥ��b�̉�i��v�k�Y���U�8?R��\��1��׷cV2���T��Vʽ���V������+���㆞Ay��@�����b�[
�c��Eac�����J�����+4������B��ܺ.L�m:��6;sǚI⥴-7��=�kK�t�S�}nGOq߸���kM��Dna>�,��N�H�����OL�u��M���:,d�ޮ�v���FU��=�Kr+=Tޣ�����;5Uc�kO֩r�Xz��K8��Ns܌w}^G'T?�7.� y�8�*q��^'Es�QC�H���r�}��]�|aug�
~�p����՞���g؝��Z;q�>�(ckӨ�-Vj�J�mp�ָ�q=��MU��>��=ru㲞$!��@��� E���x
�G��	�u���	��	��B�̚�/���4yizյ���~��m}�z�z��x!����M�4�jY����j�
1x�gV�+��u����s��fh.g�C0{ �%��8�?��I�X;t�2�$�w�N-!N�꿾7�i���PZ|�܇��>��:��vG������9jz�&�f��U޼N���{��z�pbZH����w�p(6���z ��'���8Ҙ(�6�p�}q�G�֣��ށ�7��-kϮ�-@
�L��3v�>B �,vl$��s�� �\��,���=�m�6�����~���},|:W^�uI.`4�T�8\ޮE��S)%;K!��f�!�;0zz����� *�)��M�ׇo�b�+V��|��*�R�Z�DS��p��r/ѽ��VT9�8)��'p*�W8����t�f.��Jxα"#����|1��"�|V �3�̑�2D�G�?lV|>�|�,����%�����A|w���x��q�d!��.��6�Ow�YemR>Y��f;jT�7<�G	�OȄ���bj^/�m"��M=���s;�V�\[]U>y
���h�5�P��C�z����o�KR��9����a*p&�X���0qJS{7�"�����t4G�S�UΣ���	l\�]G�B63�b/μ5<�`P��vp ��C��	����W�67r���ڲܧ����Ǧ�*�ɲ�Z���*�����4������@S�3�������N�1����Q���u�Yo�� *���{e�}D��V���|�a�=7�<߷��I���XE��˗�d���]��I��������������l�J�8U+��&�X�}R�uDH��f��23+���k���0SM-��0Q���(��?�(���}X�eZ,V���@'�V�?����H�ꮨ*#e׃ESi�ˁ�5O;��<Q13�n7d�H��\EQ��0	.|�"{Q�5ʺk�ȼ�}�)k�,&vn-�_6��	RX���ѐ���j�����j�� �����-�����W�-�ǵj����(O��D�9a֌�I��}9̽�0��{�_zB,����[K��BYPv��q�=�@B9l��N�d�Z*G}N�F(Tkv��:���A> ����م��������7���1e��s��^�ݛ�����+��M���uf9&�N�7V�KGӜv�m�����h]�(e�}��$���+���nxS������օ ���T~��8o:ut>�:<a�@�9k�uۋ)]rp������D�XB��ŚׅSז��Bz�O&>-�/7�L����EMBS����!�[�e��8#9�m;�k���
Clh��5@�xO4A�S$w�KK�A�8AT�Q���L�Nt����/~�C���Ѣ����4�	g�~��
WM�!�7�%ْ�s4<\>5&���beM�\�V���e��~�Ibv
����c���� �Z���fDJ����]�}�	���T���5��I�q]v�ڛ�T()	کq��_�v=�����Ce��Z\9�v��tE�>�q���?��X��i9m�afz��taԥ�yC��x( �Sk�Ѵ�=Q�^� %,�I���.��1��46�-�<�����󐡡�s��QF���������KAG�N��xu�+���1��<m	}F��!t��]��H�pq�?B�}9t�����i�x�L��m"��^��'z\�A��pK�7��fD�̰�vk~G+th����2kAz�4vG ���(sG��k"����f��=I�LA[>r+�Ajf�H�2���f��n�ՉӦ������b&N^�&�4P��h�
qz<���b�n���	�*/{�E�gg�gE�2jN��b�r�&q:���䗝��)��Dl_�i(׋����`Ab�Ab0�R��q��iC��Ǽ�%��*a�?��T28腡!B�5l-�&sZ Btg
.����`�	#)�����x�}����k-啋���9���J�'{�q�/Av;*�%м_`V��# �`��D�O��f��z*{7f�(p�=N�+�,kk��C�5GF�vn~������P&����卧�T���t
@R,�E(9�` ��珀�PG�֌A��r$�e�(1!�:ꋡ|���AƉ��w��̀���>�F��ߝb,�g)�,��[���>��?*O���5�N��M�����ڞ����	2�G�������2g�%ȵ
h�M�%!ɤ$R
�}Re"��#���ÇŢ���4I�2G"T�lY`<A�)�)���֎�|}��
�oN������Bw�A4�~� ��(w������GO�O�4[���6��TXc���{�ɇ"'p:r}�������)l�A65�?Ʒ�v&�k$��9��a�4�6D������o�'+�������
J���#
$d9a<��凸?1#����/����b��fk���h:�DkU�O��/�n�&qV�8�bE��c��D���J���T-�"A �R��ڭs̮��EL��A�D]��
y�B謼���Ӵ+;=�7����9�{�ԉ�FȐ�4��fGJ4'�S2�,`ΈyT�^ \�6��L�;K4��0q"
�,0tW��|����s�Lɮp	mO�E�i��tr���%��������<A&�.�>Yۯ�Ŭ��D<�(ф��U�O/Y��R�$��q��Bvh����������y=u<��E!�5ާ�o*����.%�2R���vZ�^��Qt^�K~:��g�x��n}c�݁t!^��h"�,�+����S�hQ������j����9lv�|Oh�O醜L3f���`
����_@���_߁J��T9�D�����M%���u5Zi��i�I��n���5����|(Y����˅3�/����Ɯ1�'fi�Ac�-^fOvVG��������k���v ��__,��C�^{N�ȶ�F@ѕDi,��9-h_x%މc��f��ǉ_���M\���MJۼ� *�/8w�k���X�x����|�����9������i*��h����*��.��o-̝Ч�/��~����4�Wi#,wg-�������uL|����5�&a.�*�aHP� Mѿ͸_��՚@���MR�x�oQ��&�	�ӷ�]V���Sh���*`L'����ŗ��eO,%����@��y���Rl+����E��`bf�����]�K���+���� J.���cD�R�Τ�G�~2OB�|2 @�����{0šT2���:��&����0���Y�Z��s�5���zb���eQ3D1, �b�k���&(�����aJ�_o�_4�����J&w�m\0��J.�����
Ȩ�-U�1�k�� �s΄�Xb$�A�bk����� �&X��PT� -;v�gL'tp���#-(��*��sWqd��!3�.D�.s&bP��s��P��|�>�7��s�b	 �N�n�=���S�H�����zܧﳲ�<#��:�]>���*��px1�2�zr�q�dr/(Ū\����7P�n��T�X~�W�"���g�H(4C�d�X�% �g�^|٦bU��/I�K��y�_U%U��ߵr���� ~���0��S�O=��C���}'n��'g=��ԣ�nosr �Z��������'�@�<���l���W�`	��͑�0�9 h�6g9u�_Ĳ�G9�bL;H��#ͫ,�x�3�(Ӈ�F������k.�^^F��ҌP������Q�O��^�i��/���`�hO}�7�A�!�%�_=��W�r��Mu|�//A�R��mo������ԝ�7����&%��XK+K��l�A}`uōX\��	�A�tn��'(
 ��T��z�K�+�����?���e���R)�f�� �G�Es�+Ж(�M`��P��$��gJ�8ח%脱`&Ɏ�W�HQ���|6L������Pu��<���xx�k�ު*M'�$z͍n�����|��pv�s�v��TI��#;�c�7��S��Q��D���MEZ�a�$L���i��1�F(�X���CsC�d?$OoY&�p\�z1�b�긱crS8�{�|�54�Wvꤳ8���?��?�� C��%Zbwg"YZ[�#{��r�G����y1�e%�Z��v[��$aj�}�W��`�X��ʢ�e��*�?�����gD�]4������:��;<���;��m��@�~mb�E?�h��}��}�k`}���	0�{��Ea󊷤�J�n�җ��Z�B��8���{ A�[�: �AR8�!P�=�z�u}{���?�=��R�-Д�����#u��8Р]f����=8�������h�K�����V(�"��U3;b]������(ʔ/����gw��B��C[�/���>_�. �y���P��N�(�	V�{D�����S��N����)�U����~R�Y���o����1�ߌ9}HQ`F�.4��q#hGf�����������=0{��-��넊��tGc_��'p3(p���r�����y���Jq��	��>�7�
��i���Z���-x�J��A�o�u��FNa���f뗝<�R��*Q�L�i�u�uix�~8���X�D����B��*&s���Lc��_�>н��aGƫ�����cJ�Z�q�T��rTF�YZ�k�����Qᎍ��*$��}�Ǵ�����j��S���&�w{5kM,ѳ�wX�MX�J���	� �x���뻵Pz�r'����*"f��KG��FJ/Rk�����2f?%�|Gb��Ka�� qJ��=%jS�NO�c��yko.������8�'CvP�2�瓸�-�.Z!���Y�_�Z�A���X�<#{�6�����d'f�8�v|���bM�p&��
�̇f+-�p��Һ�|o��7�~���ӽ*2��z�*�K)�^�^�O�Y�;���=p���%�����t����6Z?��7x狭�^��� M���������"��ɒiY��!��j�~�+a,��
+���:	jq]'�b�3�[��BSs��q�?XOI��r�<�Rz9 ,��X��&6�B�I����zmC�8T�Ր0%|V��"I�x#ݺ�9,~OЌwQ�~-����6�X����IhSY]M�Dx�,z-M/�6և2C������-{N'"Fx��e��hD{��2��N��_K3�uZ3Ɔg.��b�'Wi>?lњM��T�t�}��*��|k�Ux�!���N�����]�'�C�+Ǌ[���B=��4����3D�>/i�k�&�k��?��Hs��%rEtFL8^����"��џ
��p��uE�U6��n��tU�e�W:�0q3t%(�𢖔��@b��p:ߠ=���|���>b�P���ڹzPr�b��I~0�]6�	k�tJt�1>vT���]g� "A��dw:�0�cgh$&KI[�����tfx��,ܳ�fS-#��6,=���+C�X�%���A�;Mc�c��(V��jhQ�h���>���pZ�����p�Cb��O����d�&T�&p�jF�t}ye,@V}a���f�Jn�@A��	���1���
'��&٢��I�pTRY��0ij��Z���r�Q`�0�fӕ(���ӂ!����5�E �5(��Z(B�Sb.�@&5-{XXB��á��7T����jF�m���k����/2�Ta4�.�~�n'���z���)����~e��}�Q�Ņ�|AY���G%�UR�jR��p��ۃ7�rg���Fý5=]��-6�2l�۰���'f�d��Cʺ�J���r��$i��5E%��U5XM;�S+A�1���\Ȕ�j0��`���lbݚ�wd������X!�h���K6]I��	Q�R� �3�r��'���xZXׇ�5(>��l��J�JW�����g���^�x@��*�J����D�p��n����w�����Rv��;wy�ǹd��V���g]&�Z~��8���s�_v=/���:^L��ѯC�<U��9� �b�l�Ԙ�6
��~O��L�Owm��m��
�ѝ/:=��Q�[��Q���$��,(�a>������T��AŜ�"-�́G�1{H�@k���'G����]�N+������!vG���T��[�-DC��6Zzj��{	w�M@oכ^�q��d9�������1�Jk�{;-������I��H�Q!'z�i %���-�&��m7�p��r'���0�l��K�	��^;Q���g�u(���v"��Pj�]k��/��5�N�ĦIń5�J6���l�70������b}���Pi�O4`��`t�Fc[��6�73>��s�����`�!I�^�:��}���m�M��k
ʛ�)���#�seϔ/��<��5*�H�N�WZ%����=*�bc_���ܟ��l��F<��MrxC����)�cFjA�(p#��s>�7_5��ZW���p�.q�_4g��<���|�|���� d��b�J��(�)�$;�A�;����Sɯ��?�-�/�H�����NT����WmxO�`{��K�#�D�1�!	��l�r\2�\���Ӊ���s�B���Z�����u�D>�x��^d&.��i<�$�۔�$Zכ!
�HB����@Si!3�@MҖ�?A(lu�/��e\���.�]0GaV�-|�gx�J��6�af�(�?V޺���}�?���w�5�4g��}�E��ۙ���']h}QH1����ԂTf	���A��:�IPD�}�KX�պ!�^KfK����?�|�iQae�������TW[x<�ؑ�#�E�o\c��>�{$%=���4��>>��9Mݳ�Ҥl�[.�7*S��+.إe�}7��;_���he4ii��;��"Rc$Q�ÿ�S�5�hu��a*�a����hO0��Q���Qa���e9�ܝ]��V��9�Xʥ�.�����/��$����5�O�Iu*��H�xA��L��bgh(�� ��.�e~NL%�H�R�kY�984�wa�Ox<�����#��V�6��yrkN�Q��9���u9��ܒ
�Ju}��-6�`���IN%��M�����8�*������r�����@���sW�?�F���P�u�E�RAƪʴ���	
��@2�<=�@���2�Ԡd1��7N��D����Z��8&���l�rg��`��p�ϧ��,TOo�����e&�as>�6 ��'j�\��%�s���,`8g,�e¤�6�p~%��8��k��GY�.���\���^9t�̈́�l:;vM����ߔ(8�T����������R��g�؉�� �����㤹M"��0��K��U$�X`�;�K���vZ�ug�M:�Ix�L�V��(#,13j����T�P�t�Jc�6����r*��oޞ�h�y��vm��g�_i�4��~�׿~M��s�G�<���xS)>Z�fBL�+G�
P�2�ew�d��*�{_�7[�I��k���R�e��/A��Ĳg��(|e��v2�Q�P����Xcl�*��ISr-ɼ���Fz}U>$
R��UçD���`��6b�ʍ E�#9m�x����Vd٣~�L`��YS�%\����==�|�LG�<.�*�Gb�ml��҆�E>�WЬ��hl{��Me�H�]�~�E��X��؀n��%N�����B�z&�?���k��]�`�Z��ٛ��i�"��o���Qʈ��ٛ#s|��.y�L�C`:����M��Vu���z�	�~�S�5-�FzW�Q*ı��Cӻ�H6(�����^��Kˬჸ����@����O�z�]h��L�R�f�^�`=��T�O��Tg���Fu��dZ�����%�}8.�h����c�X��&�����17[m$j�a���^z�p���+����Ǣ�T\��v�Ｚ���n��y)C���Ds��O��YM`L��=,я�ڦ��ͬ���i$��#�V�Y�_t�6���r\rfw{CE;����ɵ��S$������͇�:ˤх��&���:cSuY�t��u�ɲ������"�/K�.���PK`�VT! E�h���dB��r�0&:eC���Bv4�#�"u�<�/�K[�:a�{B)�A��3�Lj��"q0�� ���J��ΌD��ҁ���޾��(�1<:@Ѕ�׶������Դ5����?�������%�������b�e����K��_��G� ͏P�J̀Ӂ#nm�$���z�J;�*w~���V���9~F�vc�U�XQi 9���T��,�����|{�/r�y�e��U� ^��B_/ʻ��p�,��(go)���k�9��0�.S�D�dgo�q��B�I��q9��.��2�ێm�*����y�Ĳ���4��i �*�Ί�����o�VTS�꺢��c^]�v��~B�R~�xK��yc���gJ#1���J?X�C��(s͏�\>���n�2ڻ�����R(��>��;R�d�~_�V�g���ulQ�����H�׍9�ƀ!��o�'{��>�kg����LC>�&��^P�i��1��	n<�Z�Y
�㟦���6�~�o��6���4��V[HL�v���҂�b�慅n�&�� � y��v�I�:=PN�����!#�zsT�E+$!�l�C��4�	�w�D��va\��ⵅƵE�	bD�+�׎�Q@dƽ��w�N����� �
��=�%M8x�A!��� ["�@�y�Ǎv})d�}+�#J Si2`m|�3;���eObGR&��-^�1m��j���{��}3=�>k"��TN�\+�ny?�1b�v����+���N�:4g��~jW�C��9e��E����?�сzR�>�a$����K�S���,�D��j&�y��h#P�8I����bx|Uv�~ԃt6�WA��a�C&�-�p��>�#���7hi3[qx������}��-ٝh���V����yQ�[o?D��7a� ¿/6������Cm�	)�柝�VCJ��O��&���`=��gʜ�&�Z�}tw�?""�P��X#׸H^�>�Jn�'�Y�g�*������	��5��)q�õo�C���|����Z]�Ht�b?J�?�U6d�ϴ�k�#��Gȡ��jr���u�L�����AEu��XYA�̌�2�Hʘ�C_@�T�����n�`+t���J�?�D��
/����I��MY�4�sh"��)��(�	i�����*���K'A��UС�P�ensw�&��F�ͫ�N�!<�@����uK���r5&�'��4���c�Es���6=lgG��Bx��R��6��v�~h�W�֚�g�X&+ᣛs�����BsÇ�"���%o���8"'bbC���zcm%��%�B�<aդ^���]��T|��~ވ;Hl*%ģ+���r�G��(v�f���j�(	�S����A���t��6��}{W(�����=xQnZ�!��**��~�uXn:����?���M �z��&�yV��[$�:�hR���Nc�.M�W�_�@�Su!2_�*19��(�������W{�x����D!���}a��<�>��8,���������C�T+��E�}������ֶ�hJ��@b��ʌ</o3����K�1�t��O��E�*4�P���	E��
�\�>�D���!�������br?X��m��I�����q�c��-AC�),�\�����
�#���v�O�����A�����z�m�n�E��٭"���ܶ"	r��H�!��xވ���1 �߁)	�o���B����9Ef�0�>�v��u�`�`x ��W^\�,*�������
���u���V2���hU 8�ቃ���(��x)&�д��(l�t�F+�b�>��eP����^pq���2N���2����7|��<�i��6��9��7�20������U��6��ۋ��z3�V/�ŋ<{~k�?C����'��2�������L<����{>.�B@ʆH��̻zIJO��Yo�{Q��䆳�T��r{�$Ǿ]��5d�=/A0��VwX\R�l?}yi?�1���qaY9�G�������{B�����d��X*��9]Z
�ı�.o�봛���T5��!F�/k�~��R�����$���@v��E��-���9�&���wشj�h�>��T�M	�K>�s��/�U�+��!	��u���5�j��\ۃ���`i�2�n3=����Z�g��B���Duͯ����\.3*���=s@���\iǠ��,� �<��S&ɞK�O8���,Ң,� Pn09�pJ=L��A��j������
mLﲇ��8������r>L�_Y7+,:���h�x}�ƌ!��m�{������B���e,��������4q�wǾ�v�y�h��U��'�B~G�}�uJ��M��bw"J�)���hW�+�Syy1�.��hdȑ�Ѡ��*�T:�4Ja�ͺ��z��T��Tn*É=n2C�w
��}�]nG���u�f�sw�0�������0w�oPyC��~��榫���]���·�틇��M��~��~�uY�Lܠ�Th�>{�3^j�qu�I�t��H!�[��;��9��<o.wH~�?����n+�1^����8�)�.�TFCw��M��K#�ad��[	�w�Ky�C�翗H���� ���B�kq
�K{�쭃�}�m�R(/���)���������m��q=�0��������h�my��p"W��
��~yL�6�w��l{1:|q��-ɼ4�Q����J��D`��W�	]�M�A�ّ3-�����>M8vIa*������,m7��<��"����{��	�l���No�v��ij�WN3��MwVVs;�若rMRf�^�^��[��6��;�۟�$X2E��r11�VV"�Giiꔠ�_?o�(U���ڢb��Wl���-m��&&��Ф��%e"s��;�|�V��[�U�c��bnx�
�1�q���u�?�ˋe�~z��ߊf��u@�~18��/+�C���� o�<^|�o>ss��
���Y��e
���	:ca�5�
΅����[t�#�X��ul���>�E��B�ЯM��iG�xq0r�pr���v���D�����u�E�w���ݠ��Xe�arl�h�i�����p��Ju&F�h��71�N�� ]ȏ�1,th20.e!j���>s^
0������-�>�A�o{��)B|��q��K����7>�O>L�^��$[��Hb��B!dC��"��m4�sc��PUƹ�E�3$��0�!f1Q��!�c�9ݍ13����]�ː�C��rBm�wnٍ�k�ڰ��g�*���J��h��
��]`�ڠ�s��I���RiI�de���m��q_���у��oׂ̿�]{u#�YwS�����dR��k�#X,�����;��>Pw)Ԓ܁��8�������Ck����K���\�O{���!
� �]�F��`�߀��p{�P�<�W�;	�~ֶ��Cqu�ʪ�BP��kq9���>�gL�V�O�[@oO�ߌ�T�6���^�'�sK X7���r�ǋ����`�9�?�#�!�[M�q��Zh(��F^t��I�F/Ѯooǅ�,V�ۡd� Ry/�7����JKF������Qp����,Y���ڮ���s����gI
�t~���T!B�:�I������OdOq����2/��0���Zs���g�W�{����Ξ�8�t�oi����t��#uƔ�������e�u����j;�������B��&ӹa�p@)���]\.�P�,A�?N?߁W���*��x0�n��8zX�"������� �#����U���d�\�☵����A
5���)��P��`܎f�bK1�-�i*5�nku����NǸc<1i�ٷ�#��Q���%����7�؈��R��Cq�����Lܙ��qK	��c�4g�l����
SP��5U��Ś�0��~m��E��2N�fja�;*�IGO��0>pSo鵆S��"���4̣����2!�}ܕL�|�i��"x�-bF���|ށ��}���G�4�ڜ �ۃ�,�φzE�s������@��~�ߩ��h|,�n��Ns,O7��IV���c�y�?F��*.��:��`	�{w(�Qt'�Ltk����s>-]�0�Z-��:H����U�>$Zf�������r:�����!�X�rv��f*Ó��LM:6G�]����'�_��ǻ]�������@��m���/=�K҈&��mx\����-�`�e�\�/!JM�M�.Ə��N[�>_�F���Q��f��X�ܺmч`��t���8��h�����۝0TJ���4Q��6
!<�l��P>��v��S�бp�&�5ɟ�Wj�~���SW�d�/c�(E0��n�4u��ʓʶ��*0�����V�yߏ�ڿ8?��������-�{x��PO�� )��!kO�i��h+��%�1-S��l�s3ߐ(!����_�2��Dvd4��u7wIl
U�z�٩\Vp��h��;ȕ����"Q�C�Ϳq~]�2�b��RŌ�x<j:��3��A�����Q��CC��{0+�)lYw���J�Ě�Q���pl�rcۍ�;�������
g���L�b-���޴���-ዩ�����VEey~r�"a���C(E�Gi��p��ੴ�O������\��#�0{�����>��&+�r���a�����س�=&Bf�q���:��ʬ�l��*%�b0f4�?��	�*`>M�O��h��8�ҥ��	B�9´�h�x���GǾ��b'l�=�`�~�Lӊ��(��r]�����e�H={[I��iu5������]*�����]���?~�p��s� �:>g`n�]d��!���C;��H�ςF�fI:�Bwn^#;%�'QL�H1cP��+�fRL�N������FaB�)�v@�8���.Pj�̡�i
��!��i��⊺�AwFϝ��m����Gyf����Y�7�!}Ӆ~�$O(�E��[�n�����C�w�OS�\(��B;�Q�u���%q�OZ ���$ԇ�L!�8��[�3G�i��� �=�P_!�R�c� �~��?�ფӏ�=
��m^FA�%<��{Ѷ>͖�p04�JԠ]��w�EZZf/�+����"��K�\�%�(��F����h�覆�7��A���%��G��fӽ��;�&2����ړ��^�8�eu�2�c�ZOti�w
���is���`�������!{oc����
���G�aC���SZ6D�nT�f�ϝb��mϭ����\��a�eh$~��
8�=��`X���p=`Fh�K�ȉ0R#ב���ԽTV�ƫ�q8Lc�:P���OFu2��o� D�������@ ��[�������s+h`�������`0M'xdē	���J7j��0g
�y�j�x���".r�u��>��zԜ8�L��0PeD8�"ڔ/rk���5��T���0y�������dP�]g�,I�,1|X<d��dC���ˁX�۶AE1袒[E}U��?�`MZ�0����됑V��0/�����w������>(:���}�����]�;������E
���b���Ѿ�9�����^��r.�&Ը����<c�8�qxӮ�	/,���.ӊ��	#��K�'L��f�ꟾn��	��@�.Ǹ�~�W�t�Γ"y���bg�3�;��i��E���Kc�6.�r�KM�2|�������n6篪���{Ne���"��^����и�=j��t��7��o�w3�P�m���^B]+��Kt��v �����h����K���=	��X{B(�u�7F���h��E*���$C��8�'�#H��-Ƚ�m=f9ܿS�Y0�k;k��k��- :��	�]���ۥ��fڄ����+\aU�D)�������}� 5;t��m�l^Ic��b����[��8rGjQ�*[9%=�ϓ%�K�*&t�h������4k\�?Vٌ`�
� �����djjJ,.�h�T��(�lr��#�v��E)�n��^5x�Day�(P���7�t6ޛ�k$�3Q���ULX�A�ޣa�\{�E��a�\�lv��*��Vp��S8Z�ώP�1�4��4\��-��Gh�oұ�_��+�&������z�w��n�	Ju�FyϋuUFXȂ`��v���F����P���#����Z��x����H�E���K*L_��۾$l�;6�$��'�`)�&Lj�мJ(j�G�c��]�86e�@�d����ho�][��9)I���3��"f ��$���ߌj^7k�v�æ�ٓ9����V���t��ݭ�E�pe�\�=��Ob�o$,�߷�L����>�3@}}�~�tQ��d�{-{��i�2�P\�`�E���ޟ��Mk�j��`���.$14��*�I�w C���)��v�妼�	内E��&5�B>��x�Z�P��[5����V����>�l�e��Rds�0v������Q�g��� ��(b�]���:yp%ށ=��a#�����~h1�p."?��j5`�VU�%�)���p��ތ7��X�rk�(����XL t�K;-�r��v;��9-�B#e���a���G�n{i�E���V}���5�tB輸�� �K�~>0T��=���V���:����&�:h�>��!8����1�qK?y:���x��K(���b��q����.9�%uO���HK.��(��QC�+7��`��_%ح��hq��G�ޱ̄��4:.\x��0#L�����c�o��x�-��P��Œ��$����"홹� �d{.�-���q���b�؂�J�	PaG���hG����U|�7���{K2��\�����ցRV�����$��x43|�l[�M�H,l�g5��ji��TI:���b�H�s䭓���/])�0SG������~fVz$Lb3�<�3d�y4s�e� �x��&/C��rO�g-�;��[F��i���@;���~e�=T��&�,�+�	GaǱm2e��';�	P�qA� I@��6��
\�G�T4QSU-aI�tN4��}�$S��c��cSd�����_��׋p4�ڦ&,8q��E��x�8<���I����u�_�f��t�����8V��W���s�{qW��[�y��=��J�c!*�k��t��Ÿl�"�����&� �6�%����Y���!<4(2���F����4���ĕl�ҥX�fN\r
��ぇ�C�>�\YC*Uj�0~�Lċ9X*w���*0T���߹_&**�u�����!-eMH��,�SAM��_��6�a9 ;�����;[vч;���>^�����*DG��mw�Q�2�;4��q�q�2���Eic}L��J��ۃ	��cppP�\8���,Y~�Z�2^߲Gbi�O��@c3b��{QIҁ��H2(n��~pڤ[�S��q����o��Ώ\&�#��Vt�����:�N��d�\�P5�8���Cg�9)�*͛=��ꗈ����O���!1�پ}� -������"PU��^z}e�ь�mi�%�w�;��z��:q�BQa�A	%k�e�[p��p�L'�v���3b.�P�VL��vrb9����1�!���#�ڌ�_yQ�I���q#_,���e�120 �ǁ���s�/��;��'V���N�YUoMH�J��h�R�#�X������p�R�ǣ�����έ
��h�ʜxK
��,s��L�@�EΆ�kE��U����	Ye�lR1�|v;��� �ȡ�8e���>�u3���-(2�3�W�k�+"���^�O]}	6���d�D5UU�������Ng%>���ѷAu�����TN�C�F�GC���2�&"���Y���އ�T=Q�}��+���o������|�����?�m+�����>���n��O���'�X�͜�,�[��q��p�I�`�l8rIx�U!�����z:�h��au��	[sNm:	W��],J��k0k�	��}c�;[�6�����^[��sf��"Ӛ���͸���R�CPi�n���d%�]s;%��v����7��0���_|&<�2�B���k��v�h��$��q��o����C�����LڜZ	���.�&͙}b���x�2�dpxX���5m�z�x��nv�F<��L�m�klB:�F�@�D�h ��2�݌��jjk��������(x�kk�1c�NU4᜾�F�]w8����kkd�<|�(BES]-���c��U08�9e��,A"���n�.��ۏ]�;��H0<�86{ԟ���PES=Zg��d��ؓ���TY)K���јq14�T�t��a�d�MxۋB&�㦌��gF);�w6����a��"T�^P�n�ɤyq��P�ڊlIő���<�ʛx�m�x<ȗL!tFz�`�S��ٝs}#fJj:�	���I���N�}�ҧ!W�Y�S@d�+�#a��y*lGD)�F��M�� &\nr1(�P$Z���LQ�$�dP�=����H��ݠU��╬}#�s�=���b�ܺ	�p?R�&O� ��|Av�5�u�����]��Cm;!�L�����TW�d}M$Q�ЂP�x��X�� :�Y�@�y���k~}ݱ��>9���q���ݗ����20����w(uIc4e�⥶ƏR%�+/^��N����aY���l�UB�L�J'�(�F��<�����+�/�;'��p',8O<�^|�MD8af-8��u8p�u����'��͠j�̲	���N�y��%�2�4��TO�e%�}j5<n/P1���]��U-;�Ԫ����ΝA1��{`Ä� �	��D��O�І�� �z���d��%��0�b6��(q�加��$J�yE��h��4޺:�YDwu ,�&�k�飝�ۇb>-���*��߿mc�e�p���CwG��Y���u�x�(&r��OgsBLK�b��I��f�P[����y�\N٩z�x�9ĉ��%E��I
�FQC:SD���V���'��e0���܈�Y30Z�$o��;v{�+c�4 ���؉��YJ��%����#y��т��pM��3�4���C�a"<�#�h�D���1�Υ�X8o�Ǎ�����͕�C}QD3
�Y�/��e�ӀI�HT��bE�ʹkf�XR�a��n�H�P�`�ъE
u���hʠ*S3�?����kv��n��uN�\o�sl�u�F<^?
&-�5�S�9����T:�)p{|�����(�}
I\z�9��5����w� �Q%�lo �Y3g� �)es9�o6�_PR���p��>�n�{R�,<U5�3EWֽہΑ����ȧ?r�5�~�Ŀ�N�c����
��s��g�ᭃm߽��g���gw�{��1�P�">}�X4�	����h���7�:x(
���\�dZ$����;j��
7�	��r��r�EV�v�[x�U�Ĩ��P�߇����2md0)WX[�p������ �x���6S�\.�l��箿	��c�4�u*p�.�3���ڻ�̈�k:�����f��/>?T�^�~�f�w9t�mm��]tL�_��t ��éj�g�k��(3.�K}�M3gBP)X�q ��!p�8ͅJ��a7�l��6�9,?�46T#c۶ȧ�oM��xp��t�lK�b�n�P+.��L����o}��B2���=6��4��*��e�Fi�C&������������T�-�Q��[F��gWt&�'g��^�0�z�*5�;x��G���}���-Z����Z��gA{�S��x{��104�Ӌ�/����0qb;�<�>C[��[{���uxw�a�������X���P-jV����Ye�R^�n�Aơ:+Ph��T$+��xr�s��X���2�V��Q��o�y� _�d��=�^���H'Ȓ�r��
��[(�917b4��5�^���tP.[B>9��/\�O|�l߲^���i N��i����$�D>�G&�E&�E��hX��ih;U>6��:"�C���ة�}�m������q$�GO4��>|�+>y����>;ʎ����+p���_^��_,���ꊊ��l�/?�{oeWy�_ۏ�3L� $@B Hq+�K--ŋk�S(�`!H �3�X�]�����g��]�����[(�ۜ�fM2s�}�~�s�%4�ym}ˤ���s=��Y<�L�j
�%yl�r�Eg`vM|=m(��e.s"Ag{
��9��U�����<U'---��ˇ/��diE9v��Ũ���
������$H�"�U�j�p�I�c�1���2s��Z��x�7�Ձ\����C�o�cƏ��e�
��c��.���� �r�"�y
������E���IN��5C-a�9ô9SIf2�-L�+��SI��*W�l�ʔl�-Eӱ8o�$�Ie"J3r�� ���I���&$B17�AN)�L��<3l+���(�ő�OIY.J�������؄H���F�W��*�6itӃ�u�\uL&�ӈ���e����L�f�2�a��dG�>
`�BF�s�@Ȃ�A��dQIHF�!�hr-<�$x����;%���(�S����#���2��	��	���)`Q�s�T�g)xn��>���y���k��>��M�A:�^~$
�sz0v�xX������͸��G1����j63���@�D�W��}�MB�0����s�B�1�{Q�:�N�yKǒ�٠*��4a)()�{�s����D��P��������e!�(t�J(M�n�<e&��,ēT��P�g/�lފD*͔L6ꋥ�s&#>�p̡8��x�ŧPP�D&��L��R̙���Q�^z����H&tNr��\.Ģa|����V!�H8�B^�XH�Bl�ڄ��<Q)�v�A���?�n��Ͼ��������K=�l���1�L���%��J��B)KZN�do�FԺ���G�[s]G���3�o��ɰ�Iw=�3O=s'V �p0�F[�����mT%��������EaR4��Vt�u"����#�w֌���o����R1�h8��F�eg;�p�Q^Q̳�p4�~��@ZJFQv��i�޽Ml�rί�ű'�����_m܉+.��Q�|���-Q��lH�S\�S;�t�I~�4FR���y�K �L,	��{)@�S�)��)�� �HA���D����H�7�b��H ��b����,�z {7��� ���f.Q�(H��G]B�J��g�yݱc"�$��pL���2@�"�*�E��;"�Mjw$tC<cFGӌ�|�3���Y��b� 2E��W�u$R)��1d���$8e6��H�4��Y��4��œ'�M I�22X��>๯ĭq�g����I�K&�3c=��T��[dL�\�K.8���A��
I1c��=ز}���"/;����ˎ8���݁6�h�m�<ɖ���p1�� ���l�B�DR�"\j&�l�
���#b;�h��@@?Y64�%�Q�|����)�.}O��!܅�2΂*�x2�M�O M���"\t��P;^_�G[���M7��쁿S�0����Ų�⸣���<���5�>TVT�eK�͐ޗ��A�dJb�	'�"�����~�N8h��;�AA�x����77`GK:�ð9,�g���9�>P�?�K���p_@�y]��v4������b���$)�r����p����i�B�,��+IR]�}�L��ƞ�XV����d�JU
�%�VRȄ���(�����@����6qڴF�g	)2O�>��9�Cp:����d�Oe�S{� �)j2�J�8�;�c�"OQ�2}�l.������~�>��w���(f�4���_�n�դ�[�v��X�s�H�yӣ�3�X��M�"Y�I�2M���<�Ƹ����T3��B3i��t�7�"H�f��nadrA��&Ma�`,���R�b9Ɛ�l��=��ݍ0�ׅU�$�0T�Q-k�Yy:fΚ�b2�=�4�l�ٙ�x<��pO�hR%T��QRZ���r���[�3�:�v�Q!��f�p�	�b��!�doKUj����o�z�9|��fȪ�͚��O<����y7��"c����=�8�މJHk��>�qE#	�ᴃ5�y�N0�L�$��I@p��\ϳE0��47}��k��a'Eل��v��d{^V.��+���D,C,�h2!%�ؾ��>�$��1$t2.��넻 �!�iiQ�(���,%!�#�1�0!�f����3C M],dx�M	��>�J���e���>	���F��aw!� �q"a"��d��ÏDII5�����`篼�`���H���[������9������0��G_�Zw�!�q�K�%8̝-Bד��sN�~�V��O>^�TM��;��[V��3���v�{8B��s�	�~��9s>�o����ØO�����r��_�������{<�L&�lY��srrb^�Oonn�Τ���f�MU±0πE͊X���c�f�I�7'm�$MF8���Ȑ2�4kNĹ�H�#mX��F�7mZ�ZE�]�4R��ۏ���v6�������!#,�u���bpV:M�8�T�� B�xMm�����ک�r&�ʆ�z������h�ێ�/�
�n8]v�q��9c�A�!P�t����&<�̳����f��	58�Xt���$���x�U����y�͢�#�c��Y�XF:ܯ��>>]�%Ӌ�4t�T��)�&����;
��̂hQ��[�u�o�~��d#��8���4�_~0�?�Htww�l����/���{�#��ꐪ�L"�������eK`q���ra��v��Fܵ���1��Y9Ҹ�Ow☣g��L*�9$lP_߅��#����2,]:�˺�w7��w>4;PVʴ57���^�'GF�E,�4"�d"-���Z;��*Q����ePq�c��� ;ۄ;n�r*�c�,�����)�5��4�ɖ7�P,
4W^vԷ��V!L��0uiT����)� ޸�q`6Y��ALE�#�$hHA&�=Ͷ���,+Q &�A�4��4A^� ʻ��S�:
�3:EQ����Z&�b�N��;�`sr����ݛn��ո�ʫ�wo;Մd��&�Ų%�p�1K����X#�lV����.8�`�P��M4�{�@����8� ��`���d�]k�3�:z�=p�"������W�,�_|Ɗ3�?k���?�U���������'�_t���+������x<�P�TK8��	qb�u��9��F�eV.VF��(B�@n$�B�ͣ�;������3���̾͢��P�ܚ�(2�!���,)aQ202&�p� �w,ˈ���E����JW˖.g�ԋ/���N>v�I�h��i�^
�7�ܜ,<|����0ƨ�-"HOS �	�������_�%�,�I������9��賎0�;p㭷cG�.�|ʱ�\;q��+���
�������Y� qP����$����ē�F$�E�@'�AK��c��㫍[�H
�����E){�ǰ��XyΩ�d�ǰۃܼ"�7u�U� �W9�3kj�[5�&����Ǹ�!�E奰�lضm'�x��#Q�P��`s�x��?b����}�YFuE!ƌ)��f�;�CWG~}���u����Q<x�S�� rQ1����O�,4���<U��щ�-����:E�Z+t�L���X��{ �t�)�؄DT4����<d���l��bFqi	�9�x8����K���y/W�DM4�������MQ�L�}ѰQe�p����B�قt4�h8�z&C&�geD9�`�;%g�\K �Hq�JtMZ�4:!�8��)���L߹3DM����'9U�q��q!=�����u�,�	�P��X�.�r�]((*Ư���{;!��@�`�[_*��'�#�,�'��k���T��&O��    IDAT��y���DSc.�$2E������� Or�ݝ��f×L�{��Fɘ���U�ٷ�c0�`(�v���s�y�_v�_�m���e_@�_~�_�V�ԤT&~}*�8(�N�$.A�VT1K��D"EyS�͆��i��6��Ha�烲́�np��F0'lF�R�7��z.ϣS͉�J�̄Kb�4��3���F�jw�V4�!�.�zD��<>[�)<?�=�D����}�Y�g0���=;�Xy��YNsά����߳ʘ/����fd�碼���l�4�=�4�م8g�ha�6D=}�w������t���۟�O�݋{�&IG���d�brB1����/��k���q�Bռ���e�põWaт���nAOw+W�����֏��}�hn����n5#������@��=�'"d9ňDu�rǽH
f�7�A�m���!�}�	8���ņ���aɲ3g��Uw�vz��Ft�/�K/ݏY����e��v&<=�X�p6x�6Vki��}
��1r�S(�U/���B
f��������&FZ��j pܨ�Q
�y3֍��5H=90���F�W��)�ͥ��Z�E�*����3�!�̈́�N<E5�M�W�Boklv'4����9�S�d()�5L_U�`Ӡ�!7;J4���DH�_1Z�1��CNSW��c�q����$'��j_3X.�f�uiRz�[�ܩ����3��1��:B�R��]��&LbƆ����#�����^rZ[�A=$�D@L�"#�/O>'�8���(u�iEE�L�2��%(,.D(�c%�%S--Y|�������wؽ��:�1��[���������� z�s{N;nɹ��<�۟�6���~����J�����S=ݩ(�i�,ݚI'Sf���.�7ͥ%�/�e�Qړ!zAɑ�\i�v���S	cS�Fd���F[��b�W�F@7�R�נV)�ãA�~N� �jH�d�I�O�������kر��8�D��6o��>�Sf�B\���ه�~}�^�TV�ח^�2����x��'�uz�98��_2��?Cc� Xzڻ���[�#��,I���;Q^��֭�x��U��o.�����lau/�3{�;��ë0썲?96B:�<�ă�o�D�ؾ	�}e�\��=m��{8	���2���B&���O���v�C�:0f�$x�Q<��S����ao' X���i�u�q8d�ll��-K�����kh��p���c�g�R��z1�K�k�݋�����q�/�AC�n̞=O��Yy.l�݅�W^���"<��*x�շ�?�(6��([w,A1A'�'�I�g��������v�� ��Ψz��>��v�4DJ&i�+�����*w��Hr��7�ӆt<	ok���vc4?�L����$�B��]άAp�a�u�r�FR�D�܈�}�(B�+
�f�8�R����"6��y���Z�T��e���4f��Mz��`�Za�,��#�� ҝ����x�ŗ�����dL�
������t���P̄n1F#���I'���'��V��{�_��d�u��ɘ<e'c�,�8#��>��d|oo+��j<C̯'�	��_x�2������vv��{�؊��|ة�ZY�/߼��������r��ao:00P�+�ptL��b�8��L�����S�:��1QP���h0��@?�-x��P�<e���J~D<��Qi��C2����L�{
ܪч���~OH\c�n_�sY�"уwp��$��Sg��y/|� ���i�ۛ����k��B���/� ��V`۶-X��3�q����UW���<|�q3�|e5̮%ba�X,�6�? c����7���ﾃ��|?�}�vv0K�W�����ē��mͭ^2+��=�������VD�>����� l�k�ͷއ��!�ض�bIN��{n�'�M{�����çϜ����񧇰�����Ѵ =�Uq�i���c��P/lv���ޕ[���x�z�����IK��Gn���S��a W\~5��r�y8���ڀ��u�J ��_�yU%2^~k~}�=��57��R�R:҂�T�p�#x���"���y:�~J#�0�*^�a�?4�ОzH)�B���p5N�	x<�����ӎ��r��t{1X�D�u.�nh]�L�<p�D����+.,��� YLz���E��&�P �h5!ˬ�!�Ȳ�X�NӬ@sq��q�aQk�G������2 �?h�mA���2B��
���@�G��ѿ8	�& Jf<���7n�/��xFB�>��D�vhRq�N8�p�q�
�����<���p� �
r

Q]3�g腅��r��O��3$�Om�{��܄T��3�x.��Zg�8<���;�`(�����W�}�/oXV��?lk�_�q����ݵk��d:y���gi��9U�+M�eB���6ـ�T��"����)뀇IM�dLք�͔Z�4�Sxޗ��AxD��e)ylT�B�fG��F��G�����Q���9�hǀT��A<^������_��m;q��娝6{;;ˤP5���nڂg_�b�UTp��c|e	>��|�a=,�	�:���d,�Ŗ=x�W�	UOU�������EE���~`��b���_r>&������sV
��Nç_lŝ�<�&)�-m,LcQ%丬���c���ֶD�d��t,Z�p͵Dg�0��� �v!�뮾+�;-��<���3�Aig�	"I�����,VH��9� �|͕��G��'�&l�݀/���'��O�L�wȸ��_a��Z��lj�d���1P�2z�|��	��y.��뮾�k����_��^@Ls %�МY �S:��QUI�7�YH�H�@p2��stj��~9)ő縅8��nD��bI 7�d%�E{c�0��d�,
�U�%�Ϗ����$�1�xB� O��4I�k_�yk�0�Q���-�� �����!��QU���.+� ;���D�h��Z�R���_'l�9k����J*�	%ȢB����BX�}|fG.��8􌀂�<�"H�d�A�,U)Y)��� N>v9N8�P�}w5d� �������B24 y2L�#��Y�+=�B$F����lb;b�z�_�ش9EE8���X���W֡�?_R��fj���cN����-?�mpߡ��3�/�����S?u��_���(^�iʑf�Y`��d�8�I�;�-w��F�8UQ�o
�D�jhl� NA��5+++y�Gxæ��(�mt#�]��p#(摀o��iNO��F@7�ˍ��0�=��O�:�Q��C�re��^Eݶ�X~�Q�_��u� �2*'��%?}�	O���$J��p�y�b�ɵ�����E,GUY)\�y�^x�m|��&؜���\r�B~�b��J���;��--�p�2�\0EVN1�E��Y![�ع�?�$�Չ.G~�$�Y^����8�&T0���$~{a��;�֠�kO�}�I�YNጓ���y3�)�d�$�Q00��E����Ð-v>�Y6���K�?;6o$$�!�K�k��c����Va �@Z�`����S1mLt����0Y�C0��W�o���8�e�q\y�9�US��֭ǣ�|
8���#��� z����kK���w#0Sw���ҐTv���=�44@��=t���������	49�h4�(���#/!�}�ͬ.�_4"2��f9V�Ie���6ւL��N��$��m]�{Hŀ1,�,�1E<@AA.+ɑ�%)�L�=�^� >�E��3�|�����/�8�;uzP[[���!�> �B]WՎ`,���Q�Oqr(dT��Ą�I'IGq�Q�p����5o�DFE�.�����
�t|V��@��:rr��Nc8A04�I�������FU�D,:�xR|�=4�I�Qj��O���I�~�m���8g`_@�q���U���c'O��MQ�Z���G�4�ô���T�+�Q �����-�x��	���>̜9'�z?���i�)�.�(��J�#Ǖ��mPG���L��k<o��04!��ъ�g�#��3�޾	P����Wcw]�/8 �S����	���'@�۱���x��ב���6�pީ�p@'�2]���1��[�Ͽ��۱�^�j�ܙ�����1����p-6nކ��bd[L�e"��2c��r�D��t|�q3<!�nh���?�"��~�()����3QU^ �Y�4��[:���h���; ���k+-p"�)a���X0w�dS��ߎ]{Z���_8��a�.�5UEp�,=h�&
�InS�j[Qy*'OG@����A����	1��:�N��p�M-(��BA����'_`�ko!%���v✓OĒ������������UKL0�'���d6Zͬ�&sel(��̔0�6�V��@(w/�dΒҡpv@��$ ��+�.$Nxh뤕�H�?&�����x��'�N��*t�0�,\����y��.�C��*�$� �>"ͭ��C�>I�Ɛ�A"=�N9��&p�hǮ]��OXf��Eҹ�8�v���3O�t��~�Y466��r�#�y�R̛7�Y�;����o!J"���'��!e���>M%E���43.Y����Q?�:l	N<z9��֫��5���;�@/%�V�!<��l�K*4U�$� �D����p�r�4ȹexv�zt��R�$fzO?�3�<g�O�%־����}��~	���м���Ғ�eY��:��T1Qenl�t	H6Z]SK�*�р�c�Nސ[[[�������T��#q6'��n �dȴ1kڈ�5%�ܐ~G�h@mM�T�Ȁ���u�N�뷑�N3z�H4���!�
�׫����7nF~Q9&�NAW/[�N�5�ņ-{�q�O��,��~{��2�
�-�ƒ�4s
lY
����[�⫍\�/�� �X��\�͝�d���|�6dTμ|h���@7���|���#�����g^���͈&t����*"rָ�1�*/Bg[���̘>�=�i���_^���#�R��5̺�D��(/B�CC�݁__�+̞:���Yy�`�gX��#6A��w3�I�l�7/+�F�7�K��c�`��E���ކ��vx�/0����W�i��vbA�z�yX:">�t����7/9sfW�o0�G^|�$	�L��P�b؟������vֳz܌I�m3sELI��3�=Õ6��3+n�PPI�:J$N�y���ҁ�m� ��p�(�ֶf1�߸,�6��4�
0g�|�rs�{��O���M.w�h���%Qe��}s�@k��9�+JZI
�u{��?e�8L�8"��nG���Y���PSS̀8�m]���t�1��8U��<�$����#���n�}�s���l+�r�q�ͷb��iH(c�u�=��Ԇ�^D%	��݉�|�I�4k���
F��A^I�0Y����w�|�T����A#"���yL,g�=9�^��ܱH�3�%�����Y��⡨�(���)3P0n*�|�U����M�yΎgM��+���o�����}������ͻO,++�W�R�{Ӄz�拺��rՕ��I�T�X;����6a��)�RP_��@ް�CܢY �n���@B,T����)S�=>�������p"ak�PEL��y����E�9��{��y14��رc���|�]|��{��pe�1�n��9��`>�_oމU/�F,��*�q͕Wb\U֮[�w׮�!��×/ANA6|� y�	������V�Ff/�y�EsG��Xr򱣾u;`K�p�������%��y�}�-��(t�I�ӦLfΎ�F<��()�FgG+��}��<����,9��u#����UU�i�lş��9d�G~A)v�5�kn�S��ލ���Ee�%<OMDܸ�1�t$"�5]m���ȫ��f�{��Ӹ�kβ�8r�����x�X�~������C^�o�݀��^\z���D ���ۧ���ت�`SD���a�w_"	cƤZ�+��%i���	�_0`H�&(/.a\�%/ά\\��1��=l̝	)�K$V$����G���No�y���4'�8��Q�x��)2�!J%��+���������ر����k& 7��L@MADv7�����-��-��x �}]X��M�8|)K ��'W��%X��D���{k��ىq'`���8p�b����z�*��w������𴡲�U���l���O�:�Av����S�o�A�����RF�K��ͅH,�pRG�Bpo2� �b��)8��c��ۯ3]c_�l+�C��������2!U��p�|3��,�
!���xB5Y���c��%G�p��/�m8�`peY[L�����.�g��So�?����?҉�W�l���3+*J�EМ��#)y%�\�p��lNGx�l���&�kw6m�Ġ�x��=���oQVQź�^��ձ���Ԯ#-�\+(��ҥK�Z����|�ъ~Fz��nu�bi�T����\�̳��hd ��ň�w?\��}ؽ��H����X�y�@�9�r|�����nZW^v9��T��w�`�����#=��|,�q�;���#V`ެZHq�L�2�d�����Ɂ��~�wW���o/:v=��x�v��������=}Èx|T3�O�E�1�׉�O;�΁�B�Z��_|���y	�y����;��bu�v|�J~w'N?�h,;t1�9��^�z��0۳������Dv�6�
E���3�ǂ�3سݮ�Y�eWc3\Ոٳ���cSk;�X�H%2��F_ ��Y���)�>��?�GI|��(�/@�����ۄ��n;����S���k�
y0y�X�q�E��0pMCwo<>7�� �]�M�KJ�Y�q��������)���l��؃�@�S0I�dٸ�䵧�F# j�]<�@�lB���i���0Y\�l�H8�(d%pN�B�d0>�h��]�֋/�$����H �?\�#?۷oF8���f�����cڬ�صc6lX�ys梼��q!�xRW��^�v�ٳ�ܳ/`��ǝx2#���PYQ�z�,'"�\�%xs�'�rr���Ub�B�m5k61G�H�҈t����Q��qp"��"�#���g#`݋�a7'�f¿�$���	a$�A$�:)&Xm$2�kj�x�r���[k�A�7��(�O����]�����	��+6��k��?���;���=���)�b.Q��84�E��iVI�4�&��Ƣ����c�8�Nn%���|���6�+'�\�����7�����j�QG5�q�`4<��eo�`9X'��<�[U5F���h��C�n�ߖ��$�n:��V6���� `w�^�x3��'a��s ���x��L[5;Q̟?f���lF\%?���O:��r�x嵗q�AaʤZ�E������i�&���nm����_A����yӑkU�e� Oc�����F����awBTIŤ�cz�1u�x,��J����юu�D�����p����?w�,DC��c��2,_z0�N;��v��-;Y��������� ,6������}X�x6&�����f`��!����1�P�+��W�����l� �peH�$�PR�d�����p B��F,�4��M��8�Ǎ`��U�b:�2�7\y!���h�Ξ�<~QM��O�!� ��������A@P����G�CG� ��jfdDZa��V��<�L;�)b����0��"'?J
��L�	�ffz������^x�1�mlgʗ��P�
a[�@&�\n)A`��!��;������7����ӏQZ�������1t�S�h܋��r������j9�&�����`N�WC�a`����#�������`�T亜���&�(,.F��IH;�����u�f����;:QYR���aS}c.Ԥ���wr�"�̚X��a��8�|<�r�H�?��5t�x����� �p(�T:��C�b�j�������ʉ���g�q�%�p�����'����    IDATꥋX�3���8��8Y?�SI��io���%�w+��E�U"%S�=3B#��(ꖀij#:�7�|���:�Q�]���g���m�ť�SY���Q0Y5Ҽ�9�z�+t��hFJ���f��G��aN�u���l�L.Q�o��/�o�+;��P�E����4�x{�Z��;Eq��aꌩ��d3���g_c:�Q�b�(eK% ��@d��"�S.C�IS��[(,��f��ɱ��ʊ����/>Ì�BL(ρMN�L�<��W�|�j'@2�;z���$&�N`�RIq&N�FV�����X�f��Ք�(w��P�t�҃���b��i���lV�]�W�6g����,
�/��x���τݦ���lq;�ы��2L�� zn)V}��nhd'�ɚ�тu3� t�#�`'�x*��HTDC���l�����B�P�8�f9p�U#5�)B�]����X�+�H8��1>�K7�c�w81�b ���ۃUO��ƆNd�4�!|�B*/>�(f�V����x�H�mL	���zxM���au������j�Vν�J45w 0သ6��<'�5�X�^�@|Ѝ��N��ƕ㷿��U����Q��{��.Ek[#�f���Q�n��m2j�N�˅1c�8�R�� ���{<�xy;~��m6ă~�Lf���I�&c��E3w�|��^�f�D��Ǜ��b������"FB܄��.�:� ������:�Ԓ�0�%)����iD	�c�<���N�c�3=:���D�fx��V+t��H)�|A�f7wЬ��2�˟ro��^?����s�?ze]�ņ�=++J��U�)e���:qk)�2UA���L����g��sN)�����~:Yp����n�]U�G�<�"m��~8��.C^�t���Nԛ=k�y��h�4�y<m� ��1�y�=�u�e<	���nȃ����'uCK;��4�c�T\w�P]S�n��/�����AF� �D(-������_6!N#��0\�hv���d� ��CO�`'tW*�p0�Նq��h��G��9H��L1�4���C\9�啢���p��R�&N@uy)�/;��j
{ �P���S�=�O�o���3д��a?��̞1V����O��.D� [�r����x�QZ1���`Ɓ%�Dԃ��\�Hd°�5VP�nnGWw?YqB�,� W@����˨��@T��NKH����Z5 %3����5I�&��,r�8�&�tB�g �C�k�7\�b�0j���"�R�$���C��M	��?�fG��0�"v4���?����N����+�4TM�"�q��/��1���lF$�E:��а���ٚ4IJ��L(��U�x"��H�[�����mH��y-��J�3m"BHn������R	E�Yl]K�q��N�Ӣb��I�[5������=�ojbHwG�O���*,^���|ww7Ǝǖ�mf`ڱǟ����7m
�d��>��]o�����=�p�-7�3�Bu^n���mގ���v�<��������!��F�5��)�:�Oȱ/�J��I&��g��v�DP4�B�0��P�KC�� �@2>Ī4�� ${�I��D�1T���:���g�yd�>��h���������H>�?���ϯ���C�� Zo�$�A4]2���H`�r�,��w����ی
=?ߨ�cI�d�H�C�4)��^4�����gLfc6O@��2�� �Hz>�j���4�>�\�C#	U ~����QXT�-��N����p(��{�?4�����F:�o~��]� ��,|��<���0e�U*=�Z��lHi&�e����d�b2!)H�������h��_	<H^�0��J2���/Ce�N�>�*E�p����������H$�EOa~�UW��K.�����3V��[��E|��SH�]��O�XBEyqd1�+.>s��=៧R��W�����������ck ��8��Cpƹ'#� �I�g�o�@G{�ن�~}-<�	�ƞ�D	��(F@�;���#�C�j�~+�ح�d�B4�F�0��,��*Tg;���u�àfh�=�C�e�N8��0���Q�e���" ;���Ī��P�1� Cr{䲧f`�Xy���)͆�Ll��!�+ɜ����$"�$�	6�����7Vcᡇc�G�!N�7D"-"%��ʋaS�Ll�"�C��� 3�Ī�d���Iձd�\̞6��EUYv�؆��ۏ�����t���믿Ʊ����2���̻��t �y�]|���h��@o_V��ҩ8�Ϝ
�c���b�q�
�6Y�;y<�m݃;��8f̝����C{c3^{�䗖�l�4fT "����!�Sr��a2�HƢP�2'�
U��8߇�8����D7d>;{�<u�tAc6� iLM*2��MH}Τ��ȵ�+�}ӊ�[������g`_@��'�zz]]�**��j���%�aΑT@&M��i$��%�f�3J��:��{�����|T#��i�����S��2$J��"U�T�S��*���"晏>��(�����?u
T1����3n�7�|���x^O|h���:mD4�UNİ����30�P0=�+�c֜ـ�b��F|��F��K
),�Is]�&��x�?섚��D�c�4t��4��$�>��5�O&�{�o��R����c1o��E����/������z���'��y!x^���jv�AP	Q����f�w��oĚ�?Eߠ�bx�g;lHD���_��c�#�p���"غ�{�����O����������Ɗ����^��㊕6�-��ݒ��	Ӱw8����)[D���!�$mڣ.ii�Y� C�mU�2�tI�Ѷ8 �
K�
� �f����<9��-_r@�� ��뛂&��'N�|�Y�V}QI1�
�����X_oi�/�FW� �4I�3Z��#/ی�-�30e�x=,�BuCN�xjk
P��qfCլx��1K��߃��An��+���ܩ��OQ���D��ݭ@0Dɸ��3
�Ię����*�LQYY�	�������=ظq#�<�tTUU��.%��������{|���V\v�(��BYA�C�̝'�y߀C�L%�H�x�� Y�SU�YS�����@mC����q��7��q�'K����Pn� �+�P\^��'����}h�o��� E�U�8p��)$7:��ל�k���Dd5�aDM@Ei����Yx��GTm����}��㞁}��=����777k�t�ªʊ[eE�I"��t$�r�Y������cNU���1�P0:���tI�m��Z��C�WB4���U����ԩ����l�_�<Y���͉�$�I1�%�N��=��?A3Ya�;�:�H!I�>�^H�2�jӷh��d�Ƀ��x(�a	�`�*zW�,�C�qհڐR���WE�w�d264.�3P��B#R]���U����N�Q�	��"��܍]�M�Tn��V��0�hf`6ɸ��q=A�f���A#���]��W�A"�J�(,��IFp�/��^��͝�h,�w���]}x�//F;��TT�Y�aR2�4��?q/4���H:��y�9��.������˟~��b����Q��B�(D�&C�-A��:��q�&���h4�o��*>S:�*��/=�P/r-@Ei�x|~h�%b���sg|��װ����8y5�e|��<��hk����9=�j�P�m��	���s0}�46�#!M��$f��ja�����<����^u�#��1<B,Hf1���
���0)�'g0��z��~/dE�.�`VE��`��ʋ�wo���%zz�WP�%����<��#�3��7��a�����O?��Ee���#7[��񖛱��=�j'���կ�n�6�S��@iY%�1<��jX�˰��1Q��f�5_\P�!��P� a���?����
�:�\z�)�!�?j���� ��F����|���8�`tC�GV4h�!��Z�$!*�䩒�*��p����������F��Vg`_@�Y]��:���.s(⽰���E��D'��.�e�FuN�QN�u�A��6HR�jlh �({�����N��~���FX����&K�Q;U�E7�X2�H���0#��3}[�q����6��'4�JT&=��؁a7�;�1�� M�6�#�"��	2�VE���4�ب#�H�h�L�5��P�ь� <B�#����AI'�$��C��XNUǂ�S�l��SQ�)��݀�?_�sG7�nSUK����6� L���睍x$�r�$0�̋/cp؃h�h���N>�v��ƍ��'����!��~�)c�=��M�K'��,�GnA�9�H�W���;���]���t�5mC~$-N���Hj9HP�F�.�y���M�#��(�Q��+TQ�,���X�\���K�Bf�3j�0mB%Z�v���D�p�Y�NW�;�E�EXt�b����N㻺v����Q��Կd8�I %6EL�)�{>j*��M�.aM�	Ƥ^Ǥ6�#�Á��2���X��w�d��)��aH&�ߑ������X3�@	�૫���A�$ �i� � Vr V=zh)����в���8㗧�j.��:|�ᇸ���q�eg���o����f͘��NX��/��v�������{w�����du�%Xqԡ��8��~s���y����%�4�
�"��|���J*�9l
�x�^̚R	��eF� ֑�EJ=�X�ao7��0�_�%��g��,������y�6��x��P�|g��Ƃ9�W}��+V�-���n�����}�������!���U7��tj�S�t�;�|yN�Q�	������vF��)��T�l��{5�X�A�u�o������D,�٢ꆒe���*��/����	':m�d���A]=DɊ��a��53y�H
*���(� �	Щ,���&A�[�j�IM�3f�Ɯ?�@8$��e�vtȋt�s:	�h ���&T�R7#�0yhs* C�y�̴%��[ ��� %����]T�F��S�D���#���M�,d�B�#v��d��V�yT�I4�8�)&	�eP��D�LG�A�u{"I��8J*�T�mE���	%8%i$`΁\���)BF`�P6X!�P��$���(�����cн�k�_�c���[�E,a�p�~���Q]]��$�l��+�FS�_mo�]����A %@ � �ӑ��&���E��.�b�%���	���FWE\eʚ
ř��݀��(v��C L��4��BB��Ȟ=I����{@�dxV�0}\5��N#l۹�� gvJ���v�]w`�֭8��Sq�G�r\,�gh%%Ũ��B[[�{�����s���˖b���ݝ0Yl(()Cn~)�ٺO>�"�1C� �7�� �QRL�DG����*du�" c�{�Ϟ@� ��ف�6n�1��L�\�ٳ�¢��Ŏ��ڋK~}��̶l����q�5�9=n��[¦�C�bu"�'P^���Kf޿x昻O����S�k����=�ހ����_}u
���璪��E��BiY�V�a��Ꜿ����T�A�p��y�a��Gܥ9�J�R� CA�Z�j֐ ��
�ޒTY'���n�F8)�#���oZ4P��`���Z��u�-���]شu7�`A���R��b%�Y�H+~��� R�]e�;��-��=%�i|H����.&�a�|�H��@
�YV�y�Կ$���+&3�4�&:���I�4s�	eRf�l9J6*��%���L*�{3Y�D�2�<e���IL4+&��%�jY�I�x�D��4�`,�`ZGZ���]At�;�y�	��L��G0�@������k#b
���,�vͥر�=�17͞�Ζz��Q�U3�	L����w�Y�b'g��΢R��C��؉n�n�RZ�Q���r�8~{�/Q�L"����P*��G�.�2ֈ,��xi��V��·?m����1�aPEVjba���GX��H\�7T�t�N@P%��L���K)$�	���g�N�҉$:{ȓސ+.-.d�&�"���7�"Q�����z
%%%��m��{�����u�C�����pz:^����{B_
4�H��z&
�5��t3�;���6oj���/�/��	��`n��*�Tq@���E���tNӖ�1Exj�]��w�n��y��ޗ�����{�YR�Y�rՍ����<Ar0���`BYT���5�kZd1`$��(9q�{r��t�}s�[U�=oݚ����������y��龱~U�w�p�s�`�(6SE��V��5�~�襳�5���(�~�/�?��yn����[����E]�����g:7'�XHtlx��i���b��p�7��o��C@g)��������(R�ޙ���xۊ	`d�y����3K�ܷ���rȼ�k���}���=����X�m��&�kFcd* �YYR�!�٩*�y�A@��2��Z�Bs+��]���9�~ija[T���n�� ��1 �E �O?؊ �K�Ķg�k�F�!��q�b6t2��Z���	�E?	�L���,�G%=�j��4�@����|)�\�\0� E�f�� ���o���tMJ���ha�Y��O���k�a�.��z}I|��ct�jd��=� ��AV�17l��{��ds��>�}o��ݨ(6�}%|�_������[p�hZ����pL
+�CA�E=�ׅ�_�����'q�i磈����@��`|*'�$��)��cAYQ�T��+Ȯ�
d��3��#�~fG������$�x�ѧqϝw��M�'����x���*"7���E/������LG�KB�~�'9X�1c�+�#a��(�.v�4C�`�		�vH	��?�8�G�b+܄�~�J��4ҭI�/����wf�7ar2���6n��IH�x�Q��ӟ|Z�M�\�'?�?��Vʬ��:����5/?��#�w~��ûF���Ǚ��_������z�	���ĥ�|^Ӕ���W��B7��-�0�	3�0��9�[V�ze�	U��^�Y>璅�p�ƙWl�dE�3⁴f#0
eH�!�S�A�G�\��dd	�7�����z�}��xz�z���Tg;�dS�"<n�~XB�8�qն9a���ξ���e��/�hc�Z�Q��͎S�@�G�D=��I�u��� �U,a)]��;ԡg,��.k6�����!���ĝ��FB,L&Q.d-x�p1��ME�Pmd�uT��Nn�m�_a��S�@A���$*��9��z��Pf衭�R;�X��F>a��Р*U�����ɬ`Qo3������SFԐ�p���z��f�Ꮋ�cp�K��D�E�p�w���X�Z�&Nk^�m�x�L���m��S��çDq~A�"r�>���]	M[���xh�(�K1���FxH�Pȓ�kw�_��W�%_Ca==��]k%�{Z���%��r�$�+
?sP*�sf�lq��965������e�K�jRҘdC��PB9V^?�� w$��4���Q[E��E5h(��?�s�:M2���"v��NF������vx���l<�b�p�Wp��/�I'��T�A2f`��.)��q[��b�XE��}+�½���L��3ϸ�E]�}��ti����W`�_��phh(6�����%�K&M���:˟�qÍ ��Q���.�Q)=�ș-�z{�a#�?a"r`��#@�3�^5o�ܤ~<{���7*|�H�F�{��b��B>���fy���xb3yl�����*�zz��х2Kߺ%�j���D���ln	Gu8�&R�d27��Ntԯ@���V
Rr�M��)��ޔF9�/��޿*�V#QO���B��3n�:F�
�CЎ�X<�e�֝��-5�r�Y �_��n���+>�s�}�X][U>'�c��Ѭא�    IDAT�)�ӔŊ�+֠�9_�K��gk�?s�V�\9��@���&X� ��9��H����+N9g��Dl^�����2MS�4�D~y�mغk���ɢ��0��p}FJ
��ǰ�:��<R�:Lw���L>��w@c�BS������fՎ�h���o]��ރX�b�d�o�%��W�2�-��Lp�y����m@&�+)uVt�
`�h��B��isl^7��X�R�"(�d�4~�*������0bJ���x��ﺠ�1K������2K���k���������'E�y��ж��/^�\�Aak���TN/�U�i�kt��Ň��k~�y���w�7�I��<	�/�{(��)o �Y�sW��B�=�W\v̡��%J���|�g�3��,��z��5k�|d�⅗ѩ2t��+�x�aV���Yb�,
�7��̢����H�W����Ȉ��),x��[�v��:����	f22������*���X�����%-�讝{��=�7�|M�8��g��c��i�0��C���*{��]������q��J,.s�'V*��x���P�%�Z���D� ��	��F744�)˓���_����c��,d�z]@8�J
�[��Uq�c����8 �������LL�y	E�Υ9Y���m*?�\�jl&3�B��2=�}_LM$�fk�������G3Y��P)�� ��r�WC"8Di�uQ�:���u���@�|��^y�	hI �Zp�i�a����<�~�SL7����7��'�\��	?��b��v
��B���C�P�5`{��e��/_�#緢��^��+C�@!R�Jp�:T;��~|7n�{5J~+
U�C���,��m�.FI�46�B�u�<� .�V"� �Y�H�%�|�ܲu2�\?��K��6-�-*B0�����)�F[��O'�����Acˀ�
���N�YV���7�Jv^_���g�0-�z��ԇ��s��5r�b�ƪԏ*�KH��_�����~�&���?���OZ�`�>PQ�c\��-�/��6��^vұ߼�#�>���k_�y��vf ��]߿��ׯ_����Ǘ.Y����eC���D5��[��˥� *˅QO��5�&�i�:�󣞰�����#���i[��#cy�=��1h�h�jabb�\cc#"G�NƱu�6���Kr�=�"�Jb���1�1��/��l��d��ko���� \'=�ߎ����>5K�!��%��y��-ª�Q���@:C:n���p|-\�*@���
y`��ٳ142*U��Vdy;bf���!%t�l)���,���0�C��$�J��t��R�T*E�Ky9?�:gc߾aqJ���B�Ve��M�5׭Ç��G�m���3��>�s{D�#�7���'AO�(a�=t�e�$s|��W�Ѫ(e��Ѕ�ؽ}�ʔH���ﲼ�8�Sx|�f,9�8��:�]�lڲ��Wg)ق�B��b�pkS��%oƋ�4h��0QC%;)��[*�*d��+����C�u�����܄�ݾ����[8�ЖBۡKP�u�:P�.���L:	|J��X ��Լ̚�+���m{Q�G6�'�zԷ��m�	A��B1�6�9Ȑ@�B�;'iN3H�ԥ\�5z���%c�'�s��NP�5�v^�A 7�O~�=����.���cشy3�i���q�Ǡ�)���QB`��)���Kp������P*L����qT�t��'���;��k��(xj��]%�����K�z��o>*5�WoT3O|A���?ǧ�%��*�§-\�1��,Ί�[!U�� od�C=���33G�7����8nI^
Q)}z�\6&2���l�����I̖��za�Ln�����>0��-B[k3V�^-�|�h~����ñ8�e/�s�z�.����[�����%P	4ةPg�b6�5���mELYH�3j�5WJ��]*��$hQ�8���@W̞5���2Όڴ,t���M�(ת2��c��Ӄ��$�������ω;1y]��GGGe��ٺT+*	Xua�@NA]T�s�|mS�e�sL�0��:\�+�Kv��PF�/ہ�yf�f*�{���A�RE<Q�k�~eLѧ�:��"N�q8lq�g��V�8š�Eݥb�"e��H�L���{A�5��\��n�3
��"����0%�b���<N �q��&���/Fo��A��e$0�d��\�[��^�1p��CkGp��[12�"S��W"@W;�_����/W	}� ��J�\g��6�_B�n,:t���uO���ν�B�� ���d�+fڔV('\��<>��.�����`38c�j� f��ݕ[=�V���r}�"��X�r:+&�M �c���PJx����>������+WU|�5S�	����CX<�yR 4���~�����u���K���?�gX�&|�o~�z��"��Q�,ة��Dv7[��[_�{^Ҿ�9�g^�yZ�@��پ�Ν;����O�ϟ�ǱL��E D��ٹ��k����s%�h��'��{O<7��0w�F�� ^J�B"�<d�󙙌���P���)�r`�����Yl\��K�a����`	%6S�&�4�x��bn��I��&�|�#���?��t����-%yJft�p�d��`�еj�WFyr��$Ҷ�d<!�&�	??g��w���Nd&&��� 2��s���Ye����ke)�s=�tf�m�R�����8��й��
Ky��t�jB�PF<ф}�c��=�$z�� g�����:@���Ro,X1�q���jZ�!��5EGLQQ�� �g�x�uP&}\1�Q�e8���Ym�Hx��G��bb�v��9�*��3C�j,�[��d�
���t��!3!$=�L�8J.-�2p�)��ܓp�1KPΌ#�kR9�uB!!��ԋ��c��U�����ZB����1J[��/@A��2�֦�0	ȬPQ�����;'�r�=�h|����~�S�~�Q�no������)9Ǌa�h��cdtk׮��x��)$Rq�YЋ޾^��]��Zx��j�.;����#aǑ�d�8	�/'߁�u!�ɢɼ� ��p�9��e{����ë��˯���+u����إ�`���P�����/��'7��I��/���}E��N(��g�w?�J�����?E�Г6���{^��a�g�;�p?�/�s�v��f/�~fΜ�&q�nk3_�P���#S�0��]�3�h�l:�-��g˧�8����la�o��t0f�Qo>v	2d䖹c(dB1�5�Vc��Y��������i�N<�r��`Ē	��IɈ���_��G3(�>�Oౕk��8��,T�
H$`65�g��,��T���+���W��+呶,1!�K6ըJLt
��Sr�,�3sc��ej��j��1�3uU�`�Œ���X(���2\?COg��D�1SSS��3Hc5���WI*�04:�L��:yRz(�T�yr
��\�aAK����F��n:Н8��U�"�9^71��]� ���:�978U��H$-$��|,T7�%���W����;dF�:�eNDP������H�v#�փ�\	f<��|E��LJ���r�M�
^rT?N;��;b�r�S����8�%�AE�T��8ܾ���7�G6 �b��$*������o9��8�����v�k��Z����f\u���ׁx����p�����_W]q9&GG`>�R	�36lKt�uˆf8�u~���G?���<���}��H��Pq��u7��5�1�-�\�Ag�"F�(�U�����+B%����u3&*�neo��,|�S�}hhO<������JǄ�n*�8�n+�C�;��g<*7.�׃����;�����!�ڰy��/u$6f5���ͯz��^ڽ���|�g�3��,��z��M�ZK��g���{�)i�Ň�.�uOJ�,���*Jn�2�3���lȶ���E���y�Ѭv;#�G�����ęh>��.��(%NF�h� ���2��UO�zww'�n܌?�y�h��p�ƒ;˛�B	�TU�#@tC��qL��ŀ�l�d
hm��3
IB<N:߳Qr7�<�j�����ĩ�n3V��觋���I�̊Aͭ"��tlLN���C*�n��D:!�q\���F<#Y9�<�9�:\�ζvy?����p�َc�2Ll��|�{�*�$�	��6U,j�����&�]gi[��Y{\�ty��;����d97����ft��D[��e� �����^r��n��� &�F�; �҂ή>�i����/Y�Y瞏�\	��X��]�Kl�8 7[�J�M��x��w��,�*��"d/K�䪐���f��H�tQ�WP�tt,8�����]�b��4���Z0��y�r�,0�rlm�f`jJ,H	�.�ȼ
�<l	���g���2�C_�<������A������.F��U9>��F:�U=7�0l��vc����ɵ�cp���7�^%����ٸ����k���	��V	��َ̛3 fPR/נ���Pw��B`Wj8��Sq�g����$�Z�T%ZA��>lUE�?b�/\�#����p}E����Sq��3_�ŋb����aL��H�����H�SH��G?�������:�O����6��7μ��3���:�s��/̝7��T*aF��:�S�i.��W�D����I�P��?@���}t;��[�f�tf���u4��>#�ܸd&�dA��I2�U�~���e��%��[��;���O�¶��蝌�XP�\A��T��+P��)r�ƲI�8s�A�%Pc�v�.��������W�DP��F���.买�JqF��udɜ}�[ l�h�I��F�LvJ@�d?!ґ՞�H����Z���C3屬b�_j�G��|oJJ0�x@*�"*l;wKf�1��<N@g)�ȨŊtÒ�m]�Q�)��]�m8�	���	�v� ry����F���jG�-�޶4>��wc|p+[؇c�<{wor_���i���雇��������B���]�W�5:��L���NlZ��}ð���U�� W^�A��٨L5$�)[C`j�'`j&4�9X���xz���.�%�,v��f��: �mH�h*:�z��̺���$T�� u�ϪN;���m��=%�1;v�7݊�6���?��Ϡ49�ʹ~�ZY,�BC���Y�������1�oۍ7�w^~�1�*���`�=��O~�}c�F`{�g��pk���JE����[k(s��q�����-�A�UX�����7:X�u�����>T���q��4�j�ö(�=���T
1x����B\)?��w���s���B�3��ܜ�����[���\-|qA��w&1�X�[+�����Ҧ�e	�F#k���2R#=�0�&hNg�G#5��C��t6<��t�8�����3��C}��XH0�tM@r��R�&�o؎U��ؓ+��JH��O<�����x��f�Fds%!��C�˶��)�m-H�/D�8�
H��
�zV-���ab� jS��i:�ۺ�Q�������ʄ�
��NDV�M�BN;�s��3x��n��Ma�>���Nh���e�@�����$�q���p�.,ӆi;ҫ�ԫ�AG�������t�I@M$C�'��6x&7lf�&�F���D^2��C�\Q*`�<�M�it�,|�oǚG���K���}5F�����v9�*�i]����]r�-7�x�[�y1J�r�vl�O�G�ھ���h�%�#��q�Q�p����=�}�GP.�}�֑�'��jE���-I$;���_�(���6��T�E�jy������v���EM7�(�B��7#���`=��'���S�ÉG�������p�7aӶ����T|�=�A\,���_�R�V����mܾ�v`��a��-���w�V�1�o�8�Ht�5!�Ӹ��Uxb�V��P,�P��a&h���KN=��](��X�v~��_�F?�t3ߏ�B]	�i���hkK�h��f2Ӭ��P|+y���.hN�8��PN6�v~�ct4�1�loEΫ��	Z1�m���gu��,�q[�_��/����y�?>�ƍ�������=wʀJ	�1�Β���)LB�v(}0��2Fa�Nc�G�q^w�.3�K�e�@@'�`�;> �B;S����Y6%�Gټ�4(N¿������i` �0��#;>)�,K����q≧���?�����|�b��T"AZ�r�]	���h���tPf�nQ���(1��+��7�Eqd?⦅��Y��\Q(��%a�����GF�9�&cE��$ꁋ�����q�R��"Y�H)N��D�A@��v�����
�6P��0m�h���R�+C-pQ�}8-&+պ*��
�RM"$#.���X	ẍ���b]�p�1�Aa�.�>����\#
|K��ۋ��6Ĕ>���ⱻn���x��G�TȡT��]���lKGS2!�h�w�?�e��$�nك�_��ܱ*+H�R�S�:��ubv��k>�q�"l�%#{�R:UMë)�+Ua������mµ��	u-�����r8�Nm�T�b�����ªS�I&	(�z�qG�=e��o:G������ͨ��|��Ex�y�C��������ՒX�N
��a��t����������>�ֶ4���w�S��˔� �}|�Gwg�~��qċz�|�,�G��;�|?T���Z(
D!��EKBE�BW?Sdq�
���3L��85�$A]��ź�2�R�ɧ�#�	�-q5̓�p�sԑ�-�V;�p��G���w�����>��#C�_}���g �o����Kl޼��P�^�?�E��7��r�"#0ҳ��u��L��(S�n���ϋ��ޥ?G��gܦ�s�����y_�����,w�LUЅM�]�bljtvse&��G@߾s'Y�J�*�v�bHo�6b8��Ǣ��7�z/�{ɇ1U(�>�UF2	�X�)��	������x�@�9������#��j�غ�)L�ٍD,�9=�ȑȥ�;N0^C)������"�y2_OyO�gp��O\��'��}r��u>���?I~�:n��&U���*�u4Ec�dk�UŸ�T�_��Ш0ӭ�t-���l��&lk�v������a��01�Ҟݜ�&���x�����ьyq\�ُ��w��FTrSH$c�^ �??�G"�O��%�CY�c�=-��qܿz ���ƍ�ߋ��n�63� D��6oy�Kqʉ/w�r���W��l�q��Q0���̀����V
�_t<z|V<���LӀҔD-m���p�8�B��7��� thN'��B�
pᅯ��?��>\��ߠ�YH�4cI_.<�5b%{�чchp�n	��C"݊M�wa��a�v��b����!D��/��0�w��w�3dJ>F'
���r����ŷeZ�����\����VT'M����ч�����Ӡ�P��MQ��8��z>Y5F����*X
90d6��~zʑ>��6�6��;p�Ky��/9e�s��ͼ��3��������l�2�V+}i��9o3C�W6��妚��w�(�> ����%��q�2t���$�Ay��� �Zᘨ��3*�3��yr�Y���g�/� zK�|��c?q��uشs'��݋Z�
��$��X<�%�ũ���+��.~r�/01Y����ơx6����ŉK�R'������5�ش]�)�2&�� �$�;�O\D��'hҾ3�R'��o�rI$\|��N�����q��pE��1���d�ŐL7	nllL���N,�b� ESP�+2NU5S��_?�?򕒌2Q�����*UU�H�K��ԔB̯a|l�m�c^?��dj

5���3��p�+P
\TϢ1�Yֳ{�Hbv���]�9�ǓX�ȣػgP8��LC�F!MGo�\����6Nz���&������b��~�}ؼ��D�+�"C�cn"��(    IDATo�;r	*����	'�`�[��#@͂p��AV��C�V��=�8��7���t];�ˮ������
r@�<׀S0�j@#�wBKqwt�|�a0�
����k�W�����P̘���t�~�h�)hN��'��DŪ��lcSE|�{��r9@Ϭ>��9|�B{{+6o�w�w=���g�8&3�����9�;�/_��O�e؉��C_��+�澧��N��FN�0'���u��
���X�T}Tr>�g+o��/;Bh4$����Y�g{ň%CY�D���w��������O��?ڔf�_�@���-[V�*W�W.Y��O�a��B�2�8�F�yUT*)��Y:��!&#f+�J���˧��C����#p'/�gޣ5�6ot��@ٝH���� �[�A�-ϑ-?�¦�mx���X���زi�(�9&ǜ,�N
�m�ػoLFr����c�,h\T�Rw'���J�qυ��J�hK�ز�Q��d��rTs$�4�z��+�pG���x��xY� �RA� ^-Wd��n=qJ�Fǻ�����{�e45���2�/��P԰�o������B�D���X�;��B�#�ϳl����ZQُ�[���YX~�+0Q7���,[�Y(�"����w�~��^����A�#�Ö��[_�$I�ȏV�y�v�!�=?�+#β��#T��e�!՚FgwLX�y7���Л:p�]�btx��I�P�����s�:�C;E[���SSԘ�|��wXYR�DI����{q��'�m�X�����ɨ������PD5���7 }BJ� �Yˮabb�{�Yn��~d�5	�8vx�ч�u�>�_��s�)�����5�L����"���oe����{vo�+^y�̙���
^������Q��O��?=@)?�#�}1�9�R��ͷ�;w�jX ��������� N����N�-���%dI��IZ�4Ly��c�|W9�%5�j,�+0)��E�9P��Zeӻ�>��׼��/�mp�c=���g�`���7n|��?,/_�t�;u��.���i�I@D�;��3��8�8��OL���rLT��^V����gg��?�����I�-�����-Iϒ�+f$՚����&��ص�����#�?�lڸ1,у^䴖4�#[��F٩
�@��N��,����CQ���J�c"�0��la|�fd֮��8��KU�?vv�	��s��̣@��uf�!W Tأ��	��:�FF��s쎏�7��\�|>�J-� Q@������뎍�%趶v	��ft���j8���މ����*�%f�%����y>MZ*���v�۴�=;)�t�������R�b̈́W�LdP��=��H����t����1|�Ocq҆M#�
p˟���ͫa����TCW�l\�7b��n)����^jȺ*n��.#�o$�9%.��^���kОұf��(ʢ�759���,���b!KSЖ�I���pUw=��vc����mՅ�?ZW+�xuOG�� t:�.kg+1��jGd�����"�֝w>�ZM[+ng��e�nKA�8t�|,Y�@�>�L��ǟm{1�+�/�<,jxu_�ܾ,]ڋT:����b��[��>���1>��j[�<,�
�E��S��ɡ�_]�
���I-9�(�Q8��)����r��К�4+�Ω�p�z���{8�BY��Y�bI�)�����	��K/:�͟>�?4����ï���@O����<�p�%�A@����w�iCJ@�U�P�X��3tk��t���q��D:�1�E�U	A� ��m)MKvސ���]�7Ρ��/a�O�8q�����R�5Ԗ��c�n�������G�~�:��-�K� !�=s�ڳ�*�S%tU5P���8%CМ@ײ�2c[�ܶ�n���GJ�ct`#�ZF��Rf
~����]b�Zo��A��q%��]�s��d���<L��6K��B�7��UU��	�щ'$��4*���\���	�ʅ�>�:᪎Ύ.L榐-D�D4w��/�v%s�x2�Z������i޺l�q<&*
������±�<ݛ��1�л桽�	��|�˟�|+���8Z;ga�\��ދ���ОnEv|
��uԑ8���C�8��7n�!'�=ق���Fl�4����R��tSCWW7��8��.ep�M7a��0�*�e�H�ۅ81:���N=�(Q�_Ё������b_���Cc����SmoF|a�x>�ۮ��U+�)��9�E{S�.[/��9���T�!?��op�����4Ri_��2���	��5��i��wtA7lX��f�/\%Jpd�������ם.{�7��6�Zz�w�Sa�3���"��� ����|�\r�RPod��q ��	[�q	�:'�͑�c1��@�"���b�K�L=-�<�P����~�}�����@�����,W`П�=_'�+J���]�u����%w:S��# �|�Y���c\avzta)���o P��|0����!Cp����'����פOOh>���|,3��;vb�]X�a�n�,�KP�=wN9��]�_��w�Њ'Q*�(�b�A9T� �[�nCk?����T���8@[Y�@/�ds��G-�GGk� :�@T-����3q~^���'��?+�/��
��$߅��y||��Zx�F���9̤����������۷W�L���Su�eϗ����4G@��ˮ� ��U⪚�@��C�7�6�9��WU�*:RfÔ�ܳ0Xe�(\�����H��0�S�G���4�A��u$���Kdl�a:J��Ȥr��#���7adbÅ���qر'�?�w�؉�dQ�\F��U��'��~�綡���xO<�*�<-בnn�W�P@G{3]؏8�KUa'���k��M;�b��$�Q��Z��Z� >&����O t���hoI�����U������O������(�3X�t��avw;&F���[~����سg/�<�x�^�z` ���_�|�Q��QQ�ҕ_�1G�Z����q���ú�{0<�)b�\_>���qEH��e��_|�)=L[h��89 ��`l�WA���Ш��4�	ɖ�GN�hY�'�S+��8�ێX��e�n����^t�R�=����+�����V�Iq^P����	�졇�3M6�ܧz�����(YD�ǥ�"@����~�`��W�$��<�3uE�Q��}D����2]` %kP1)a��@I@$�?�r��̙�5?U��[�lً0w�\��W��KWc�S��]N\ƨXr��C�Վ�E���p��Ӄۥk�:�,�rPsET&'��5�t����PeN3��A#�b㸶ak!�H��H �cd�!4�̦GU)!y0$	R�����[�^XVg���⍕ 9g���d:%Jy�:5��J�^��B�""!j2������j��ѡ:qԌ$`6!@�l	�r����Hi�B`-=�?l)�K�5�����%��Ǧ�P���GRw�o�n����s�jy$�	�:��sd���{��o�ޝ��U_�~�nz��旑L��ũ0h�1I*���H�pd���2��/�s�6$cIt���箸Cc��KvL�J��>�~2.B9v��8=ӘC�Ba����.w&>��w���D:Մ��f\yŗĴe��|����Х�P.��k�Ʀ�0�oGy4������`��}��G��}S�)\��O�}_�b���l	��A���o�d�_��ʮ'<���Њ����)Q̒�����[��{䬂�8M�)����zyt�kL��k�o��V��Zx	�+�,(Tv�5l�"�s��/��5�8w�2��ڷf^���)��}������j�����\2�m1_b�dv�֤�UC�U��?(F�_���e��F��z�oȠ2+��v>�D�(c���	H2��l5��bC��kQy:�jjc�#��Z��܅'W�C���9�$Ri��/F���>��˰h\��2�Í���e�rZ�˗�X(����e(��y躏x����0���<S����vT�.�<�i�#u�yl<�x\o��  E�~��Ƿ���gBSWS��ey��(s/V��j.��n�|';�]��b�*�}T���4�)�1��3��MH��iA]K@��0j���Dv�h�t�.�Xfo��2��Y��Y���^�.�G[#Pyp�
x��D"�f+	[�1�
���,A]�F
U���
y�lY���r*������iK��t��mm��Ąn�P,�#|�KSQ+�$��*��_߈��.lؼCJ�f,����9���!��V���U2�2�Ⱥ��ܨ �ם�]�.�пt��?��^G�W�O}�9�Lxn��ǰk��P��r𥫾������8~y�o�_�
�XK/�׿z����5k�~�6�z�������4T]�k�8�xP���-9B2$σ��6�^��&<��2K��	�tVcd�*M�CF;��>�'��@g�#:�ԫ�iK��%�R�m����z�;�~Lb� ���m�dj��U��<f��.��߿)Y�j�E�Ͳ,%t�RG�N���E`&�iȘF}���~g�}G���3"��oɶ��q�(ۧ�tt'�y� (�r�t7����z�� wm�!Jc�Z� ���#3>!�}�qN{��%x�o��?�~��_�\%PC��i���4(]�h�?EW����HS���J;w �k7�BIf{�:�Q,��>7�N��+�m5|���Xz'�G�2׍���7���y�S����i��܆�F�kܩ�Da�|�p�������#`����Z ?��j�
�P�N7Ao���g"��S-��(4J�:7|y}������]�Xg+M:����bygR�&����1h+/6RF\l\��*%�51�	+��Z;�e�0��*��nl^�ȗa�iMn�[�e�hi��\�9Шj�Q�.���M���5�4$�\Q��m')}�L�(��μ�0{;�KA=���S��Oed�d��x��$��LX���O=I�n��C����Z.�#_�c�=�#��b�
��ae��+8��c��7����KՀ0�N:�8�͛���Ùq�ɾ�g}�NmuGm�EF�z�#aídm=��1�&�M\�ByaEe��!�qEM�z~�-�f�E&P�~��ue�^�IS�\��s�?w�qP�<��i����>�>pb���~G�y�?�
� ��,�^�zV���pἋǑ����N�-{�i���R�"`!l���@�Q:��e�t^����/�����	.�R	`��d��h2���&��!�Bu	&�w�6���y��	�}�U+�wݏ�n��c��/2����雋�#����dKp������\Ϭ��/D9�QcFB�0gVP��Ԟ�ЊTG'P/U7m�u���'~�(���x|Q)��+o��.
��B��/nQ���e-�k�[�va ��Z�t�b0��?7qʖ�
j���0�"��Hr�L�ҭHǒڿ2�^؏��K�{��l�G�t�f�(l�$Ņ�--�iM���HϞ��ZCow����-Q��<��X��hI�a6�2S��zu�+5ĩ�� Suj�İg� �w���H�O?E���Ŕ���r����Dϝ��g$G0Ά*�a&��a���R�*�B��S	�,�G�d�B-�]�]�`��}�I�e�
Bf����}�j� (��4t!'�2�D���P�O�;C���:5����#��Ф�^��T�qK�l=��M��zP%EQ�z��@��v���� 䋨�L��⢢Fy>�D �EĘ��a�2�G#!~\Vx��`���4�1�62��^]������/_px�4s��_�@��B�Z�t�d�O�	Iq���N@���F�=b�G����FO}zv��G�$
a�>ҵp��3����� tE�e��|l�_�a(��c랰�Yrg�Α����p�m�����-�_.WK��R$��k�6���\�*��T��\:���0�{ѱ���
lLMT�f��Q݃�����!zT�*��z�f��פ�I�K�Eo�ą�p]�iY��~�h%4*�cC��r����	��P�&p�K�k���P��䊊�OrWX�T8S�>Ɔ�ZM[��q��uT~Ճ��Ba`��
�;��`�s�o.b�g�j�j�Z���Ş=U]��������4�t#[*�i¶�VC}�vī<�Xں�?�|�J�dB2o��VJĚ:E�޴Hҫ�!�L�v�֪����hغ� ��AE9�A����nT�fjЊ%dW��T.����ZЫP�J(�B5-%�g�����.ϵ :�7$$���+�D �A�Zh�#_J���@15���|��R����j̈́����|@�ZY�C��^1 ��u97��y~�_�v���Ke@�A5l!��	�b��p*�,�Sѐ�F��k�K���+U�"��t�	�t7��u/}�?_|���68S���eП�=O����[/\�x�|*������;o
�sS`ɝ��7V3�5Rrc��=lx�����(*�G�&,u3��#mv�A�x�S�B03u�9����x?A��*�L]�2�c�<��j���X�z���j�:�.?,@_�a+v�X�	�K	�R�F�tn���о�PT|U ��o>z�������H�:X�J���g���UA	]j�G��-ľp-B-�Pio��~�;2Rf����Z�nu�E�ň�e��<
�E���Iʬ�'k�x���K�ꮨ}���A�}�۴ ���_�ff��UU�=�}�X���c8�DZ3tk�<$��@�W�U��������B���hM5��6��6n@��$}�+H:,\��w	 Z
0��S�d&�ꪁ���^u5$��9��x�hn�P(N _,�7�;�`�ݤ��\��9pT	�Dn*���t'6�@�Z��Ѳl1*S݇Z�#�f���u��ɄEu?���f1\X0�D8���� ��X�fB��_�w��Tq��{����9g�}
��P-]8����b)�_�aIQ��q4R�P��]c����4r��iF߼�hnm��9��T�TOAfr�6a���X;�J�ݶD 	�ň��Ԡ�������I��m�^�v�+�|�u{��i[�y��xf �9^���9���5���C�����R-�)���\�F$=�z�)E�M�ǆz�Y"��yuF�b#
�D3ԑO��pI��N@�Ζ�KQ��b��M�r65��FF05�bYa���x��uص{/���I�Z���x�K��ۇ���g��[Q��Ѕ��̃=C�{g�u�bT}�c��	�n��q4�.ܱ!TFG01�W �rbhikC��]5��3�<&��jU�.�zLՙE�u1�o�=>�棬?�z�-���LE$Y����W�W��_��(��I�Z���Ԃm;��-gѺd��N06I/�40>�<K�SY!/ʈ���c?����g�y�"L���	�<��C�����×χ�D�0Q|����ō7�P�a���8��Wc��^���o��-[T+�ܺ��QF��#��?�65�c&.xÛp�ވ�9����-#�xp�F��ڟ`͆��_�|��es�2B!�tؼ%���sX�q+��f$.F� ��u��LVx�� ���Y^�Ba�*�%��V
$)a�C�\����fuy�(����ཆժ"m��3S�:�`�);��O��q��1�sz��Yk2��7p�8t�B����p�1�#����
�S-@*���������_݈U[��N6˵A58�#؎�\,C8JF�t�Й����[���5���>w�c�>5��
� ��|�4�O�����۶m[��}?�N���^��Px� � ��ESd����x��%gY�����~jB�jd/�0km�9���,�ҝa��Y�0�%�U���ˡ���.'��ً{|T6�ΪB<��^��yq�q������/\yJO�Nb�	�4�cXj    IDAT0��-�r]�G�-��$�*:::L㻶ah`;�PK��������V�`Ⱦ�;4$��Ϟ9%0��!�S#Ef�������E@OP%x���Й=����C"���G�[e�G�`���45É�e�\3|�{����B]G�Ȩ�21�� z&�Q!a��n���f#9o>
�ӲQ�?�#����w�}�JYJ�a*:��,��W⁇�g������p�O���-�������J�T�0� ��^���q�׾,�b�wm�n�Ӌ��6lٹ������sp���P�طc;�Z-����a,S���~/�dKhZz�@���n� �ᆮ ��hN��	�d���D�͑^�T^��c?�$4�u�&��<?�F�.Brn��΢��e�T-��-�L _,�T�bb2�J�Z���P�oF� �QE0� �:<NFx.�����} �4�_�99}&/p��?�W|�'�4�'qVt��z$�v�w'��{�QA& -[9*Z�y��G��g�z�/�mp�c=���g�`��ß~��v�
�����.�q4]��_��S��n��H��j��9��ɢ,��.����+,�D�͡e+{���J]8|?������Bh�b���v����:����p��'P�y�uw��P,�{�����5���o#_$�M�W�������g��u^?
5��p5,?׋���4���CC�pL��Mp��~6�$�VB:E_��;`s:].wzu#o)�6z�ӫQ�>�Zy���/t�����K���t���z M�P���$ҨS�2D�VulL�LAӒ0\V>�̶��W�x~ck�ni���Aӂ���>Ws��cq�ůF9������C��)ق��p�8i>vN��?�9>��"a��_��(n����}���9:f�Tm)O���XB����\���Q�x���Ǔ+�^��Ö�EG)z�?���𲗟�e���~�;o�E���9��Ga�\vŷp�� ����ѪP�y����{��PG���D@g��]s.�͈������rC#_!�ND�.�#Ĵ����F�z��Pc��3�s�c�wJ�V+.���X�J�N��H#_vQ YЉ��	��"��J@%�4pq�.�G?��tZco]A�X�����&A�؅���E@�~8�&�~$0K'���N0m8F}��3���>}��f_��y�m���@����9}���@;P�����]�3��:K����3�I��|˟�U6"�,<�"-9W�޽Ј%�O����s�K��A�����$EA�ĩFW����c��m�w�ѕk�Ԫ�޿O��S��dD]�8��G�{Ɗ'V
)�Չ�</TiIS��tQX������i8�t�8Բ0������B�����U�$ǦSC�{C�� �E$������dzi=��U�E�̞{��O�h�"��аg��u���NR!�G����.Y�F�������L$PwR����8���&�o
S0X]�aЇ,w�=�K�b�jכ�^u�qx�E������_Ǯݔ�M�H�p��_���}x�񪗝��O>��u�k?�Yt�M�¾ͻ�ljŇ��9&JSC�������럅��q��O�=��h��Dݫ �N������&��Y	�|%܉	��:>��Kp��B�\|����MH-9E�V�MӢm�0
Ő��W`�5���w���.�h�r�P)�Ñ�P�!��}�S'�g&��?��N��^Ι�3}�dk�%�M$!�&�zG�5�&�WE�(�H.�"Wl�(`A@����g��N�3��<�3����ߋ�p����'$�;3����|�Sx�>�g�Lr�����K~���0���"`���;��s/��Uk�!<�A�3?couAW����Q��'�/�$���������_}�UU���^�cש���bb.�p�W��o�?e��"cu-\Q1v�ϑY�%D�<+?�b!w�y_8�?8w�δ�O�j����N@����=Ғ%KBa��֖ƅ��@�'e*)�#RU �<��QoΝp�����^y�=������-�Si���0�+'��׏^G��:v��I�#��	��Ƥ�~~dpH�=�J���Ͻ��_|�l��2���P�x0⁈�g�.PդC�ƈ��҄��t�S$+�MI�I((!h��F`�ѳ�h~���;�g�J��x�}��r~$jP�]�;c��?+7a=�G���7���*g_y}*�G�[�V��B�+#;n�;wڴ�u�o:йץ�n���M�h� h1��<[�`G��ud�z�r���G�3�8����D��:�Q8��㔣�c���з5�n�C��iJc� w%��L��/�c�8ϼ�&~��P�c�$�P���wM�ј���^�9����O=!ϝdȁm�0<�DˤIX޽	�R.�i�r�hN=�p\r��duo����ݻ�����j�d��C�[�).���l�G�Hj[u�^ꦫ�vy����
�A�zn�\o���[7�����a�nl�Z�X�l��ׂ΀��h��r�aBǰ���1s�,/�7�GC�X���W����/Z�,�|��.	����g�e��� ���}غ�*�>���<�4<g�L�S&��c�_^~IVW�-��
&¡�x����
:�9N�|Тq$��w|��n;s��Otq��͟���}�P��^X�fM�m�7��l�DbPE:��Nq&�;ԗ(�q7�G�\r	J�N?�+�X�41�2+��;;soo^�i%��̈�t����m���(E�2
U���Hj�dR.�5U	�Y��}����K/�{�!(UM�VuUB"ʖ\>2%��.	b�~!JcjƍA�����6�����Y�"�(!�}3�B�DL�e��oz��T�tNdn{�h^5�S�G�2�e��"��s��������ol_f�3����k�k�g&�ߋ:zeP�����KQe�Ym+BF�F`VI������y������|A�d��G��� ��#��
��\_��ǌC�Q��Q؂S�8��qF�����à�b�
��1O��\PSइ�ӿ�㏞�{�=^���#����4�P�i�M��<����؎l)�}͝��kx����r�j���+��#xu��9��-8��p�)'�*�"p;��ݻ����E��ڸW&Â��CՋ��<ύ�-��T��a�a�����	Ԯ-�w垯������[L���ۚ|���� �r��];3ƽ�T�I�?��b8`={6:�[��D}#��؏;��N%��\���`8>h|�y��\}�Q�R�B:�?��ظ��p����s:v�<�B �?���t�����w��]��|Fȉa}�HTpCCJ��{w	����E"|��p�'N���_�,��3����|N� �4r7��{	�ýq���T����Nv�7'�ѥWF�}9a��`*�d��]	@� 	m���E�&�:�fyN4�B��^)(hk)�Gݮ����W�\Vtȴ��Xo��|s	��^�?��W��u�8f<��} ���0\0�,��g�Æ�k���c�r�i��с��1��uJс�!&�,�d���2�[��2�4����Z����'���Maj���Х�ӥ�q��y�����8湲�,'`��GT��ބ��!C_��jy?Y��</?�F*,�gꟹ"��C@���v���h�xv��j9�FvC��YNxϏSU�_}c��;R�\nA��K��N��'r#y��ݻ�dc?|mH�sRD�������p�<\x��x�W��sω{��MX>�#P�8�4�����]�Y�m�C���ڶ����o�x
���8��s���
�^��ٝ��o_��cc�����GD�h�͈Nj��������" ��̎@-��\E�1��|~��3�	����ZٶرQ,y6Ȣ0�9q��?��W�])9��暆�o=Q!Y��fMԷt�m���]'���ow��;?zY���t�+�;X|t}�s8z��ʙG�
6b*$�7oьFV}4D �)������[q�!��&!VQT����{/�͢�)��7�|�m¨ښ�.:�s�=e����eo���?<����x��֏��r׏��%M���S���Y�(*ռ���
`T@���
E�aS|��>~��J�K�}p��9�ycF�{I�^��zń�/���u�����=�e ��!��B�Qg���6n���-��ӏ�m S�cLs;�j���)��M�Pt�z��x����+�H�~h�m���B�~c�� 8�<|�<T� M5R�z��S��& �]?uޔ�G�ܕ��K;W��O��=u	l���ө��J`��%��=��Zy-��5�=�G_gq��T�5��̥c���BH,����LX��X����J�J�uT ݊�����2tq��͛�T =<i,"�-H���+;E3g\z�03%|���,8(9;i
�O��\/?�<J�$�?�8��9��_�O��Y������+��"#�����hj��O=������[�򶋉c;��d��܂�)���SO�?���=�ęG��#=܇��v^}��A�����d���b�@� �f��}z�kb"���D��zPu&����� t�^��?,�d��|�b��� u�n��u+��t��*�>�8r޾�nh����p�]!�FiN+�DB�t(�s4�8z�\~Ƒ�@,� ������T>On���x �cgo��q,]�	_��70qRF��V�Y��ZNd�����5��?]�G�-b�N>�����sj,�i]]��ߝ��9}mW�Z5ʱ�7�w�	�{֪��d׫��A-	
HUV*����w����,Wa��[��z�� �GC�8�;CZ8�����av�d�{�/iͅFǰ���7��%��� /��lnnF4����/;F]uQ�P�������ԆH4��,�Ԯ��6<��$��ϙ�R��`[;FM�Bұa�խ��!�
E�Va���b��F>=�M��erc�RG�9O�+�LfR�`a�vyQ�s�d�<�`a#&;;`���Y{;Δ�B�M����T�)F�V�>1�����1������bb9~�.IMqJ ����������%đ�סg���T��+�	�
�jE��EHF�AG������S�#7\��Ͽ����.��8��c�ۮ�`�o�۷���q±�b�ٻ��7�g�=+�`ds?J��TyO%�:�|�B\v�iΕ���/b���j�1{��P_[��)v߻�.4���1G�κ1	�<�,�.]�@4���,����`�N���ЭB�^D��ag���FWǠ)6\K��-E%k�=��*��d����W�zA'^&�Wh�=A�5�<�J�7���/#\Z��sv�I���A��
k�t�x�C�*�?T����,hV���t�`�
�.�/
G�V|Uٚ�B4��o��~�c�;�`��~���`p�DÛ d2yԍjB.c������ۡ|o_xډ�~W}N/�;��'<����	��v���t���$��=��az�ڡHP:+�>ޝKZ9�S ��YNB\�bE�*%P��;��.j�
��`�J���2r��y@�lP{v�z�ch()�LYㅍ�~>�J�zOO����Vm�F]C=��0�Zs���H,�W�[�HU~���������4���+�ۆ�ɓ��t�@~�f �JEiUb!X��F$$����V��i��H�T!����,t&�{Œ7���rB]e��u�e��ǘ��忳��:vW����Xw�@`�'�:��
4��%��۲a�I&?��0Tf(���r���J���_ �zz=G��:t��P;о��2���˺���^~)�F��/�z�0�ZG!���kK��;��c�������F�����~���W�\wE�g����H��Sq�-���I���+q����x�//ᥗ��o�-�1DB��4c ��ĥN��O:��S�M� C���3��8�[�$FA:� WA�.�v�R<Q����=� -�+���ܼ��G־�����E/δ=5 #\��lA,�O9�Xw�~�Vբ;U�u�?�44X�X�XX���'���I����g���y	�}�Oxw�:���<�'5�4r1d� ���{X�i+ꚚP[U�O�iN��[��� ����SB�����hy��f^t���}V׵�����N@�t�������76���m-��g��حr�J@'���*ma]�h(��v�o��*)+v��3��g�Bt��<W����*�������P~O�&;ږ�aKg�G�,rEx�x��We�Hn~/�3������.,[�
o-y_��ӿx�H��� �7����[��7c��Ux��O�^��l�p��F��e*�V	�b	�����u@.d��d���e�(���O)�L)�Ŋ�A�#�m�D�?!X^)�_2���W�z�'�퍵y���q/$B9�������
����%�[|�٥����B�k(X��rC�j��0JZ��Ѓ"�"�;�okѝ��CO{֯��.�����!4�	z �.�K:v7g��E4�QF�#?�{{���yt.�p!�j!oY�f���/��zꈎ��I��DΒCa����S;��/Ǆ]���`�HfG��ko��?�B��v�W1~�X�<� Cj\���b�O�q�57�7�Gb�d��Rg:�t�hf	N��h�	�%Ϸ��[9oR6Bߗ���e^^)}\�Qy=��WVR�����S��3�k>�t��a8�K{�qG��C�C���E\{�}��;p��W�y�����C���G��E����F:n���`��5(6.��\̝��<n�U��/����j�%[|�0Gn\Ѣ��_>7�i#?��U�/�Ǿ��|���f���v�����?���;|'���/ȧ�s�/o2�����V���
�WHi*w���G�� ���m�6<��3B�aW|�'���]���U�;��3&py@]N�*~�Cb9b4o�H������m�ߥ�Ђ��M�3��-ߑ�
�F������N �s⌀~�KV���m[$�b���b(A46�!c�(���-۱i���,�D4����:m*F�ܥ���
�,�|JM9�\C>�b�J6:M�<���z�4�I9���5O
r��{��~Cg7��w\�?f�Sf�	��u!�n�Ƚl�[ٽ��g�#
|�|$��%�ŔE�'�`��1�}�t��E���O�?�	���ݗ�"�=��Rf���s��ъ�	�X�$-q�+�`�3U]%Q��u��*R�A�I,GQr4!�G�톐��~�R9���k0�`!�1����2�ahQZ<��:�� Ǵ�iSW�$سl5P0�\� �M0���~���h�,�`�d�U�j��
��X��|,���e��#�hJD�u�f�r1��C�z�����V-�L
`�Iq����ie}��'X��X��	:�_�P�f�9���/w4���7�U	l�q�=a[J��1UFj,�}�bGǩ���0��BdS:~�����W���ѭ�2q��&�6�QO��t�cx��%�\w�N��.,��)�MJ�B�r�{�P̏�O;�'��9��S���S������v�gtП�a���Ʒ;�ƝÑ�D<��^��)]�Hh^�'�kMSo��Ú5kp�W����W�z뭘s���\de�hzv�-{�6�s�t���f�����†�"��Ѡ��v���<H���ׯ�����A�����r1�z��װf��ߺC�$���kj��9�n��A����\�ᴗY΀wTJ[3:�M��&�%���%@A�3��G|����/�@7�	V��ւ��j��q980�d2%���I�0�}Y ������3-t�bpxHΊ�]w�^����qcD���(���5'�<��"���^8���:4�� 
��p���+�ҕ�"�'�P�i0�afr������ZT���)o��� �ֹ�ǏG����x    IDATC�pTX��pA�0����[|�m8V�lC�!�A-���C�SPCt�wquo��m!&�q��x�l9������:�E"�׎���ݶ��[��l�錰�L�q=���g��?ؖ@R[����},Jָb�$��G���I"��A���)�,�D�J}������>�!��ܽ����%~�O� r�""�tEC
�(�Sp�i'ᘃ�'�5}Y|���-�C�T�zA"Q���p걇�ܓ�F� �L��z�&TWע��5� ��`W�����>��>'�aS����\�xӞ�����He	�1�㼳O~�Y�n8qZd�'�>���8�O������?�}���'_�5kִ��uk�1g�Cg�,��G"p���?�&:(c�\� ��쬗-[��=�(:;;q��s%���t�p�˟3���:;�X<���|�e��
���pUW�\t��"\M��-���7���6���� �ѻiy���M��փ�۷c�g+�2]�DL�>��#x�c ��qr>��5����$�;`��&4O��#f\�t���i0�C/!gVu�&|��xuw��Tǫ�X*F�џ�=�c�
��J�F�`UP&���������*$���j���'�'��.�A�*'�7��~�"|�<	�๼��R�u�]H�҈��PfpӫۛZ�й𢅸�sQ,��v��۷�C2S��EQp5��*�$>���M�?�f"܍�<��X)���=��6��N��p{;�'L��M�\��F�ڤX�&�P�P̧Dz�.kE��y@sJ�+,ń�:���W���:�iؼO�$>� h�|�l�D�!�O����ek���ȸړ��՞ �Qd�I N�F7#1y2\���䉅\)�a@ѳ��;��h�[/�P5p�Ap��{�X�����K���
\~+�O~v(��i����������2%�?儣q�s���º�����1T��l�F(��� %�z'�?_��0�h�K7u[V5�q}d�.�b
�����O�//^����6=)��Q{��]�1����M�%[엫�jq�Q?~��{]u�.
��w��/8����9}�-Y�j�[;�ƜQt�]bGY��{�2�΢�v��Te6n܈�˗��3P�Κ �ۨ�zjއ\�h��3aLAmm�3���:��^{��*���L(��tvM.�x�ؚ�z�d���oDMM=�R(�ͳy."�B�P¦�A,_������8����1#�,�{�ato���;�b*��^n_ZG�a���]fJ�_I�2�}��]]��}JBa�7�E@Sq�]w B@�� ���D-���p�73e����sr����<�#�6e����O��w������W��gDkHη�*�{~x?�`pe6m�e�}��C0�:ݐs���^ge۸��W� �M##W�qʙ�bE����1d���u�h�2uO�1'��MF�
C)�l��v�z��,��H؇� 2v��uaء�%V�T�ՈU4=�:�WL�0�X��gW���0TK�_�a*%�|"V	��C���"��;�e4�ya(,C��8�K ����lA˅��0���kr0,�kP��V���i� EB#�{LN�Y�y�J%��,b���*��:T1��8	|VA��>;�pQ2x䷊��-�3\+��Z21"������۰}a�UH�)`SpΩ'��� QU���n�-w?����Q�P������[*b��Sq�i'��9W7�p%#T1H��?ۿ�e<��ȸa(�*�& E�_�m�h���Y*���LA�g����6�N8����l��^w>�Ox;��g��}�؎�7��!����\���N��L�e��v�Z����LQg&##v>��9�@�vy�N�Xv�$��jk�p��˞�ie���σ�-��m�E�'�"{[���w܉��~TU�
��`��?G�e���d+ׯ��� �Ϙ��/�N�&3w�� �nي@ ��H�P��c��������M���m"�p�L��W{�^ʓ	��N;g�~"�H�����/\�1�m��s���gqՕWyt4k�M/��hno���;v�4I·x�}���y&��I��)'2�w�h,��>�0��5C�b�;�?���=�o��Ȇ�2Fӝ@4,c�o�'w���q*]2m�|��X�q��1�7�jQ�5����~�2,j�C~8�%�B�!��ad�z(�T�$A*�Y����B&�y�ݰ=k�	�`���#Ǝ�r-�[R��	�*��*��u�)��F��>8(�.�Y�Id��Iw�����݇���as%��!�`�L!���g�p���'5���!4,���O�D�Iv���:���K�v-t�C'�]c��ݲ�B���M8I�t��1�@���?M�@����g*�Z-�LJ���N<�0M��tS?���/1PtX�˝��,XXTs��s�h����8l#�P�/���pH��J�`պM(*��Q��3�G_ޯ.�3,Z�SV�0�:r�#�4ޏ�Ɔ��s�>��o/��3m��ʏ������O�e��w��T�un?a���w��٪ ��(��
r�"6oތ^xA�I�sv��*��lO�l�_9G�̷����de>��ϗ������n�d�
S��.�m�'}�b�I���_?!����G�	?O g8��ۇ����k&�w>"�*X����{�f�VhZf���P�a��*�|�����M =���g��!�������7}{M��B%+�ݫ1��A���*b�*�\�w��#$��RtT�Ǆi�<q�������׋�xB�Sw�w/-^�H�U@
�� s��rˍh��l>+�v���{�y�}��	pi3KR�h"���ӦN;J��#X�t��|c^zo	�h-� ��d�+���U ��U|��6z/�C�HW��
hk�<p����P���p�/�U�Q�k���`� U�NҞM��&�|��	غpT��F�,ax�J���fۥA	g-J�OQCСT:w��U���� �n"dY(�y�@���`���{͂���v��4���r�`��n��HW�"���N�8�|�S�PV�I�9>�ne���*��P/�ߙ�N�%����U��`-
\5X�{&�{h�86���߿�����I�+���A߁P@�^H�ʦ��J�S�X���(~QH�נы�r�D�P� L]׹p8�B)'�3�9-z� c$��[�:X^s�A3.y���_��/p;�S9��� �S9�O�N�.]ZS,��ۮS��qW\&�0tCƳ�8�U}�����9�{��IgQU3J�i�7��X2dWˢ@t���9Mkk+F�TI��w����Qκ�/]Ӡ�R�J��d9����t�ry�X<�H$������I��ǿ��L�DO��n߆}��g�{�5�� v۝w`��m�ð3:�C#��)0N8���n���#~�t�=�W �)�hZ�q��W�#���X߽
k׭DcM��x^U5uض�/��7�]��d�T��}\���K.�HR���H�
��;<�U��㕿���P
~�c��˾�*���/�nr4ME�����a钕X������YFbQ�YD�a\v���}ש�¦-)��ށT�t �:����-�~Gp�yMR5�t���)"��R�ȓ���Գ8��p�W�@���ry��//�ݵ�%k��Ia���1o�t�Y�{�}dJ
��(B�RI+P�D5�Hz�T.b���5���A�r�-��&�OĠ�
��q�t>��1�1��C�đN���g����!�`H)X��$���j��'��Q���'#w��m��{(��1�HF�6b>��p�Lٚ7"�(T���T �c�;��Cy*�?z�T̅d$��5ٙ����/9*�`-��w��u���7�Z۰�'���z'����Ģ�� S>o���B��,e�E�@-���~���ۆ�M$R��H6'!t�Ӡ� �tz8�#i�E'�j�U'��?�t��~
����]�Oi��uG���ug�/��%K�D3��{�1��P(��ݳQ����
���rLh��#w����SO�E���NF���;d5ϟ���Ɲ/o�DLF�Չ��\�`	v輀�k����Hr2��uy'^�s��;��z�����J��fy456�_����F��ؼu;�8,@��
#%��y6� H��t�@~���Ku<@ooCݤ	��";F�dl+m�Q��Y3q�g"
`[�F<��0m�Ihmn�d-��-[�uݛ�N��y����S��1��9��5Չ8����~h�(�vv�o/����ǯ��>��Ǣ!��~:&N'��:d��;������[LQ�6���	���)��c�Y�a�:�!T$s�6k?t�>/��?x�a��h�9�%�2M&>ڸ��C��-]dsj̯�q�Ep�է�?��5���#g�T7�>n?К��_���_{C%E�e�=`��"�d��6�*�,���}~�h�-D"�9��iiD�Vg���[=�CׄI�L�~Y���=>�c#����� � J��L����5�f��eR�ס[���z�g#���YϢ�����)5h�[q�����M:��@��>aU���,X�$�j�7\�W.<�q�l�Q�����ދR������s@�Z�����3p斳p�Yu}���c� ��l�0�>��/?�W��$6�(�s0�T~�H�"t�rԁ�x�����w��	|�5�N@����֭[L&��<e҄�#�H��8���~	��e�J�.[�?��;��k a$��虺�
y�;/j�:;ϱcǢ�*.���G1~�xt!���3�aG�ݹ��!_,�Cb�і�HP��_�!�Jg2���TW��g���-�F�����Ĵ=v�"\]��:�o�y6��#L�=E7�`&PD8r�����2O��팁��sAY�󪪃�H�x5�1�oGCum��EC�z�{K�ek���P2-)��\l3;:�P�gQU�ԉ0��U�
����1wޡ�ƽ�> �d���mW��r]�b��I��.��v}7���ho�T:���\�I<�9{/��4ҩa��c8f	���ee��"�s߹�}�C�z� ���`�p� h �N���˽�߇���;��������Q\w�7p��GacO?����X�7D��z
Sۛ��/-@u"�d���b�� Lr#�gJ:�$���n�J���U��$��,r@/e�X_�G� ڛj�I�˿�4U~wM��,PMD�(!��'nn>���ؓĿ]
y�������uv"KS ѡ���r�و(��8tO/�� �;bpˀ^٩Wd�ܝK[�н.�����C�Xָ<�'U�Ɂ���3O��{�Dm=������ �Q���jK�@�ѡQo�d`_ �� @+e��qf`���O��B����Ej�E��"�LK�����c��9���W�2��F��\�a��y��y���.��1.���g���Y��N@����\���\����֦k�x-�f��@�u�^�̋N0D�k�.��C_�~��8z�>�!+t�"!��hʲ�k^ m�XԎ��NEډ�h�59���V�a��h<F1��׹�}��u*|�|>?���x��Ţ\{z���ko╷�b{� F2)465�.D��N�Y7��l���Na�<�/�x�-M; =����Ns�l�x�;@��@u"�ֶf�oCm$�Iǡ���D����|�]���CQ�08�*�"�homBo��84w?L�4	�ea��������؂��`��M�WX���>x�]�)L�63f�!���ۋ�λ��"Gk���_�0�c\�o� E1q����4��䠼��Hc&�yǝ�u})|�;��Fyc[5 �2����]��c4��B^R���7�q��������I��ٿ!�2#�B�Bp
)�s�ua���!T��7n����ۯ	S���P����IeL�c�� n)�]���Xf�;����k�_�5�dl� �1sJE~.ӹG'/��E��F#�j1�5q�� �w��F��jCk�G�)R�	��(y�n��
"[K�� :G��f	�\3�8�l���2rw˻�:�W��ޏ�RF���I7<������1R("	�s���P�ԆU�S��?Ā�?Z��}��H�\�*�K�T,���N�E7?��P]��F¨�	��p|6�b4���b�J����|��N��O��ǟ�Vm�E� ��|��}�|�҃��$צ����=�����}m��>g����m'I��l���BJE:5��ՙ�D�HUE._�mUW�Z����6��uu�Ì�{�P�!��>����0gh	S�*֯�y�^&w�ӺR@��E�#�Ury�����=SvR�UW���Kj̩o���/�/}Mm-�k�L�X����!�ɢ��w���
E`��(E���}!����h�<^�₪���>��S���gᣅQHeQ?�	�MuX�n9�:x���;����z���}��7O��~4��CYX��xMZ[�}�:L�j�٧�
S/bt}36lڄ~E��h1d�:2�<��ڰǞ���W^¤	8��C�b_7�����7O����H�J�"52�Q��؅U��bbW.��"�&�|F���勠&�{�IX�-��~�s��*���5�e��xZ?��P�M���$`먯O�'�܏�S�`���{��5��e�����N	��*�z�eh߈�x��(��̮6ԍ�ƒu[�upH��󪐊)m��.B���x󵗥`�{����~���>l�U�@Z*��KH0W�����ڄ�}}�h��ql���+�Ū5[�+�,W)������8��XT2��t��50��:B.MU ;t10���q%�����y���w�qsY���5?Sޟ�$�u"�l�^���I�ayr<��"��X,��睍]&L@}C+����7n�%L���β�L�)�C�o"��O������|A���J��1�
Y�#AW@Q���a�a�����\��Vc�޳pС���᎟�k�� 9������7oϳo=����Χ�	N`'���������_�{ܸ�;C!���>FIG:3"�T-B8g�ʭP(�Q;�-��a��R���L��ӧ����9��(��=�X^�������z�ǚ��ݡGt��A�;����d?�y�"�E��b�m?��s�`�r��{6�Ϛ��V"��m�$$�.������4��
�B�G��J
@m���]H��� "�W
�W�~��-j�j0���=p����s���/b�	�e�׿u����c���&bL?=����S�@�WQ����7ߌ-=}��T�tu���.S�j����	���ga�Ţ0�u�=q�=�c�
v�~Q$:Z:��8��Vc�Asq㷮����O&��ނ�W,B�f�����ޟ�%�qo�8����-�]GR�b�&�H��1JШ��rx�{q��=�����3�c�p��a��U�4��q�6�q�IG!��O�7o�Vt��.Ù��SO��߾��?�,ŏD,�#����8 Q+@M����⦛n ;�?{�A���7��@����pM!MC}M������f�i]~��`�3����G[�4�Y�q�%)��!r���Q���\[F�I�R�'G���'��}+����|EV[���g��~0yM	F�kfx,9#��������1V��6nO���~��A��>e�Q�D�WBM����j��T�`�aT-J�ako��b9�K�6�ɗ�\&/��E��!�A�@?��!�{���>H����籮7��d
����̂���٭;��>����x;�S:������o����%��vn}]}Su5�۶��ى�����nCb!�E�3�]�^�y�1}!H��6c̘v�8Ø�8�//l�0U.\��s�}r��뼽�'i�	��v.� ��	��{P�,��
Ӷe�������ʵk1o���l    IDAT!�e�ݰz�ZK6&N������Ç�mp!v=��A�em���#Z[�@�z �71X��HZR�΋��9 hf3��+q�i����G;w�>_r9�9����[��S��hoE��6���_�`��ƿ]���zWȁ]&��|�C#X��<�%��8��s�^�s��w��]l�^'�=v����,Z��B	�}![���AgWҙ!ԏ��K.A]u2CItv��;��*�֩����M��g���(���\�H��^{A��m�1�h���.�TM�p�58��#0�zsy,�^#fD� oj�Ĕ��h����xe�V��_ ��(�RXp�A����rc�>���ٌ���3N<�A``}?�bh���*�x�'p�?BsS+��.�,�t��J���I���\�H�	;�xu����a"�㚋+��o���L��}*�U�O���c���:�jM� �*!@¨c!F�H)���
�q+�9틂C��^��3���c�{�z�C/þ���r���@%���e1i�x\��|4ԎB,Z�-�\��{�sB�݀��(�!�^Q��!���҈�b#��c ?�T;�37�JA���bņe�C��3Jz_�xm�S#��<f��w�=9����d\!t���__x����091���^����	�����ӠN��v}�4�2'\���N$b!ƨ޸�K`�$J/p/)�,�)��SVVIc�K�G�x�u�yt�b�i�y4t�_,˔<�:�]��~���%��yq���enL,K��x���`�n�=�`L�:�W�����i�Г,��߃�TZ �����ҡ��
���цz桗ea�����D���*ng�fǢ�4�#C[q��98����ӿM��[�nǃ��P�t��)��D,���eK���I���ͤ$��,��g���aŚ�ް��Hx�Q�������W]y�ح�-�у?A�P
鬎M�{aM4�����3�e�z�q&��D("X���w�>u2����+�����G�	�����!b$����
�[C)d6o�o�� ��0��	w�u;��1Y�@�Bik@<p�ns�>�,Z�	Ï���谁���2ƍ���%���?��;�6����=3�W^v����u�	hhh��7\�Џ7_yA|櫪�<��Ev$-���MEw��k��ƖV8>?z�J����xE7F�(�Y�h~D�j`UoXl��QsnJ(OU$��h�J�C�s�Z9���ty���z�ȭL��b�����@����_&W^����A�2e��ҥh�o@Uu6n¥W]��吜l���׬���:��$${6 �s�X[����WT����%�f�E� ]�|�ߪ���߫j��U#��ah�&O¾sŪ��}�C[��������|�ٳv��������?h�o�=��>��7�q]�H�6��ibJ�s�D�q%@�hw���k����d�Y&�xyʟ�m�g�S	;�\eO腴T���^񵮤��B�2�;H!�3%�39�J����,o�Q��YQCl}�x��gнa�:�xtN�e+W�v����^�����aK_R�|qh'Z2���c�C�Y��h����k�iy�ZdO�edJ+�ݦMF�����=_BS� ��G����ò���Ao_F�[��3vA�8U1p҉G"ư��T&�W�|�Hݛ{�d�j�܉��4F6���-8�ģ1��N.�C�����H�HgM����-��L�>�t�a�8 �:Z�㙪*R�4��Z��7�o�u�E5�"5�d��@@�B�7rwRY$9r'cߥ/��H��x=��o_��}f ��d�$@�ᑒ�^y�,۰Y�� b���ƕ�����7FFl<�����م���x���0��W_u7"ؾ5���](:�{x;�j+������Ln|~oʤ�~��;���kW����#;��3��k�b�V���:�`�y�{�~;nq�����&Ac]*c�9v/w�.\T��^1��X*�;X����UV�T�m�����Zt������Dm2k�t\v�Ũ��A}}6l���@j��4@c5@��Ƶ7�9�ѻa���+b�L����Y��s�``���FO	�����a���7#Az�M8휅xw�v����>b��osg�xb�)�/>mF�K�y�;;���K��3ҡ(��e|�0��dW�� IM��29�h����rf�L:�p6�]�*�i�Z:�'�p����h�Y���d	��l�p�X�{��ȝXB[W>'�\8,	-�^������M[���V�ڀs/X�1�;�l�j�&�:[t���b�P����X�C�elj�>���ױ�j���]�������0i�X��6U����x���ol�䩻b�ƭx�EX�z#�l�8�GF�%0uRƍk�f��mCXcƌ(�L����xg�r�\�%ΐMS���Fa��8`֞Ȍ`����s�!p�X�g��Wto�G(�@&9��1�hi�¾�����f>�u+�`�	�m�t4�'^��Wlƍ?x7���_S�5����g���V4���<�i/�2P\�UB��s�<�DD:|�BFw�əH�0�J�9+�0���|^X�-� .<�z�����Nc��lݼ7]w#�9�h�x�1RP��~�W��Mݛ����1֬y��>|�I�S� |�T$2.�x��x�/`�%�b�=�Ē�[�ބM=I�2:J���{��x2�+�7C�|�� 򡥹>׆az���41�)O�*�^qd�W\NZ��>+�
R��s���}"��t��*�n|Ё8��sj�o�Mۇp��+��1=$f?`N�b`�i�q�~3�n�2UȧS�E�ҝs��)�<d��. O[d� FF�B��
���#aOZ���셗bٖa��o˰�?�ށaL7�ӎ>�kN��s~���\�U^���n;�����+��{n��ud�m��*Nr]�Q4乌�"Ilܟp٥ˀ�g&$m=+S����%���M����==����
�WHq_�6�#�&=���l��gR�wj�U�{9'!�� ��v�2%�D:��{�����eشn3,� uM�x�נ"���LlK�������!t#�� �p�m�b�I@�.#�Af��|e@��+��#�;�PЇ��vߵW\t6f�>o��F2i}�AHf���v^x�l�2�b�@ Hs��n���8�kW�����O�&롟>�G���$��;��ބ�z�;�������_<�,tt6㏯,µ7}}}Ydst��:F�p��o�Q���o��'�&M��;��&��L���j�~�/�s�pI�b�L�ߘ�S}(ad�P���C��P_���|���mh@��C�](Z�`����M�,�pH�^U����n�p�E砳>��d�Y8����>~ؑ����ȥ,���t�eX�t5��G�q�R��Ø0q�������щ��) FR�ؼy���oL�uV�ۆn���<F2:1Qr�槽jYR���,���m�T�����(���^�ޫR�x�sN-��U����@+�䊪��+��b�t`Y�x�:S�t�$���Ԯ[���=_�P�C--mX����%$3ԭ��`�Y�X8��q�~���_�B>�����F���ԍ7Gu� �9����F����>���d�@ �BIG4�	o���NFF���o��赑��ӎ?쌻����z��{>�'��?ǯ���`���3t�<���W�����e)/Na� ��I�
�� �b&U�`y��Q�Ʊ=;z�[FA��e'){po�ͯsGN��\o���M��n���Բ{�
�ĝ���@���΅Eq��Œ����`�K8�S��ȣ?C]c;���CK��f�����P�y����U@E��C0t�S�6���,y�@��=�P�j�;E��nx�;AuT��mx���q��ǣ�����c<����;F0��uJ�:��?�0ƶ��|�z<��S8��31��O=�*n��(9~lܼ]�1�������#�������g�¼����'��E�q��o�Ȉ��ޔd�+v	�0p��/�����p�6��������mmCҲ����Pt[�{��%�N`őu�
�t�V��tγ����[n@uMW~�k��6"�4�b.MN��wX,1��C��ތ�| �?
�f1�F����A�vÂc�ctM��f"5�E��Z�"'�x��?������5���]�-^$a*�J�ߠ�Q*��eR�O��~sDc���܇[o���"�S�f��H,(��QR����N�$Ѡ�-���'�Ӌ�W@��a��+ ^�#�2��2�'�{S,�O�8���dJͯI>�>����_���U�ol��8��/�XT�r��0>�R�?h{����S��_���-�+v�G�Q�	$$!�L�1�`m0�1�`L2�`��&� D!!��P�3��s�P��9Ճ}�{o��g�/W��XB�鮮���w���A?%��`yY%�_�����C:���E�9���
0u�T|�z�}9tKD"�bg@j��]�޲1xsM�I�0�`��ԟ��S�l�7^���|� �{B c����Q�/5u}A*���\.;�d���ٌ.�\.Q�D�DU��Z�ɵ�r�Z�����M3Kj�+��t*��1d�I�vƂɇ5JŲ��]d�������2�\��#�Zq+��'�K��!3�Y�څ�Gq����tu��$��ƌg]�H�^Ą��1i�\X��{�Y�^��g�z�f��rw4�&	�U	���UW"*Z�*�5����`8
�$�1m^�e��v�D̝5O?||*�����/���Ǐ�;����|w%����œ�Q2�Z2�?|/
���+�����ł��p��b�{+p�]���gw�wKܲ���<<��#S|�Ǟx���,\�]����?�F,��f������W_�Lb��%���f4�����c�b͖z������e�Pf8��9Yh�TFv�f2���f�CDy^^|�9����_GG,��i"E�᪗��(p������
/�xϣذ��;C��].m<�� ԕ��	G���4��^����G���.��6q�e�� $�v�*���`�}���acC#w<f̘�-�6�������܅*(G�P7�z��zy�A�p��m��o��)t�6�Sݴ(f�6
:<n	U�E�B����R8�8$�Q"��H��	_q�"�<ݑw�8�����}�'b�Z�D�ƔE�/�cb�Z�1��W]u%��<�WU���g�u!�Q��� �,,=��'$�y�U������X�6s�l�И"�N:Y-8q�^�$1[W��W�Ɩ�����E~n�� ��s >��ɀ�;0�$4�z�������������������wx2��o�Dº.�����x*dYIʊ�9�?�����kf���M�������d�Q�Af/W��dCҖ���>%�.}�IC�+�Pz\�T�s�A�rn�������v�Q�4�#@���'��u��SEM�>2��8P�6�(Z��nv����Fa �C.FsC>]���p�/~��,@*W�_l��y�Y��v��f���]2<5���t���>��t�C�5 -~�<��mL�P�g�A����ի�SOCU�X<����`��G�J��v5-������ןB&��Ƶk��gkP;f,f-\�7>��=�"4C`+W��D�A<|,��W_��O>�C��1<�0�Ep���!��zJ����8��۟�ٺ�}]]]�?"Y���>���6t�% ���t_��kI�t�;�6�h�`�(��z����+QR�!�3�6�~�x�i����bY��??��w�#i)P�����V��0F��a���l�J�xME��vmن���k�NȖ���<.7����;��aŊ����F�h�"��������	cY?m�*�;�����؈P���Tr�KC՜�����:��9��TLg�.�0�LNJIDNt�Cv(���{�}�$�Θi�?�#rБ�����u��:�w�H����x�*��N�ה#.���8＋aj
:Y�
�	#ǒ��p�QG`Ŋ�8��v贱*.-�~�T:�d'�d2���ޛ���
$c�(2�:�������G�f�/���1��a���B�������u?r��>�۟����oz	c�X��p����(�_׍��g�T�X,�c��dY��j�'ibf[[�E��5�E�.-]OR!�[AiQI�[��a��	������YGZ�F�%O@.�g �P���X��[����PÑ8k�=� /��p�m:)ZRV��AR]lKJ�Ma(���c��;��J��CGAi%DO}��^��;��a�{{Alǡ�21UxkG�_S�I�H�``'��c�u2�q!��ts:��`Ԩ2,}�1��7�g�BgG�:�<�A���X�z-�c���*�S�����OA����V,}�U�]� u3�a�����+�J��B	8��#�Sq���G�Z8Ҷ������hj�ēϼ M���mH�Uh�a�t�X�h6v�܆<O�����U�σAUf�3�f��b��r��ìC��{ǅL"
�K�$ou��햫�Lip�s��-(�W���@�e���;9�w����:KpqK��4���DKC1��S1�F����o�C��&���@A� m�����CA^J��H&z
��*2f̘�/�~ʠt̏��*s�ҥ<�kU9���6�?��m��y���,��������Q�[�j3P��:DJ�Z�N�NO�}�E�
=����$�FN�8�ܸ�CX���T�}�ф���-�ɝ �ؚ��'J���QZU���|lڼ��k��I|�\�g�X��,u�X��^&����ĉ���%0L�GX4*#@'��A�,R���苈�4���#�c(2�ʲBӦ.\����amS�{bhii#Y\��/<�/�ſ�2�����g`/��O؞zzWW�wp0uC߉�,떅��n��'����7TVV���+W��<�����t�'_l��Õ_O��*)ztn�R��[�U�ؚj�]�]۷����<?<n/��	�G�jn����hh܍��ͼp�.77/((B{g�|�m����M@+*y�a��
"KU��c�Wk��IVQUR��/AYa!,�@~~��� Ô��㾿`�����R�}�&$�
���S_u9�0��U��0�-��ڰ����2��D���?���(�{�q��E8����tv��e<�iǳܶ���������S�o߁m[�#��Q���՟b�&�R,
�%X��<�=k*Z����ކ�`�g��[�|�O?��[��X�sٝ��8��;	��|-�ÃВ(27���O=�7?��ǍH4�ȞL�����s[�y,gr�dFs���_z鴍��nl�����9{:o icBY�.Y�����7��0���@FP�q��c��)�U�L���6-�<r�_�U�q��]]���^��^�[�P���yHD;`YփϜ5�DJ�S��y�x��9�����ƌECS'V��J��2'��ܝ����`광�Ц�*V���|n�� �K"eН6�� wAf�S����r�����g�ǜtK����h���#�NݫlBǾs�b��٘4}*,(.���[p���# [A��Q�$Lb��98�G��5�!� M5I�,�>s�񸊾e��6(͐���,�c�BfQ�4t������r^���h�5cQ7s!>�Տ����Z0c���u؉�U�{O�k{���={��=��O����:�����`0�����m����7�_����荵7?��;�R�H�Z�L=���<�v���=�����o�,�}޾};::�PUY٥����Og6�e����O?e'*��&�r@zx}du{�)��tK`�|>L�9'�z*���L�����(�bTVTc�TL��Ua�ix�
WT=��ʃ�=��mN���0��2dA&.7@-�1���Ξ    IDAT.G�2��D��0��	ltn�/��L���=г1\��q��c�g�2��F	�Q����Ȓ!��N�t���
����3�ܶ%6y���������	ݠ0)� �4R�<m<.��ltu�����Itc��x�et��2&XN<�`g����g�$L[���J��o�_��f�J$`K*l�<б���(�|���O�Hp�k:�����ȣEyE1n��t�E0{�<���S�7<���}�Вqp�!(=���������.��fҴ�#]�w"��F�!�@�����$�eK�G|��r&O���/��� >\�6��zp�i'aG������;��������~�9�汄���n�P�f�.�xSwHR'odx�@w��?z22���BJ��E$�#�M�8J�>R������J����{���e�M��;:	:����Fr(���>��_�i��5UX�����+ ^غ�i}4���A��1?:_��>/]�o~=�̝�ҩ,��* ���!�\H�B,u�z����{��=2��#��1�P;}>>�ԁ����V,�?{��'v�^���2�o��{���r���u�Vu��Ɇ������ͮ.�򗿸��g�]�19k
�)2R0�H(ȓp��?��� ��+�Fia/��w�<�Z��v/)/�:�	�<���!�xf��N��$R▅Ǟzd$�$������zt&N�
o0 ^��L:Zyb�G�EV�ҙl��yӘ�e�M��@�����i�rtʓT�__�S)� �����ݰlx}A$��#&�h�<c-���GUM5����Ջ�Ͻ��p�[��%�M�83A�Y�UUW��ο �&�=�̓H�S�d{�ɏ�T6,��C�Gie9�*������	Q�`�{�#6�K �TL�]���=��#� 	n$dҚC|K�)���B�盞�3��Oz=H�(A.��`؍���'L_��/�;Zq�	'��3O¶�.�x��,1���8����+�#Ͽ���������LDcs?^~�]�ڰ�P~��#�p�{ �n;X��G��w7ap �`���5��h޵;v1��<2��������S��g���̮񕷡.���F6�;��k#���܆�����J3��K"N�;��� �}���[��X
��$<�ҿ�vw���$�q��"%ÛȘi�eO<Շ�@�u�i�P>xB����ӝ�B��г6[�R�\Г8��y��ч��O�ë����MS����GAVx�N��h#:�M#���녙�`h8��}===m�x��ND��EX����"hmi���Y'p�13Ñ�ep���_�����y I@����ݟF���k_]�ȓ�n�m����U^�DUq �^wz[��T�����$�����IM9�[�pG�q����ww��H�aIQ��D 58�_zє�D4���@u_R�ӥ4)�ʞ�̔'G~�+�5�g��L�������d}���5�Ї!i&D[��֯.�'����1[㶪+�B�Hq��PEFլ)PKГ@���%��E��KG77��D���p�Nڌ�5�K
1u�L�̲��_�v�
U�d�#T}.��O��QXY�F�0�I�+z�wv�"E��i��DM����L$:ff/�ɯ��:��>�~lq�[��I�ug�N6f�	OѨ�gL�=���,���V�w���"��)[f6;�x�iӧ#��X����0�6vïJ���s1��kw��{�K�A0uL�)�տ�%nR��ｉ���m�((�@4�Dmj��	���q�)?�sK�rYt1Q�ե�q(q/�ǽw ���A
B'K<tI��M��!��h����N��[�	q"���Q^Z�B��y����%��)w���sI��3�@υ��t&�cL�>�Q�6��Co�
*�1��N��`�2sZ7����7A�}�)`VR����1�`������٪�QmX�Ɯ���Br�a(��F�0�����=d@�ɢ8�0�M&�v�:,_��C�H6K�&M���QӰj{/6��Bwo\���3O[t�	S�)�g��{p����"�Gx��������=��+���O���F�����!O1p��'!O�"�ӁHO���2Esqh����U ��U8��,Y���q���п�1zLW����{�� RY��lS���
��
N�b�8e�g�����4�pDsS�8L�*.��t&���tbu'Ӑh��b.�Nfؾ���N�2�[�k\�����\�;���&ٖa�I�Nr:��t5y<\!/4�o�a��$0��
d-H����2ҙ8��
C� �TL�g�)GV�V_3��eb�
w6���T���+�!y<��m��KQ�Xh�1��b���#5m�g��ٌ�	�#K�d5��Qb�;[$��e&H9�a��릹k��e�!��PUU��
I����I($n@� ��'����R�^�	E�A�|�9������q�Ï�TOU$z$�x���^���W|��.��mIɠ��DDAA����!�b��YH�c�f�г��q�ɨѣ1j�x��o�ڈ��aj�#KA���e�y�<��;6���(�	�̠�4^��i8�6JJ�pZ��S��c�4�1wdk�S�?��|�	D�*mP���22��sn�wx���9�� -Y��.���E�
�,Z�
�L��O�O�9��|.�i|���J0m�L�3���:�@�x��#6���\JQ�m���klش�Y�T5�u�=1�R"Vm��ζA���P[Y���g��_X��=Y������=��B�.x��n�4U`�iC�'�H?����_!��=2���nv�D0e�T�ر��***x!&*"വ�a���<'lh�ņ6^����He4�KJq�7Av����˒;�
����3I���WR��Տ�p��"W/ن<G���aZя���Of�]��N�v)���e@�IJ� �2�lodc9�J&�\�%�I�P�����`�]H�N6lHu�"���m}�#E�+9:QY&>r����+ʇ�u!:Eo{'0� �:���Q����!KQ��U\��qc�+
�q�}���-We:ivD�#����P"�1��U
�������D`�Tpr�U��%� �2b~[��悮W&�6nqЏ_�sj+
xo����
UɎ�]L�B�PD\�x)V�9���oQU��M���^B̒�Y6�T���SN��� �>��&/�q�Kq����[o�*hزu��ZQ��Ԇ�eX�]QV���nŌ;�&M��Ys��у;�y ����H6���d���-
6��5u+�M'����m�71�D�dB��r���.&�f��1���sְ�1�MK0S)v!�s���X6V��B�>(
��&Tٞ� �gL�
2w�44����'� )$�gq���p̏�`���ã�,^�`_?�T��Ä��1�{�y��Q�ģ��$���l�������2
�G�b������`�N��g�ї@�������>��c'�O����c/�On����=O.�p�3Ͻ���E۰��xB��T����k/�P�V�����D]*�/��?�[�o���/^��g��$Xqq1>[�	ƌ��¦�ɦ�$cՋ�n��@m]0-�&C(+C?��I.&�Qۏ�=�W%�R�u'2�M�i,ɀ�k(�h�nv�t�񋧥��P�ȵ�) �%#0n4�U���d��B�g1��	NA��*ɔh3�nb't�^�)c!��#j�
���tG�M<���b��j�R\,���!7���C�z1�݋t� ��a���)��xp%M�YU�R\WAja>b����>�%�t����kSG�������"�LG�D��T�sW]�SC牶Aܙ�זefw{dnP��~�ſAmY�����C��Q\��/A��0f��U�y���W���O���k1mb�a�==H�*�li�,�G���Q�u�¶d�����[o���/<������ފpE�0,�@6�DA��7*��}ؼyR�,�Μñ�D������K�`4	�$S#s�躒o��N'�Q�E�}�Uqt�$�ͮ`;m}� �}.�7f�3���]h䆖uf�-N#�Z�;#�QgB�-۲,�N��e��L��[-3��ݳ4�'�g7�^��9q�:�_0'�x$�y�Eh���{I��/%�(��@aq�4Qr���b���s���ƣ �ť�=�ePY7S�-F^|�����h鉣0l<���p�q��O������п'�o{�6�������[�}����4�D�妑��G�e�^�u�5��h۹	A��D�	'b˖-<C������/�̙3QYY�����$���u_�B6�n�b	�Μ��;p�7s����V�xC��)�*�1�Q�NaDHr*k5��N3ur8jC2�,��QD�Ԗ�! ��6Q�x��m\2�&�����x%jB�`}30���mK�@���\z��v!+	L��T^
N��E���$[: ����4�s�/�����-��%��B�#\]�F;��(bݽк�� � �&Zpf�T1�\��_U��&	HN��������<��~���Y�_F�'4���
��9]cnP`�4����llʎhԖWi�L����!�uaժU�V�<rW�V�������b���(��u��c��~��K�;�fC����E2���Pq����nG�c����W�Fiȍe/>���-hjm��C�Y�PO?l�@�����v�j@K[;����&`��\��[�=�P4�6["��iCH�<=���1�"9����N!���F����L6�#!F�Tmӿ��@���~�b'���	�9�"k-2S��3)�`���z�����q�	$
��O���;�=����i�p��G��O>��� ���l*�J�E6i����=>
^�P
�1�w�cx0�L��'td�I���~��}Q7}6�R�tCZ��h�O�� Tͥ���ť�{`���{��������`�2�S�˃_����]q�a�
�ZF�({Qr�Kσ���CY8���n��b�m���pIa���:��;�]7���Wq��<��UԌBB.��uH�&v5� �&A��D�U�T�r%G�� ����ÂC��m�""/v�y�67-���� ���(~�X�4bvIO�c@�hL	J<�!�H"��:���J򆀍m��P8u<^7�-�B:���A����Y�qN�_��'Y"�Q;ݦ��,������r�J��Re�#��V�ӹq����1�d #��b�_8w8Y�)�#�6�l�oí��X\��l�����ad��ӎ�PS��p�,w鋠8��9�l��ܦU���I3��m�)��΋@a'Yn��u�ъ �x�A H�%��1�,L;.[�©~:2�\� ����Lȴa��w�z�C���]]���>�x>[�1�&Nf�����5�G;$������!jƎŖ�����ߡ�{Éw�� hҶ��{�ǝvfNt,m�h'Z:����1����'�e#�-[w�]H$�=z4Ǝ�#��;w���񮢈��j�R57������#t�h�5o�}x��m[z��_8��A6�4H�t݉C@/�De�m��ZO�,2����c�{�&}H�#܁�Gc��'�	�=�~/T��^�����P2�d2�K�ʝ<��{��pQf/\1/=�ZW���$z"B����~q���9jo���vO��K@�'��{�d�҇��_X~�n�]�r7�BE~n�U�q��CI�@6M�[54�FwO~��!�������k���/ěo��`2��ωD"X��BDR4���w�(n�$@W|(�8	(+E�6:�7��;Cs�m9��ʀnC�,�$jC[�3�O0��C@���j.b Nz�*�`�dx+JѲ%�h
���@,�d���T��b�E&8�~��;q�߃�A����]КہI�)�Sd'2�R�r�U�|i�����^ǎB��vFC�Ɲ�z��N; v5������v���KX��$|��X�q+�|F�I��^��9�lgNk�n���,�W���E�t�N��T�i��0Gk>��`#� �x"P]鰸i�,�n���ǰ4�e0y��3�ҧ�.�L=�l!�L �֑�g y�45���"<��m�^�%D�<���P�F�tT'��0~��x�ɜ�i{'.��*4u�!�6�[2l�qȣ����W��9�L6�QDZz����K.�����ogE�H��瞃c�=[�l½���$PF�ۃ�.�fϞ�5k��]wߍx<�����\s�U\9?����,��t��y�D
���v�? ]�I�4,+yJy1�� �_0G��|�|t�5��!f��,;&f2p�g��%�[�C�hsG#'�2��xhdQ5z�?�0�%��I�������>�������s�Q��|�����w[�������{n�'g�܇�?��g�8�+^��Ase��A�L��_y�֣y��P-�'LD,���_��~��ƣ�1�F���xfN:t��'L�֥&�A�gʰ�ygz�yx�Bش��(�1Bi)�	"d���ij��i�Coc�1��Z��,B�`h��X�Z���y��d3�ѫꊊ�	�WV F�ϴ�GS��j ����T���@���?�@՜鐋�C�%��[@��ٖ60��[�"DS`V=���鴲)�xl^��U������nkF���mgִBd5.�3�ɜ�f�4Cw�9��̱�x��f�?�ͭ�ܥ8�30<4�W^|.g�F���� D���@�!n\������9!5Nv=���L*������9����,X'�tRG(����8?�H�;�����a1Q̉��fL���tݥW$��Ͽ����M��D��MvhVMZ�}����)�Y��i['.��J4��"�Q�_�m83h�=H�M:�U�юhQWĀde�k1x=&N?�\v�o��p�57��g��kDc�믿����^���7��/?��{��Ѹ����q�UW�F�2���on��M(..�+�.ý�?�Ξ!>>���N�t�����f���w��t�i�����֯���h���s�("3��C��Ix\�ob�)1�<�iDA-x�l��|f3ve��lRK���'��s-��������GL��R������3�9��������K��B��o��\���?}��ղ��ܴ�*p�6�:�
7\v.��f4lZٰ��J����$a#cZj�����seN�l����{�SM<U�u�b��v���ӐT6m��z���J1��x��T�>� �Vatg�r6tɰ�"�l�dt�V�J��\�\D��Tn���������r&���j"�^�H�gP5O�f�?i"ι�B���}4E�u����XQ���XO"ͭD��1�E�8�_7M�Y�4"y��6�Omc*����nd:�������aR��Z�Y�Bd9�#`�eʎd�7�T�#~�4��$i��A�S���8�x�=�M2��̀Ǎ�qu��c8���ʝ|�)�D�$����Ѩ�K,�4j<�mR�)��<�̥.�J�����͸klã(<cd��M�@�Z��o<./�t!E�(���.=sF�1�6����G1��A���(-.Dyi�M�{�o�։�}�Z{�6hCBD:f��Pٹ�㸸�K��hA�"(*p��.�R���Ͻ��.��s�+��p�=w��������^���kH���B�rۭ�W�W_{>^����W^���>���;Zq�n��u[OPl0��gjD71����D���3�AסzU(��	�G��3Oƪ�cx���V���k-8��!���Y&+8X��eK\
^"����c�`�?B��~GV�߆�(�R�͌���|����[����wy��wy������'V��>x4���Iu��6��0}|~��_�PM�q�:�#Qf��"�t�����#`�ū��ƪU�yVHZض�Nz��܃�%�e?n��O�,;w7C��Q:q��0�&9m�d�~��;=��N�A-S��A��W$H}C�n�
��0x5�    IDATM'Ŋ��V.�]&���7S�Q<a"B$���/���t�j��@���Nd9F&�Ys�œ�>������؂`e9�"Q��z$	��t5�@O�su��%	�����2���,�W#0��g��]]ȴ���d���-؆��(s���Uy�M	xd����F�=�be٩�Rqn��a�����:�������:D̢�W8��sf!T^�X&��˟�Ё� �0@��XY�Š�LE[��M��k`��e�lVI�Y�+��I������&�R�|�iO$�T���6tA~�F
��"�=�,�AՁ��n�v��u����HCPRT�ѣjQPd=�@l�Ջs.��-�H�*L"*RT�������fl�#A"�lE�>�b
��sfϜC����+p�ŗ����K/<��p��!���;���o1���C�-�܂��a�}?���x镥�2Y��+p�駱Ū������m�e�Lh�T�C�cń����sS�ߝ���2�C>̟?�g��K�(�!q@z$ƕ�_����-�R�I�}���IF$�)�� �
���%tGRH�
z�:�YA�Q���������/E{_�;:{�;:����^��G?y�句2��*tb-{��a��J�q��0��c���솑՘�N�T}R%N@gg'���0zT�׶oߊ��ZO!ft]]{�oܺY��{x�c��]�'��	!W�q�]ݎ[Ö��xdk�>"G�y��m8�5z2��Y3N��/c괉���lB���v��(����q�s�"o���DO[���l��.,�ͷݎ�W�D���׏΁(Z�:�
jkl����r���"�	֗_�G<�!M�֩��e�;��7
��5L��mn��57Ni;�W�As�Eiq>�<7�F~(�h$��|��̹�b���)$g۶mX��:v�k�l�2���r"٤I�`hI�E�*P������@<�T�I�r����Q^;��8n��#HR���\n��Nf���+׵�U��=!^�o�F*a�o�H��p�a��h@yY	�J�at5��/C��L��<��z��-�5�đ�zH��aw�b�i_7�koFc[):��-"�Q��贅OjmS�A�Ҩ�.��$��|�`�|&0>���x��e�O�hw��GL�6����7�-M��B��k���� ��p�]ws����`��)���S����-������Y����������ܰ�Mn.F-���"r4,uKht�7NvsFU<{yP$,]�Qs�1�%s6��ϏmJ�A�j q��nL�2���Ɵt�qc���w�{�;8���[^���c��'�)1���<��xE(�0��
�^9�L����+-�$y�V;U)4��9zIi֯_���B����މ��b'v��]7i*��\����vnkh�䀖�	8ִ}x����"W)�^&���rwdkW�$y�πnk)��-��;n��XL	��x��W�HGp�/NC0�L�,���;���̦-dKJ�n-�T�5uc��ׇ����
`(i���ݽ���7��a���u�000�X<���Qxi��hl����V$��T�D��W[��J�s��:�{2飩}M�mU�9��?<t	�SCȚi�0�O�fb�s^��B��Yw�q6l���4�Ǉ;３[�T.\��d���z�>�ܷ�;�n!K"���&��B%�p�T�k#/����-�	d4i�����]�p'"�7��@���N�(,1�s6b���!L+����/Ť�
+�BW{6|�n���eD#���CWg'J��B�E�Vբ��7��^�u!�0`���G�k�O ����:=#q�t��y�5�{ 	)TW`��Y���Gc�֝<�f5�%8������EaD����q3�7�����b8gb\Ye%/�����v������F[� �)��燎�*�\e��	0g#��;Ѩ����&� ��K�Mߜ�Z�E2��	�䝋���0��	�1ȣ�<!�P��<aT����=����O���=��{}��o��.ybՏ�x���i��)����<���FU��΀�A6�Q, ������5�4k��T�j'��֭d�؟�N����b��󢯯�5X�z�eb�,�Y/Ϙ���q�ۙ6z;��Ld<�|�D�ѡ;�q�=�;�D���¦
�����v3�ίBkk�=�W�X�~p�<�w���c�)&T��܈�[7�(��:��S�$B�|�G`+
�C\��q'��.�N�����'N¢��Q^Q��_�᠙�_{�6mCk� l��v�|������r*���0��n���8ge�-�{�Oq�Eg c�F"9����V��	Ԏ�T:���~ēi��2�(����=�\$�I� � �pՍ��ΉF�[�v&"������0��<�lhB��	֎�e�܍AAF�E�]��rd}n�M�S:ҹ���?.�׎���s-e�?���A�
=���a��j�t�Y�R₝�b��z�^�e��p��t#���!���}ڴQ3~�#	���00��v6������\F8��.I-!V��Pe�%y\����L�L:��k�9���q�E�a̝5^���:�/��-�6�s�+V`��]������ݰ��/������	c�S��څ��(�6"	$��
�*1���ڜt��Ӄgђ�$�gHgn��5�y�,#�4�;D�d��QM.��\Cd���	�R�F��CMu����+~���s��ܿͅy��^@߃'��~�_=��O��ѓ����5t"iP^E���S�j�Kp�0H���ц�`�ۺ55U,I#2-,D�! yPuHh����6�")�H�@<|�O���?��mI�@'ݹ#�2�xh�?H-���C�2*���i}����0f�_}݈�^x��;1�d}�a<����!�q�������#ϣ@��#[�z��Τ�8�BIu�[r8�z���HJQ��W���c�}�a֬Y��¦xc�*���g�%�{, y�eᯫA~]��@S;��n�G��{��H����MלǮ}Cq4���
�ӕ��J���_����>,}�u�\�	,�FFә�L�h"%R+��;���h�"��C�j���g`?v,�Ds�n�2Q ή����P4n2λ�Vd|a���E��� �?ߜd�JxB��N�,�9���	"Y�3��l�/}�G�3pYi�ɸ��_�Ư�' ��X����-)���o`�mmE�+ഽ��a��{Mh��2�� �tH2�a�u�:>N�
30�o�����]����C~���w�}����~�y8�ğ B�*�hom�s���	Mm����C��w8��R�����c�DMu5��l�;�}͔10�B2E�>G��0�ф3w�T\���x�����.��&�+�Z���gK�\�>����;���ȋ�)C ����̓���;8{|��K��K�����=��{}O��=�>�>��qϽ���LF	0��2�u�K��J�(�A�����ʁ�T�ĭ_үRHU�B�M:�@���~�D�����f��?�D6��+/�,@����t�D�a�,�$M˝|���� q�hQi�S�妐��";�s�N�2����HU]���� JJ�f����t�6c�>ӱh�\PȌ����z4l��� ����V&9�Q�B��aaʬ���61�%���J�3k.:�IY��[���~��?_��&"����Au����ה#����">a�m$��!�/�e??�\r2q�x~��߉�����W�/��J��Ͻ��=�x�_� ��o��k����φ?�C��[o�����1~�����݅ի?ńq�1��#ya>�d���م�����0|����{���#){a������J�S�U�\����5t���sMmrh㖼�|F��Vt�v�Y�x�9�zP$d5Q:GԢ��Y1}.��9;	�tC�(v7������ёI2m�+p��}�!$_v� : ƃb��D,Z0m�[���9���0)�ӕ��W�"����p8g�T\t�yضy3��l��]�-���� 5uc�+�B��*<n��j����\�DR�z�����:	N�]� �g@wl~�,w}�dҬ��'�ON�0����.��up��G�߉�͵����OT���0d,����>���ġ�sǜ��ŋ�������'�b/������;��V<�Έj�[�΀ȳ\�BA�f&�t"Mw�i�eAˤ���xvGgZ�3��/|//�����c1H��&.�\���!-����8
�N�Z]�a��PH�-p�N-]W;x�%3۫:rj��#��S\"ɝ�Kb��Q�%x��'�b�Ư0<Ћ��7b��I8���0���,��R4lߊ���C43�y���u+�߉e,"�̢v�$,8�p�5�]����Ox�=~�X̞�/���ɗq���`����O�̈�<Xi�v���_P �׋��!���K@��_{4~���!�0ܮݺu36|���N9��G��8�|�i�˯��	p�<�x�|����5����_��~~*.<�<Dc�X�bƏ�iS�2��ZȺna�����ޅұ��{0����$�22�/@�5�э�I.��ѹ�I�$G*t��� �eWl=���֯%�q�N�@"'����<!����PP�#F�)C����2�]"o(��Oz묞�{��E�}hk���U�q@��&[�{�[u��XOQ�t����`s�f��ǜY���_����[� ���ϣ&�hs�hm���J��U����%/��FF7a�
|^�wBy>Db�q΅΢�����L�c�c���*jb��f��#:H}�&�2;�0�3���M�?��)��y�h�	�Y�.�P�~��/M�aQ����7<1��g�����_�CK�����]�=����<���[���ǽ����I�f2��0)��tV�ƊpZ\��-I����'mSWQd��Z���;���:��Q��k�d��aS�F:�<����*4a<PV���C�,rtf ۠TH���r�ej�*6ܦ�X��q֚�*�U0s�8�q�M�6�M��ڰ�;�����3I��8jGUb��Mضq\�	!���<�C�*;�W�3w!*�&`s}�E��~�Q]^�)S�����-���Ïaݖ]�P��U�;�qF�HP}y�!���GE�ֹ���bUƱ�/����s@sc��Zд��������<���\��s�q�ϕyII	~u���l�}��z����^���xwKV~���z��7����&FR���lmlA����s��1��JX�$Y#H�����.x���<8�fD������A�A!8�*YTy�g�$1����X|��x�6�iM-j���ߑ̑3m��jֶ���wt!���$�et�l�NIjtSek��� ��L=35L�8EaӦN�%�9}=�����+K�a[�n>��A̝==����BYq>��<$Ri�� �|����cI�����_�*sp��7ގ��v7w"C3(�.�?�ϝ��H˝ �zLtc�ڄ� �f�t.��U�����4'�y������\���/3�1@�I�)*�Y�������.7�J䰅��}�W_���M{��%��}z�o�m���>����}�N|�ՏZ���q�2��������8\
�*��cN�mR�Tճ��Mf'Nˏ��($q�h]���F���z:���*(�����"4q<�p�BU=��s�)#^����+�??T�eA�:^��:����#�M�����xbZ*���|�}���fNG_YY"?ߏ��a�֍���M�rԺ'�pn_�T�s�8�0�����e�c Ս;���M@UI#EV�hv����p5���D�Rd���f�vf��))b�%��e�4�S|8.������n����h���3�c�?]�=X��2<�����;�q�z�}�����Y�v�e���gU�3�<��N:	�}g����K�?��=��BUAs{+>Y�S��޴�~{�Y���`�Z䤃)�Nd�}���-��8�I�s$X��{N�挰��V
�a�ΠwL��t (6$3͛,�*,Ҷy��y�Ul�@!ڜ��'I�����&5Ȋ��t��I�#��������=���6��M�O�9�È6l܆M[v�wp�u�Q[U��3&���eE�1��6O�P>�"c�,>^�9Z����Q�#Ũ�ExiٻlM��ڋ���G89�?ۈ_�ϑy8;�9�8}O�D)j�~g�����&�t��r6�̘�p�/�O'� ��Щ�� Aᅾ��S��]�挿�Ջ?����o����oпգ�^���n[���9��7�|,�Z<�Ɍ�k�x����*�hb~����|�E�lp�hԓ$?o���t)Z�u�`Sj_�d�Ӣ��4$��}BU�<	j1���+<���)�4\��*�P��Xɚ��J:./�wv ����,��CuS|��������F��m<���hڽsgLä	���ފ� I��ؽk+�w�b���m����8��ˇ���]����-nޱe��0K��_Ŕ��0��e���Fk� �z�1l�ق����t#(#��T��ǔlXY�My�\=zd ��8��'��eU�����݆��f�7v1;��������x����b�G���k�b�
�v��أ��`�������sf��w�3N?�d�m-�2e
&M����g+��?�Uk�F��1ˋK~�'D4��Ȑ_;�dj{��O?�`�0S���)/�6!�t_A�g�Su���]�e�����D�ڬ!wRǲt?	�w���4ۥ{�x�8���"�$�� ���n��U_� E�Dn��P����ঌqb��W���O%�,U��e����.�>3�P_�/���oށ��V��T㺫/A9�m݂��7�0��ǃHdU�{�&g}�}����wi�{GjH�A�����5���؉q��l��D�$$@!	uiW���N�3O�9O�x��)���Ds]�0h�;s����9��-�5������>��'�~���rV.]���i��9���?B[߈��{�vcsx�$$���;��lMZ����1[��31�+||�3�$"a�����d^~�d5!E_��t
�ͮ+�x<�H���Цۨ?��R�2XpWp�c�Cg��������K��s�ʲ�}{�T�����3�
�����o�����g^z��D��M�#��1��ja�E�b7�p9=��ana@���SZ�e_)���q�μ��K��h"����j�)�-S��v�zy��}�T-�átguѬx�H�:��<���!.�5xvb��t���2��N�a��E���5���'��s���� ]�mdi��x����a\c����e�y�ݽ�ãxlF2�@���$��#���J���,�hu2���U0���k�h��c����TSQQ�p$��~�+�9����"�}��Ҋ�^�M�IV�d�IҢQ�E)�*�b���[o�wlPDD�F{���������0i�T��o���+��ʗ��%�Ü8v�eK���{���L�9���mR��ׯg����{v�]���:A3� ko;��C�ST�B�V����G�y��
}�4�m�^�����m�O��Ȥb���b�k(L�r����')xV�C�X�*KK�FB�5���u��(*�)��v�'�g,��T����y#VѮ���K܌�*�ÐJb�&��� %� bU+��;�&�>�b#� ��A�8��"�R9�L�V��(�������N������Ճ�e��T�T�/�xn����0olݦ
�d���TT���ʵ�|N�}�U��?�dt�����?���p
~��s<��K*�����tW-ӷ&�	��� �Zk�� [�&C�5k�r��e�[;4���uR^V������$�Ѡ��wE!�>Jc780��]��2�BA�N�U�4����U�h�ē/���@���a,>;�g�ݿa�ܯݱ�!�:
��~��t�?��Woz�w��*�ēE0��|䚕\�d6m'�'0<��R��    IDAT������(*�F�HHD�t����L�\��Е�.2���>����x�h���l��*#�A��a��mj�]_M8�#����V�/���TIxB^2Z�
)�I1&��q�H�vvcL$���(��mgBs=?��_1�9L4<J�Hǎf��Ŕ���>���r�h/�x�!�!� '#�X��9׎�#�%��Y�0i�~�~��G8x�F�Κ6Y%K6��ξ1�{�rFg���!I�ϧ�Q|�բ�@���W��4)#CCX,9��v>y�G���7� o�]u*�������vzz�������u�V��`�f����6�z��1m�ڽ���U-�Ar�W_��T<J癓����2�-��v(-������hd(e���X�e��ר3�Ø���B	\����?JRrѳ����uk��X��hbFќ�h�������3̜2��-�������3�l��j�]>?c�%�EL�:����B��fy��)�=Nj,��a�����W,�b$����.�|�=�.�2�PI��TW����U��xu�z��V���R(�L�f�����P�)��G����/�c�΃�������ɒ-9r�C��������� ���Y8���cO���y/�X����i>{�:L�<��'7��G?�h�@g���y���+!��BW��(�1�M'ȤB\u�%\s�*�z�!�z��X(���jW{^����\�af��XRbn��W`�8�pXW�C�j�$}ɪK���ɓ/��x�C���{�=����#w];���(�o�Q����.���a�_��?~��^���x"oτ�X�!.�x:M�n� ѱ1-�3�O&���LEI�3
�KqU�<����Hr��U��C�NN�<����n����r:��ر�;�:@4�`ddT!���1��0�h~������̋�y���Ҋ
�j�I|jk+��>����1%X���l�3�����T{8u�c�N�:���s(/)&a1f�:ĉa���h��A��)ͳ�؅e�a�eWRZ��h8�������9�ށ�WDmu��̜n�N���7SY3���g�~^�e�2�8m$�u-RS6���5�K����s���+���o�-�eq���g7�8E0���A'���>���;��'4-�� +����I#fw�����l464PS�@,�!�HQ]]Ɏ7�q����Y�Y\|�_�f�$�E%{ݬ^<�iZ�&����[�y�
��'�b,�����ʸZ���vp�
�߱4���Ml}c'��z�͚�~�>�}���l�ͷ���d�j�e\y�2|�B��G�<��F�پ���b>�ћX�x���Ƞ�����c�y���o/��g�L?�+�^��Ls��G��m�N�-Vݷf���I��1��+���~�#������.~��_���6]9|�k_b����=u��_x�� D@���*�1y�G�ol��uͭx���x䱍����7��/ܼ�|>E�`���{��?�J��g�8�4HO�vM�S��¦_Mޔ��n��(�����˖�c��T{ɧģ1����fS���E=�N(WC�2��B�ͷp�,v+6���k���n<�F"<��.�u�LY�	5g}�����[7�{d�x��3.��������_�?��~㿼���[�4�[���T�u�'3��G*4B�׃�餤�O&���d3,��qe�w8q��"(к����Ϝ9�E��o�����=l}���`dh�PX��n�gL'n��g�WW�)�a1�$R
��8<8�2-)�r���}���z��b��0���2��Ԗ��;>˂�M��hk?EGw��#�,f7e��6:�Oxt�[9$��@82[e�*S�1�6#�p�k�����ib�|����a�z�l��)4�k&������ws�Tf����~���DJb,5RK��
]lao���t�#����o��� <� �艣���VS�Ѭ9�TF�}$����3��qb�N������i��SD ��0���\"��]o2i�l5����[5w��V�FF��b5�����R;~2.��eKq����*#�L���r���G�D$kb�7�ZW��(S�ʅ�FBg�����QZV���.'�#Qҙ8.����n"������&q�i����po ��L�8�|��ߢ����|�vB�<]}Z��C�ԕ�`������gto<u�4���_1iJ�B�/���{�W����:եM��Rܳ�K�Nb��?#I��*)����ǻ(--��O}��N'����h?u���!<�b����dեk9z��'�x��� _����g.'��a�9yyǻ����(���d���j��y�����H�gІU䤋�N��+Wq�ݷ�l�BA"���1|n�f�˺��rhKGW9�'B���T0��'.���g2��u�ΘO�X���~��`��A�ε�P$+{W-_p׍W,���,������������ϼ�?ӂ~���n���{�+��q��b�A,�55��ճY4��@'�bs�d�L6��@?��rl�l)P���Jפ�̘1����r:U���c�Y�rӧO���N�����G�&3�n��yF�ge)F��͢ӧ�6�DB��G�A���v���㚈��ف9�nOs>��fn��G__Gy����a�����N�fT��1��6fL�UC9�x�$�	�N<��h6p��q*�K�fL�9���3����m��l��U)����l����;λG���=���C��ޔ�U���Q��$�:�Я��� mgOr�'n�7ݠ���A��a��Cш�ҋ�^e1�,�H�v��͛_V�8��㩤����T�Qj++��u���". (霉c�ϰg���(��53�0�̺x%w~��T��PY]�ퟺ�r��$��ةP��ecƂ�^̃�n��nE��(�Un��4V�0���'���'��,_6���a6?����]��R"�(M��y��TV԰��E:�������eU嬼���x�7���E\r�|�g�K/�Nf0��\��r.Y�ď��q~����p�������7���/9yB�$���?��7LgG��!�1;\�1*}6{��4֕�ޑ�Țm|���D(��sq�G׳p�tL��<t�w�mqXv�f�J�JJ9q�4�6�Bg�ӧM�ί݆�k��,╭�y�W��36�hٚ<�za:/���>w^���Il�4����K����-�m�V���u/�����=n:CYY����*W�!Ԕ'�R��\-��FJ5K�>w+�]K�@�g~�&g�#tF�l��K'����wgN���	�;k�+�|znqaY��gu�L���5����+���;��9��L����W,���Y�I�1:Э�N��Ht���ܾ2%i��A{�ĉB|�٬�{yy�N��={V���e�tz?v򬚭�}�]�C�ŬFt�-�l����OR�L{N��c�0##m,��#]Z���4U~��a��bN���U�O6�����?�aFG�p�5$�	�?Ʃ��x��}��=�Z�T��ѱ{��MoπN�c����4e"kV�������u���M6�6����.�t��K}�xN����7��h�hRR��B�E8���~iI�Z�Jt�0�%�����Y�j9sfO#��(�����ب�uYY�J�E��ꡫ�G���n�D<�{V���ڔ\~�e�UW���Q\\DCM5�����VzF�[_����n͓��0i>�u�,�h>W�]�9��駟�h[�N�W�^ɔ���Ҽ��^�}�Ŋי�K/b��y8��ۻ�ٯ�#�5�;����MOkL��իt�2k�t^yi��\�����p��Q͘�Bt��C��YV\����\��=�yg�^\�.?�\���ͥ���u���o�+��W߼��,�e7ȖGlx��m�{�C��Ŝ:�C(�T�8+r�hn�RTB�|���\��ތ�,_��Y0�X
���j����K(����Y]킣#�ز�}�2<S�{��&�J�4��\��a���P
��E�<B���v��	_
��L�q��jHr��Y����=N��AUe�>K��?y���!��k�C!V�5Օ�#��&�+!�\�eE&�����cOq9k�ZO_$��}�9�>�hy�[�XD�Ƒ�o�k��Q^^r����r��F]V�.��'@:�XR�ܱ9E�$V�����
�1��
�������µ�|�{;��}=�1C,�!:��OeZS	�N�H����HG��R'29��e�?�x��.��@xR�e7)ž���E�)a���W�9�y�=���鎫���si�6�~!�	YL����K`]��ɁO$��78�jbR#SWW�N%U�,F#n���R�j��͘�����)��5�ߧ�e�ǫ���j�5�C��v�uK�iٿ5)���w%b��u�Sg�P��Q!{e����c��=�C-+	�1�-��)M�?i�g�E3-2"񨰰����d/^&�\&�8�)D0��i����3��s��$7<2�HhL�F�E�9��xR�G,�`3Q\^D]U%��gI'��}&O���񇼸�F#	,N��	���Q][�>�g:����njj���1i|9��<�ēųd�Z�����o!�p�=�e��6LN�p��]_���b�����9��͛Y}��,\8Wݖ�^�{�h��j�U�p��Iʫ*���R�5!E��/�Ï=ζ={�{�8s:�p�T,N���ʹ��:��2;����y�g�W�=���ۦ7i�J�ʕ�������(&K�]�!�&N���b��.[�D�@4)1�a�KW.��7]�͘Sd��)��{�@,GU]}��X����sF`G�U��x���#��4]Ԍ���C����,��;��`��KlYɥ�'�\u�2�]��7=��n��)q-��2<���0m���E�{*V�N��7����o�>����C:��:$��i�`)��7���k8N'���݁јQ£�-1Ĺ��f��=}n��c&�r��<.{.	{#�y\}���&?q�4��������^(��{}W>o|�[O��ַN�E6k#aR�E��RF�I�$c���Uv$����ˣ]�����^c.�$ª�B��_��옥����{��G�u��p׵0u��w��C%�L��F��R�=^?V���xƛM8�6H���D��:{������Y�,syҹ4N��IS&���윓��Ǽ4b1+�B���]n��2I�����3E�L�3���rn+cc���f5}��(��䑣�S.Z�L>��X�.�#�O��,����.w>�PhYEi�B��d���n�U�	-�MQUU���|��Dʚ���%�=��ͪ9��HkΤ,g9ԣ���x<�uir2��x�V�[�����d^�����(P��F:�UŁd�WU��;ngJ����g7�zH������~�&���^秏l��)R���W�f��*ʝVZj����T����(�{�l;�X����P�4��}{�Q��i|+�L��P�XF�~�l00��;?�!�w��e�De~ٝ,�6���2ꋋ9z`??��0:6���W������n����L&EKC������e��w�\�f�zz����KD�������6b��j�s���,Y�X�nM�V��=ȑ��8�>�1\�<���Kr�{Q��]�JJ�W��SȞ霒ׄu���
��8F�S;��D�/�&k��U���qV.��-7\�O?���L\�b�\�����5P�dEÐ�)/F�p�H�������A�����SV?Gi�&��1�4�������dߤAr��^�3��l����r�N�[6�~x�c�#��1.��m���������<�~G6g#R�(W/�J}���� #�}�29j�kq����US]�����^�ᰲ�Ew>w�\��+�~��>��S��k/^�ڵkyb�&v��ǩ�a�58J�(�o���IMsM�p���>��B.mp\V����.'FJ�^:;9��!N�w��N6��x>YJ4��U�3	��5�nI�h��cu�՟�tZw�B�K��)��͉�����L�qxK}j�bH�����q�t�z�l�2��U��|��^�F(��S��+�].��8��z��5SdXCV��-9�yLfc#���9������"�P���QY�l��j�c�d0Hc�S17��ϣ�a<Y}X\�mv��Ϩ��42�I!�9y"����L��Ёv6>���x��JsM���zm����w?���X�ͦ��~��\�q��4V��}�V�۴�o���+��R�!:����i&������MC�c~r��GS̛���������o��'~˔ӵY[>K�� >���<�أ{�=��}|�S7�>��i!��,1���{۾���޿��dކA�"F���a��)J.+**֬{i�ˑ�Ǩhnb�)x=NEF�bt�9|�G�.Ô�\���f��w��\̜:���j�ʔ�(���v1*�@c�x&���s�t[�W��F��7yqV�~VШ(�fN�U�9����c�C���p;�aÍ467��R�o����[�X�[B�|y��Bc��6<�b�]�����^����,)�S��*Y����93�%k]��<�M��Ұ
�$�A��6s�����OL��r�~ >ƅ�������=o��}�߽���Od�V2��� k�0�҉1���6���FIY3fNQ��T%���O2��	]&�iӦ��x��<x�C�q��I�Օ�����5���!�=I�_L��"muPZYM���+֬���&��SYQ���~X �R�٨{@��ٜp�T?�7w288��$����Х�Y3n�|�$(�h����Ƌ�Z�Κ<���b��K5���:1:��K+q���DKs�Z�F�ct��s��q������[
���l�t,��2�7t�*��J�j��j(-+��'S�L����L��L}Cm�p4��A�`,��EK���IO�ܬJ��Pr_Dlz����2}�$Z*��;�,����]b�,�3�sxK|���P_�:�����DB��/��U���������	��5q����r	v�n�Nz�Y^޾��pT��\B����o�����zr'��s/[κu�()*V��)� �����{ߡu�$j[��3���M/��3c�4��[���<��<���̜9�%��h�l�<v����Gwo��=v'_���x���M�2��f��I�r8���ɯ�عn%y
7#	RW�㪵kY4g>��䤛H%�:w�_<p?�?��KY�l	�&N��o�{}�Cg���|Xr1��T��3���|�n�����|���1<�ZcuX	g3��䱲���|�;�DR����� �`�B�Q%f�T�֪bf4Tb�F����*c���n��lA��D��tZ�����l�˅���7ޯx ���x�e�*��-��
$���5;1��V&����YLp
9p?z�K��?�F5�����W���N��r�~ >ƅ������������g��%3&������i`r]C����SYY����sq��u*+n��J`c*��W2͉[��bm)����<����=���K�)�n�n�4w��K�0Y��,���E3g�RUꧼąӮ�	g�oa��D���guY3C�ߌ^��Ͽ��8>�cId���q=�Ƶ4Qdw �"�m�������dd��V�X����uJt�?����3����=t��l�J6\s�2�}�Zf�utr��q6������	UY�$W�H��+��`��x�g�q�BA���Z��L��[�$�vVKaB�����QI�ɚLiB�}L�������LB�Gւe������[�����ٳ�0M��\�W�la�m�%=E$�5����HW��B2S�A}U�'5�雯Ɲ��}��6>GQi	���'Y~Q+�X�=o�Ä��
�/?�)��:h�.���R%dE�&v�x�ͯnf��E	�q�l�Y�\S�M�����5ki�����������3d��%�_�J��~�I����-�(gϡ�����<��#�<{���j}F'5O��U���mh`�p0�Q�{�Lv3��z�;��g1��j�;e\=+�%6:J0bɂ�2c�]�:���?A��n���nX̆yfnz]5�vs�W���󨢜1�    IDAT����!�6'3g��{d̀9'��yu����F�H��~� ��h����n2���++�v`M��RTY�T،�Ԕ�Z���V�'I�K��� V��OO
�tw�<d�ƔQ���m�ٽ{ݽ��j�&锾i�[��?�"k��>'|#.��"�_F)��#(�4!m���=O�9_�d�W��}�	��VC�����v3���A�;���Ǎo�dߩ���\$�5>̲�UL��1�v����U�~9K]s3gL�xU����_&J!i�J:��5q���G�<��Ü>y��b?����$���?�&h43��b�W��t���i����+YX��%�J,P-f���v��t�d:������1x�)��F� y��A	�<���b�C�%����=y�E",�=���FJ�V2������.>�#��>�4�������S'i��1�����|��q-lzm'�o��H,MVP�%>T v��E>��)MN�%��Hҙ:����W7�E�v����&]i���e�p��/Z�ukWǕ[��*�'�~�(���h���s_�����q�]T���]�����d$�%k��{3:8�֬j���P[FSU��ps�}=ةn"O[�`���E#Av��Ś���`4p�d;���:�D��k�0c�$m����8\6\w��7w��WĔɓGxzӳ���r/[�d��8u���>Z[��PZ���׿�O��O~�#��l�v���c<sQa:�>��αvť�W�K�y�-��1A�̚3�����Ԃa|]��؇qI�:N�8��YKS��<��ttwq��)�4��X���#�3r�/���]��^����ϰjn=�x�7����=oq�M7���\~��$�`8#��b��Ҷ]���vƢI�N?�h��UO4F���!\�056�'#����V��v�q��\y��Jz��K��bl$�.�������1NƓD��ٽ��{�&
*O��`�eױy�~�?�p4�9���~��$o,�H���ڙ1��*� L�D`0������+_�����'������>(_��@���C%?y��<�)�2�Ӛ-9�E��4�X0D���(-*��&���U��n1����hKQ
��
z*�Zs����n������9�޻
���*�����!$�n"K,ge(�0�Ir̫�DF1���he3�q�
�7o����w�U�L���2�%_=o$6�Ng�T\�gKc%Vy�Y�6'�������ɦc\��2n�e5=I6>�gN�����뮻���R����/����[��k�t��)��`���r~��#t������ߓ�	]^�(&���MIY������x���fs�FE�t/mrI�m��e��\�b!o�z�W^��!�9�7����:�>������2�,���&N�{��ȥk.a���􎎰��	���脞˛	�v��T:M,a\K-�E6&7V��/�i��ۨ���{
�9}���mm����*�:U	�ٳm�(��eߡ�l���������_XM� Nq�T;o8��={(������iS*���2���2�Ɍ8�=��Fn���Y�p���49���=]
�O���k/����ͱ3�գ��)&	�˧>}]�����kX�y�6U����X�5�h�}��܋����䖛n��ZX{����`�x]n�)��3[��3[p�Ub5e����9-jݻm�~�{�Q�eE�Z��2�+/YE�ӡ,�=����[ab(�o(����jw��G�	2��Xlk�L��eb�����)2Cmy	�/Z���뮿A��L�p�M���"��	�ʃQ������(�}�!5�!�oU4N�_�ȫ�r�D7}��C��dB�m�!�)y�i{�0Z~_�%`Ǆٜ�ḧ́V,����h���+*i�����
��=����ǎT���:��&�2aJİ�,�R�7 36�!����N'���WZ�e	�kI90"� "Ú<y��˞������C�l&��p���9|�'�d>F�p�L.�W'����h� �����JH���X6���x:���$m�Ĥ�1�SVmV��t�Ij�Y�,����&d��St�حp�U���e�<�����%�pT�.���3gs��I�|�j�y��qL�vS�ڪj�\���q��=��7�S�gq�u���%ML�)�4;���7�����kY;��0��X�8546����E+�S׬g٢	<��6�zn#T�Wp����J;/��.���u�Z����Ù��6���5L�>Eeu����wO�Ԭ���Po�:��}>5����ԵT�w1��,�=�Es����N����`����Łcǩon����K.���j��tq��	��=�>�C!��\v	�^��|*�όL��z�Nv�cv��$Ҕ�p��7i���z}�ڻ�g_x�D:ɭ������2<0���D.�P$��h�qu-lmUe�dfv��K�b#���tXHu��/��W���o�e1s��%�t�Z����y�x�eN�wr��a�\��O���D,H�訾��My���v������7��Jq8L�~��^4Q�kw�>�O~}?#Bh3�Q��_�~;���L�^���?L��T���Ec)Z'N����D6�~�ټ���E�Ղ~���e�E0qb+n��n�0U�5���C~W������Ʉ�R@�d)����/�3��I�ZZQ̈́��gx���9�5��2�A7��� ��� F����?PZ��͚�'?�,SK��8�n���o)i~�BA����o�-���]����	}����������_�L0��)`Ʉb��=gq�TVT(yk��%�T����N%�:Y��L�RХ��+OhA?}�$uuux�nb�F
ʘm�rf�F��$i���@T�>�(EVp���2�hO�ۆ��(���Ū2�M&�������$��F���Y�9a��9L���j�v�d����s�D�ø��0f���c��ٶ�?��A�y#	a�[��9�,^�MI^����U�0��
�ӎ)/��F,��xv3�
��@ Hy�ǿ��e���5���U�����߯�:�	yMȄ����쒥�La�gIFٰ�2�X3�������`5SVZ��}����=��Ń�W�T�*o1W����2S�50�Lw/o>A�p��X�Ԍ���1�C���b�|b��V�(��{4 DH�g;{�Z%��JC]^�'��w��H:�ۇ�W����t4N]e1���x�V]ό��8r�f����H��$cq�`+|.��kH�ի �L�<������c�|sQ�Mt�ʢ����j{1dMڸ�76(c<i2�3�X��{{�2e���<ӔLp��|��+��l� =�"�T� ���}�e��>#�K3o�m\F�⼰c����$�-9����X��N�z{��͘��Z����7����FOm�œ/�D�f���I�)ĒM �or�I%3�	"��2ԺlT8�d�Az��P�����s�p��ex�����֣�5 ?_���68�s��	6=��2�%xf�ٌ�:��pZ��:�c��+H��ff�t��u�^�W��n�9
j�]�^�"C������]�`M��"ݸ����Ђ�'qm��o�#��z��{���W�y,���(�g�#�$Ę�0ALe��5�f�ʕ��5h�N�9C!Pdp��Y���?��|�]�viB�h��Ϩ���]�K*�NB2OFHl&;��Q��fsI�6y���Ql:͚4eϛ�H�,����q��V���&F���>��pNcIs�����V�g�������%�B���t#W�����|��_1�ɑu��7g�*��d��"�>'�uU�q���}��I���Gl��dm.�yY���43굒�.�v��HcR\V�����0�H�p4�`OV����5���sj��r8ȧӘ3iRcn��J֬�����ع�Vu-,Z� �^�v���������/>A���'����m�����3Icsz����_�T�|V!�����S/�y��
qOlk��R�h���$.����2ܲWMt&��!"0m�:T*(���M-x�N��
Eb���buz�J��d��^��-���\�)��IA/,f�kꔤ���h�wd�aI�9����dܸVU���n 92HWG��b���cIE����[o����*����M/�ȧ3L��f�Vl��J���3'5��zM��͋۸���X\%�#W]�u+�QZda�['����zI��L���}�Q��ṗ���Y�|%�V���iVI\峥%q�dӵ���z�-v��wTx�LllĐN��١h��p4����Y0.V��P8�ix��.��Y� �=�<p�ǎj��\�9.��~<����^��ف0�#�dǐ9����ҰjQ7�鑪;�g �����]m|�fC��5K>�~N��?����P�3�a
���M�_��������f.���9�ᆋ��ˇ��Q���R�2͍B��ٖ�.]���� �V��I1��{��̙Ӵ��ShRY�n9�����\iq���XFY�6�����G�_Sf��Yɛ���fl�+iq𒒮�-�y+��ȴ.4��4����hר�d*�0��`�	n Џ�fbBe����i*5q��0���/�I۽�S��4)L�a��VPYV���g�`BK�Z�z�~\�b���*}�(�D�X�@N|�M��]�����d"�����±�ơJ���/�I"� 6�YY����-p�s$�����2�/�*Fx#��d��;b<����{�p����!�M1�����Y:w�2�Ot������B`��ɛ~��B��D"Jø&�.�>ߒ׻������ �m��xȤR�n����`�ϫDѵ�aptTe��5�x�>��"���ct���ُ]4�Fc�Hq��=�)��b�h��i���"V�&�����~F���'�b1ZkmjQ�]I�������KC`�bO��z�LV-�Mqi1�0�lz��<!�}O��������.�;��C�`�Ǐ<�#����)�	��/�#�*|��h;?��F��f�.�Z��_�<U^�6�Ol�Ƴ/�ƭw|�ŋj���!YC	I� �B2K���T�$����D�����Pc�!�X @x,H8����Y�g��:NWc�1��αٝtt���٥b�4(�{����N�I�=l}�8g�B:�gS�<	�]Hq�#^��[,� ����@J�b6as�1��8�����f���ږ�.@�:E�BA�ӹ��wr���xj����I�2Ix"�uK�QfIcI�!v��D,��i�j����	�U�c(�0�XY�#�x����n�ϝ��\�����-�T�`����+��%�̄�*.XI%e�II� Bs�x��Q���E�Ҥ�a K�`��LsٜNlR�� S�O��R�mB���z�kv���r���_��	'N��ûM_$N,o����q�u$��t�>��%�]g{�H���2�[_�TI_�|�a:F1��mn��r9ѝ�T�&���dBW��h�h<����`�I^����E#��5�u����6��')�|h=fO%��6�����u,ϼ�������r2k�<::�ik;�%Ý���o���{Q�o}���m�=��k���HAO'cԶ4�p	�)������n?��,+	"Q"�M�Y1�!��zmu�2����B
�L��P�/��p�*B�RХ�1�MX΂��Ɉ�h"�˪�On�N�$�p��AsC#V�:�X��8����$�9
=�A ^AD%a�z����������D1ܑ��[�.gټ�Z�F���-m֢�.Y<���.!���O:c��:\~/a���x��W7��C�V�[�P�~�{����YH�#̪�sח?M}�C���x�����򵗱l�Ŕx�J��%�����<�\����Cl~�	�n��禮���$&�M�tu�Z�b3S]WKm]�zwC~��($;�����^���g����q��)��2�9��񮀦��y�N��.�Än�t��E�'޿V��L�ٌ�`H��7�+�O���
����P���o��������>������x*�%Ƒ�jZ=�>cS&Y0��eIdr�W���ۆ�뤺�F̄Q>��C4�]�*a��c1:::�L&p��5�ؼE��\$M�SBI�8r�J���0�'$��Jn�)ВC$�v!�I:�H�4�L/�v�z�@��L.�	f�������~Y��gt�݄#��˷~�+O��l�'�yF��,n?K��`��b��>��[����´덝tw���h��y���?�o7>�lWqޒr��"��@�&���c�$���oV��ф���""{A Db��`5��!1XL454�Y��rزq�|�/�Ϝ�S�i;�~�˗�d�̙���λm����oj�K_�$�H�y���<J���ԩSq���Ny����"O��BoϠj�mV�t!��67����IB^&����٢�)��//ĭ|N�T)��CiI��0SaR��	��p���{��x<IgW�]�5b�$(����@�b#d���b���آ�V�L֐������(V�f�uG*���	ͭZ�m>�~���~���a��� 0z2�u��#W�%r����/���b�a0�l�<�.�OM��s�#
q�6VSZQJ�d�{�x�g���[T�G�o׭⺵��T����{�|�\Q9�p�9�����o��#O%���ͼ�m'	���S���j�R�ci��9i��dL�i����~K<8�)j�n�"=5pڅ`����O?�x�����X-m�C�}��E��SQV�,���f�q�{�8��v8��g�h���Y0���`&#��tsa*��]͓�a����P}���8�6�4|��+g|oC�A��^W�BA��	����]Ϳ��ړ]��\�s�Ra\� �L�gQk�l�l4�Z��1��be�����������RQQ�ӯĈ
�]=��A�������t�2�-Y����������s�R�2�ۧ&2�f�>g�P�@�܍f�0��Ss��LF��*����Jb��Ϲ�-3�ᔤ�t
��BGO7RЋ�،y�.]̧�]�-+{`q�+ؾ��Bgg���|���s����ƺb��zE0X��-����;y���H &#YL'eU����{ɦ���6I�tw��0y|k�T�˥�N��u2�%�xJJ4--���}�Z���j��<{����{�D�BnX�a.�K,���(=}}��_|��3�Q�ĳR)%Gui>������(�pAV�J�#MX*������UЗ��Ke9�ގQ4�����ȋ������1���>?%%E�wڢ�4+��.�L&�+)�Lr�\�j�m�)0����.�:��*%/MF����.����s�*I(�.τ ª�Ҫk�TPʅG���R\��ɐ�`I��q�"n��2m;;��Җ-��m3�M�6I.��n��7Y8g��@�_�;���{JS=�_����b��8�?��!�[�������ۨt�h�_?��'_y�ȿ5bE��I�-o�*4m�(G�����-JmF�-9��X�"��G��TWa�����%�����񨉑x�}at,H4+X��}TT��9����Lg/���ݮw9t����0&��tF9�h�q�x�jI5��2��K<�ш�唂���ʟnX6�Λg��3�����_��?�$���^j}p��Ǻ��9	I�q����H��H��A40D`8��v_I���uLƼ2�SUQ���l:��2��'�_���0�C,R���Ì���o�>gD�J^���+�u_�H�1Z�$�����f�g����χJ��X����+�E�L�L"�;�	�)�Jv9X����J��AfiQ^w)W���FxZ�>�W_}�׶����-��>��%P��%���ةS�{�H��n�I�I�3��bV\��!$�|�x6���%���ۣ��d�Vrx[�Z��%��*�k�Y4�V<�m�VC�勗0�u<w��ǜ:~���
�^��cL�2���O�ke�.y�F��DՂ}����g�1Mb���:\���٣�E`^��sij�uO,r:qué�v��+�laB��3J�3N�q�q5����㣬�B������B�Sރ�S)δ�U���r��\�	j,�    IDAT��+ LV���F�\��^	��]��=$ծp@m}mv�.Ey�9&���n#��@� �}N#4���&"��3���v������%P��2e��h�\c,ˮ�����{o�������ӓyxz��=8�!&H�8!$"���	P� �d		"a�D;�G	B�Q�q��q$[!
x������guUuu=��<�F�u�l��vUߺU��o��������o�{�{���Z�Kg6�HJO��>���.��勲�d����~랬�JV�����e�JD�A>�_~C~��?+~~Y
�ӽ�"��'B�,:A��}�����ҍڒE�́�H�Y���(�> �\�x]���e�d��ɌJR�2ۊeanFff�P�E�E��;we{�'���raeA�f�ew[?��}��������?������㽾�^ߔ�W_�������7�ʍ{[�ܴ����T��!+u�0AָD
�`�"ͣ��N�ݴ���_���?�����Pz6���d���͗��g>���}����P��#�I���to}EV/&�jư�.J�{�AsOcE�c<�^Z\P�NC-���+S�B8�����7�|S�Ə�]�;��W��(s���K�G�.�?/�sӺ8��p�D�te��C	�TZm$�8��k����󠘙Dc��a���=�j%�=׮�c'�[6�[w��ݝ��s�:����̄T���*��-i�L�����d��c
\�����]ռ�8c���7�.ۏu�;FRD#ǉ�9�gw#9�zN��u��G����H_��w�J��Q�(.�Q�E���f��B��c���ܿwO�66uⅠ)~]��t��1�g`����2??����#��c[�]�R���`Xȝ;���L����\�����̆͡��捷T�*���/���������m�����]i���B�vG1�cuO��!o?*�)��KwЕ���?�t�#מ��φH�s�<�[��]��4�tL����3=�������'������*�K�$i_V���cG^�c���y�f����mo�>4����L޺�._��dyaA~�/|P����֮���%�y�5����t�������¯}N�rw]�hZ��Oub��?�y�3m��ᓿ#���_�~�h�ĉ��Gv@/!8i�:��duaZ��ܒ+S�`2MumyA��ֵ^&��H�#���D�nj��)�����~o�Cb����5��K/_��G;zq��5��/�._��mY{�X|H���9k$�NS�B�ݢ��O��+x�$�Bͅ`�O�t������\E�{S��Q�GQ�
]�������ү�ܗ��H��Xf��[��=�+{w�&-?��O\!�磱��(@��]Y^R�����G�J.��߼yS�wv5����V�z�|�~Q����n45��&!T�s�/��/��v�R����x[TL���
8����R��S�GÕZeTTa�bȡSZ@)	�f��锡�F�FAGBT�C�A	����޻�Z���:8�;�g�g�Â����i���o��|�G�QcHuC1�C�x��T|��ѵ���4y������,ʧu�;�����յe�A��JCqV�'W5��]�-��^#:�� 8�T��mS�rs$tðG%�U�-�V��pz�ϑ{�}_^yY`��سR���5B�Pv�hը2�U���4���{A�@��ފh��y;a4�sߘLw�(k�	W�l}n��U�j�pE�E���H���рs�X��d�������-��Q�IП�����:t,��a^�JIh���S؇8����Ov���j| �@0ce9�d�f�U�m�U���>wD�T�5���OnPTm�Gn��@�
䥭�+[����R�N|p�u��Bg����~_h�7}��ʱ�@y�m�Ψr��	[��7��ߘf]�)��Γ�c?��ӝ��;�Zy��g�,v���������#��D�wc�Oj�r�ɦ���������٤�Z��,�%_U>��}�hԄ��%�Nd�)iɺ��t0��ݥ!pp��[�,�M-�vƧ>��q�&j�JB`��܁�/�s&��C��������s�T�rO+D�H?�ӣػ�*�c�"$g]�P�o*��$MT�jbx;�u��mt�ft5�s���Q��5����w��H';�ܘ�=��W>9�r]޹�$�|3s�U}о�5M�`=r��A��s6�Է\/];V�뫜��W������6_�9�����mΦE{�s&.h�#���M�̗�N��@
�t�lU�)z-:�_�0U�>��I��SuN�V��
zG���K�b�ӯ�hS�Y3�dAgD���%��{)�(��7z�g�Vq� �!�O��4ɬ��=���%�{l�=������ݙ��xq��?�+�� �]��m�VY�����5���Ӟ����>�6Hu��� <U̸��Sj�O��ς���ٶ�CV��F���?�-q��X���e�I��W~��;��wi���t��:���8y�y����]j<�=v��BB~���(��稜����	P��L�Ӆ�4��o��F��B��̏fN�F�p�@��!^Ǻ))�#aLS���/��x��<��E5����$�����er���_���mִ��)�몋�Ov�	�,��+�]�k|~"s�t�Sh�y^��-2BA��WAk�ݒ߱0���$[�u�+<o�gߖ�qTE�Uf�T����l�g���Y0�!vM ��y�OI�W������}|Է������:267#�8.)�4��������Լ�Vf��.��b0ߊ�����]�c)u�KhY��Z�d?�O`�95��-<�qJ��Օ�L��\��`�C&��x���a���f����~����?�"�j���W��R[*T� �͸��h0���G}~/�}��
�FB���~\U�?˺��~Kb���	�+"��&��^�>>���g%��dξm�p�j�צeX�5�Q��r�x%zjv*�V�DȖ�9��H�H!օ����*#�N������sq�V�Ј�+���d�3js��{����hsg Iؠ�ݣ����>�(a�6�q��&�9����z��I���� N/��*O��9ͤ�������kq�$_��mQz�nQ|��Ԟ.;�X�����W��˩������Z�뀚�r?p�'{�k���ZG�J�����$�B���VJθ�u�y�W�¤rm�������v�l�R$��p����S!8%%�O�	<�6��j���1*��:�e[�d�<"�� �L���澖Z���wŇn����\��8�Bl�]Tvizg&�m�	<4������DU�GO���V���i~��.��'D�vr�|�P'���aq�ն��	W��-6�NB����ZR{��g�߅�^��>v��jo�a�	/�ˬ�Jk_ �.։����w4���\�"����a��OA��^_���%��F>��U�V7��?���d�)g�鷢�
�1�eږ�Jc���0�j;Ծ!� 8Μ�˰P5&�~w��!z'>���i�H���\�P?,N[W��>LW����^�J��������|�jSW�<ÅK���C�B����������a�W�+	�\�_�)�6`+��t���ԇݼ�_e�3��R逡�]�i�]���dYq�lGOiHᯒ1qq6����ǭ�¼���8������	ZՁccc	W(���wM��`F�o|Eg�,�%{{ K�9Guk4h�ÛjČ�giF�@� ���hUjd-Pg"J��9Z�60�2b�A��YN�Κ�(��Y%�;'|zo�K~�(2H��8��QD��6r��g�r��.,�����_y>�&�e�0����ad���EL���=��eZK��(�㰌��`����ɝ�Gg������&�$\Z������TFͱZ�V*����=^��;j�|��<<-jA:Ң�-���p�r���R�Tk�ɞ7�5���QOA���q�䫟5'b3{�={k��Sb�
!?��b餿5��OF��8%R�$�/iAwgpO�?y�oW�Tv��آ�Y���uv�t����V�JmŒ|Xs�^�wM�m~�+���^���[*�/�ɼ\좋h:bC.�J_�#&��A�l�[��7�W��6�<�q+�
�j-�Ъ���g}��ӂ$]41���#p�`a7��r�!z��@+�ȕ�jv �F�C���~�
�������B���#�	&��B��/�O_�e<�O�W��r���D��,�ȰBat�&�~��nq�l��xz�.|g��Mu8��PK7��q�Rޮ���M���M[I8/��R��tV���vzRq��4~�������䠮��R	��![1��죈���0mTq�~}ꔢjԤO�SK��ߧ�&�w�`����uXx�Ru�(-�M~�=���[�4�3ǉr����H����^<�)dwq�K��A���\��OO��W����aH*�e�x��ɪ���hІ۾�}]E��2\�`g�|h���-n�O.Pw⸎�$d������'D�	�y�E��ؑo'%-씁�7c�ֱ�@?ȧ> �V��\��s����6�x�9���uv��Dq���ۿ/+��՚j�����ќV�8��}Hؚm��ih6T�&jt�'���������P	L�ɔS���r��ǳ��1h���v��[m���E�ӯ���c���H4Yv�ǭ?~�j�|��U�^H̢a�T���B��\�=,�t��EA-��5�LF�}nR�� =(�!ʫ�qW.3��s�fX��8��跅$�6}��/�QK��hI�0���ä��8�Nlyc�W���L���IP���*�) Uq���N����T��âitm�
?S��R5JH��	.,fxi��4���g.F����0n�/���p�"�f67��Y&vD'~F�_�+�ˈ���I�AK:����D}��i�
�)�J�����G,�þ���61�D�,��\�,�\̝8-bQ+7D�v��}�A�Y�@�y�=ˠ�c@G�����]��8ęĭٔfd�Λ���#y�p���l�^5X�>�D�,�E�Aj��>���.��t�k<��ْO�X�g�"���:1�)��tuh��z�<8��*f��L�Զ@0yx̾h�W�1:+����ȥ�ƍ��+G�]ӷ��:eȸ\j[���PK?�v��(��d`�$�����+�[�P��L�I;��}cm�	�}�������b2ݧ��#cX��#��"s[�9M�!*vq^�xd�ǽ5�3�-��!c���#,�w�����U�p�覶>�2���A��[��S�r��ꓚ:����H[�]���j%������Pս��=�6m?�qW�ƮFѳ�1ޱk����s���+L���\m�
��=#���e.���"�䪸c���P^/�����ޞ����:\���!���(�pS+�ȼ]]��Xe�������$3Bνٴa�vq�l�z$j�޹�����l�9̤f'ٝ�T�!�����_#��ZD�,�Z��3^:.A`o��Z��(��gy��,�$��wuɎ�����A�IC��q��@O�w`3�R�c���j!ؗ0�N��T�*��Z���IcnT߅�w���|L'�Y{���x>��Uy\NT__^����A]F[�@��DOD����z��n�8����Z�<�s�EA������Vhٷ�~�ԥ�W��-���2�_��Ǣ更C��7���@�h�A���6�^2
&��=��k�If����2�i�މ������;1ǃ�͝{%��w."���N�U�7�"�����B�3-B������3T�1��b���B�]�G����2�k��r��w/�cu��xk]�ޱ�m��8.3h�c�*�C��!��e�oc�QT�l.>����/�23:�8��ly]&�S���ls�N�ݙ]5��G��0���2��԰<>P09���pH�zƄ��M���_�R�f�q�v1�ſ"��L���Ƙ-�wKIh�]����8���X�jϛ-����y�L����#��r����Ci�{M=��Yg�_��*ߧ^��K��+	wGl7���u	�+�:~�����^�]��8avf�+� 5�T��Q�1��.
M4��}������"�,q=s�B�un�g	����|/�Q��|�lV��!�{��|�Ʌ?I+jf�j���Z��*��.�>�0rӿhq��U]w���A%b(C�s�/7�|�R�{vx��j�z���c?�+~��-H�7*��g-��Y��GV�����Y��N�E�B���4׊�"$�sE+����k�o�&�h(�^!��bP�V4"�G%�B�����Q��p5Z���2����h7�*��P�]@����p#�ؑ�!e����Z�]�W��7�(�Q���PoO>�N��#��o��db��t
V���{���r11s�����LBcĪ��Tg~���oŊ}���M�<�n^�������n-�"I=ĒoS}��~	2��b~�  ����Ӳ)����} �U��C�l�~��	�3VI���x3���	�1-����N��'
�z�����3�^ȼ��__,P&t"����h� �b$#>޻�+���z�DC4GF؁��v�D�G�� �kOAᴷ�iB��O)���|��l�k]���k��K�ǉ=]2��P��0������R���
�@m�j��pz��\�ݐ N�+���6>�8�k%�oS���E�o��ϾE��pt�+Qġ�<�y|
�.@����q�_�'���+!�L �^��_��4 ��)i0m+Ї�RG���nk}+�Ā��ű��_{���g�*�C�Q0��T�Ʀ�Ac޽`�XDn.�h��������u�8����5bۚ��+־�W"�h�U�U��sL�@���/JO���3@a�a�xH�,�'��D�).lM�܂����T�{� �#�K����!����ü����u�d~H2��gr����L�}+[{�Ds��$��ňA�L
����2��I���@�:�����H��h�L@l��o�  ,��C�W=�@��y?����xh	`}Y�9��7)�Ѽ��t�o���sÈc���Z����w\UG��ܜ��
	���m V���L��15^�I�a&��#�P�}��=\�Eu�ap����<�!ȑx͛�����Xx����=�AB;QFA���w��M��%��@�n��ś.OD�YbOd���\�7�B�fbH:xA�^m��b��j�](R�-��y5��'Y,��n4p��bV���y1Avn=ݔ�#(��	�X�:����:���?��+	}�N�V>���k��G�]J:�M�<!�[��M4����i<I��H���	��������4�Ԣ���? |�.��J�}�mK�~y����\�y��P
z�
��	��Ra@�
�&��'=i�r���_˱��B���|��!�h��~����4�G�}]�0��Gw4����~׈լ�\$��Վ1�h+( ��H1����oI��o�-��F�(;��؜�^ᷞ��6�^ub���,�p�EWX� �@M�7e�'?�Y�D��јox�"��hL#%gY�Z1ӤճIQ��w�=�"{
��1��R_a�w�-R@��f��H2���_h7·D
���c[�DƐ����A9�:��2ꖟ+�QF��d������
QD�3Z�{�Y	�V�:7��O
��d7�Y��j��!�3���dX"�v}�a�ù���������"��Z�#�]nx]��kЇ���F�M.�6`5�]X:oؑ��a��0�J����L�D�@4�28�-�xD<\��/q[�*J��W�k��?3��jN��B��k�����PqqF6��#8ch�Yd�|� ?�Ua�D�+A���F�~wG�_�5n��1���{T���C�~�۳��c�9R��!GU$o��(��u�V]�ǟ�f-3͈I�~[�@d�0GJ$'�r�����ԒUnNt�����XX����C[��>�Ԥ��1�Ⱥ!8��妌�(�G,YB�Aߨv�n����.�@�v��v� 5@�D_���#)#�4g��p��d��7qo� Y%27>�gK�s@�7M发>�K���wg�a�Ӵ�3�B�̵:����Ԧ��!�ȉEA��}^�W�omR�����f@Q�ᐋ�E�I��n�2|��{s!c��R:G4�:�H��['D R&N;�ޥֲ�Ls�d[�������a�����0����i��08�<�v���l�&� ���E*���x���G8���z��x�ȷ6��4Q~� �d�"���\N2������L��r�ۋ�?�����W$ОbDb���ԯ������te.�e޵��ؾ'-�A�:�j��nL��d����BGI*.�o���v���=�	T?�FO
�/���Ȁ= �vV�5����oB�A�s��ѧ��!9\$Z\j��5
_z:�+1WS }�v8ۭo/4�������d��U��� >nWo`Q�%Q��{{B�F�0Ln}ϱ�e?��ݮ��6 2vcD&HX�rd�#6����X	d�z#��(��Q|LO�`�)���k �F���萆��X�M,��A���lL�trf�D�H��B�$p� ���D�����-�嚛�kb��C�K�G^��T��q� PK   ���XZMZ��� d� /   images/c9083cab-aae4-4f9e-a621-fba1f0ef8f4d.png�e[\],<��;� �����www��www'�ww`N�ܯ��sշ�a/��Z�#U�dѐ��  ��g)U  Z ��C����<��  �I��{��y�V�oD�f�M��;"p��(~���9ȭ$����+��<�1�a�H�W3���TTT\�l�a��ڧO[T	�M����=m< S���ʭ���cvkb�f���T�b��/�G�禈��
8���)|ِ��m�I�A��������A�� t��xd��W���{����j�fG�����m�x�߬�=d���u�E�}�e��1ki��i���/���s�r��l�_�k{ߕ_g(���Q Ó�$�\|+����K�% '��9^���}�ݡ���8��C[H��廚��~��`�E�?l��[Qy��Y�߾4��z�_���>ng�NA��97���m-Q���9�}C������G�{O���#��M�����F���I�[���������� �2r�H¡$�Ӄ�ѕ��V�	n�uQ;��(_9���x׵.�=�r���g{:��{ �?6n��-���������ýg���Rd�����8����{�����j�F�c]E�|NS�'��l7��k%p��#���&�ߤ���q��s��Zqy��޿t��Z�������0�۫6��=x(��$�8
P����1��z�g�!�g](X9�.��t�9�ݭ�g*- :fu�yp��d��Y�m������+��8<���aZ��5����;X�?�7���2�E��lݳ������eX����*�$#˲G�QX��Y��#$-��I�h�Bs�~Y��߄d�g~/�-o���O� ����������*���h=r�M��p�p)�� �Wj�׼&]��O�[��T�=T8g|�Pf�h � 4s1'uf�����k+	K1H�Ԫ-��3Uݶ_�eɇ(�$iZ��F��&�]�����,�zȷ&0	���c"k�bc��s���^3��v�G���8�Wm�=
 8	��nIJ��}F�E��1��j$���ʛ:َ�\P�=.O����B��]4wB0>� |<�Yj���0���ͺD;A��R&F�_��چ�ulB�N].�r ���9~�	��+)Zd}�&Na�`��O/ZL��T�F����a�(�$(>n�Ρҟ]�Ǫ����Z����X��Q?y�r�.�p~���� y��b�p���;ӌ،���}�e/������BS��P�h�R<;�S�6l/Gϋ�G�=�p ?���6;��Պޖ%<��w�Ð�|� ���Z}MiRR8PU�:��[��>``�m	dg:*�E���~�Ul�l[����(��;�M�WNї:�
��E��W ʓ4�� f2M3_'�P�J���}��1z0sc�x\ Ne�X<�Av�Z{��Y� 0��k��Eը��o�Y��j�x$��XPy����]Օ��m�Ҟc0�{�^��� 6n�� N���H�(aL;	��Y���6��𣴱���H�M��r{�P��w-�������?ygz}���ܾ{��Ԥxq\ڀ�-_�1H�y2}���#\ۡ\d��!8�� 9~n�������� ���OD?��QR1Q2l���$�X��aq�RCq���0��k�B%7�}$���n<_��رK����:����p�u�	�o?��b���:�1�o�׶5xkͻ��7��h���l��tJ4|�� ��N��6�$�⥓�P!��$��=������C3�A�ʥ�"�~���rr��p�/\"g�mIlb�L�p�C�_	1�U�Ӛ?q��.��7�ܦɫ��9F��B�/ؑ:��]�f���<�n`(lR���s	xa�P2�P�0�<���lB���3 �-9��G��1Q�%�@�^�H������;16�S�X|7�TJ�^�|�l>��I�),��փ�q�F��R��x��'��k��UM��6H_��X�>���v��ů�Aۘ��U��8_�cTv��C<!�ӯ���ڹ�Ua󗊻����F�����ў<�ڢ��4%X�%j��{��\S<1=C�+D\�38Jv-�oZ�TQ����4�(����T
�	��#���.Oi�R6Ѳ����4�\9?g!3#'K��#[��Er*7����w!���`�dMwv�W�_�Ʉ�߭���+K��-�'����n����/�B��T��f\�kqӇ�Yn� Llb�@lS��gS�����s_�S @�M�����J���|Y�����g[u<��cBW��V�G�*�0능���,�}���U�Gp��)�κK^�6��?
`�G}5��kՆ��|O	=�%<"�����2r'[S#�e@&�V+� \n��>K,a�Ho����:��_��	J�Ψ��9S=���x���/���8�mϨ�8S�fAJ�E�,cW��٭�룚�'�[�=o���{B�U���X�i��+8��<.j��,r�g�� �qzz�ݞ"x�H�`����p�1�0������?�m���7զDD5����Cy�����x3�k15j3���� 0�:q}>Dq7һN.�A�Q���%���i?��]�ޘ��ؼK��<*�h�.���'��%Ґf���T�A�ov� �H	�/PYi�qJ�d_:+�En0Icf����2ҿLg�{�(G�B��8?݋�}�X���8��(�?�����R����}��%2(�#E�`�[��t?�]@-$��{����<K�X�&��ɉ��|D�ۼ�����+�cթ���*��ٞu���N��
ܓ�^'���IP�p�E��G!�;o֔�4����dTӛ�� � �;�U\�Ҍ_
����}3��)/`A��j�n1ז���Wk�"��&���6�(ڮ�N�9Rə��ӹ_���V�1��鰞~��������>�?=8Z��m�tT�7�K߅濛Z�,��0���U���d��^6��~~+��_�W�aŏ��@u��F��z�Շ�����1���$�R��m|�J/�a�
���Z������V+�H2�K$�Ѹ9!F�ܪ��{o:��I�6Lӑ[%���bj�z�a˛J�]�TZd�|�9����%}/C���/t��k���jQp$�;gc�*�k��:�-�k� 4r�m~�z��C[�ɩA8��	��WhN0,R I�}b�\�!#����X)T�c;�N�6�!N�0�c3�9�E��D�� ���0V�`��JQlL�e���P|� h#���;�:m�,41����/!)Hy����q�╊dC��O��6e/�l/@��O$�ʝ`
��nѻ�M�*2��\ǿ�{�r�t*��Al!ϲ,��ga�˟z���M����H8(�]����Y����;��L����z�r4�i�"���F�r���x2ꀦp��(��(EK�]��n�b_���Ůә�|<����eg�w&���Ju[�9�
�?��4�MEs�v`I�=�_Bj�������j��{z�6�x��<�2(n[���x�i��>��<^�LNW�7 [��c �j�ᾉ0aRB�ǓH�N\u*���x���i8�03#��y���N�!�/���b) "��H��Tۘqd(y�yNJ�Es�6�f�k�XU
3��M~�	��R�4�W��R��u�D���Ez��ᔋ(b���mR[�̂wuRQ��\x�nl��u����᣻qoY�/������V���O�/7l�Ğy�����]�f�:o�u���ɺ� b ҏ ,$��|z>%'�,���A��!�Q 9�pb:xbt�]傿O�����0g4������H�.�"z"R�{g\Vg�36kH�J�Q�:�+�_t"([��6=�>$�f�B|�fH �	�"�o��׃˹/��2�����4g-:��)�<�Aj�rޔ5��>~к@���p[�Y�t��!�$��H�G֪�,H|���)ձ �����L��.g�5aw���3���ޭ'�b���y��R��Yۭ���IZ�ӆ���Q����Kp�k�xF���;-�jN�e��t����Yˠ��b��
��o_�xS�	�;�}���׬�o�_�K!�A��68�S�/���o���ݾk/~au�DmC�7���1d�oF�(�R�T�0���������E�v%oՃ){U�;60�3'u��þ�`$+Y�]'$}�*���SM�(x�^�*�
�k��NRN�B瘟��-�{E514���FR�8 %�gϞ�ςҫ��������n�=_/�%�Gp�Z��;���!ط��|�S���7౬ǥ�,Bt�Q��cP�Jn��`��W "4bC��C_�a�uR�2FHqh! "�5�yi3�N�5���0�F^�y��S�*��b��Ysx4b����:f��#&��&�b�:��)ՙ]Z_&)c��95��$���ј$&f��%N�.������]j;�K–���˷~���g޿~�S���/ԙ����n�B��z��r���h�Me�{~��Rd����Λ2�PD'P(��}�-�����Z��Tv�6�~�6��j��%�#)9�Y�	�&��1K�'� �!d�Iе7b���;�����9Ug���儯d�&ל�1?�Ƙ���jZ���l<��>�0��$��E���6|�+e� ��z�+�泓%��p�I%��z����jqhh"j���|�����@�ܜkH�5>�_\�Ӵ���z:m��;A���y}:��uҚw����+�	-̖%�Ԣ��,��I�� �T�F��}��C�3�\PѪ�@�ީ�!qG�w��(�?/�3*E�{/E���K���rE/B}?�7��ʗ3"�;E��U��r�J4(�w�

�\��n��s)s�_>ih<J�-@s��1ѣ�����ȩ�݃]	�_����ю����io=���� 7=�����3	.M�OE�e�W�ZqD�D]�{w�)V�,�F
J�$��jڡ�{a4�f(<��p�y���9�`��Яgw�쓳0�գ���b����̧�������H�����R%���[$��{����b0���,M$ނ���T9vam�MUv���ڋ���5��'p�v�Y�_ծ`\=��̏�>ICihw&$��u嘂ѽ<N���g��z�
���z����L�3{Z0���,5;��`���
^��3rh��%�')� pUL|�N4�9`�;a�z�OU��}MD2�&��^'�Cm�&[Iè.��m�t��h���Ŗ����II�����F� e�=H�Jꗯ�o�Ԡ��'��^��s<��I���d&��<��|�&3w{N=�LW@��w������ɛ~%	���g���h�Sޔ�5�L����	�[Q߁5��'_�̕��,����o8��0kF�s��-×�����7?�*��$��톇I�HH�j/:[>�z�^c�wk-���Sw���i3�h�ZO+�X��23$&��v3�(�E��D��l;G�=�_�~(H�8�\��\�;$1�%z���Ӫ��X��)���(�q�cK�K7��y�JH�m�t�O�(
n:����A]w������dCj$���4N�բC���p%�q\ؖ ,6l�����Exs�\L�d�%8��R��O������@�$u��%�+3��y@��m����@���H�0D��cщG�9����˦W�U���q��Z���y:�\8,�ɴ`�:zά���TZʟ�^m�;�f<D�$�i��@�������?.H��D�Χ�z��Xgg��$uSN.����c�CMmw�PM�|�s�ɞ,��pfeA��Y�����a ����񨙽���������ȋ�xJhE7;�~l�?��VBl{�g2
�j�U[��TN�f����bk��;i���$d�%�6T^x��P�k0{h|�\�U�Zf_���"-UǕ��uJ�^�m����S����..�<i
J���������<�Hݓ��S[[[m�o�V#�v!��xD�Gw2j���KM�r��b&c�w��cV������Gq��n�
��3~��fZ6�93���X3��o��n�7�6�'�!C���.)��J�}�f��=x��^�y=�d��ⵆ�a�P+�
���Q
.O�	Xdj�L޸��!~�r�� ��Af?����NO[�����7Y�+e��i4Lt����Dc\]�Yd	@�� ��%$ӂy1�����K��0��=�����h�
E<�ze+�fA�}���4�[b��]�@Jf�a��_S+y�Y��3��T��X`W-TO��I����Sg4�n)8|�*��Z�7r8�=� 1�S4�@�Y�J�Sr�k��;��nη6���|s�W��=�=�#��,��J�>��y�*w'z���cx=�w�1,RFI�%��4�X������kO>�M�c��*��9���*���9/�TN��<����9�����i��T�;Q[!��ޗ�z���Q�P� ?,�=|��D�Gw�E������H��N����sv;�,p��T՟ܾ���ǆ��ǔ�A��K�G�:�p�?��.�W�~���]{[д��l�F�J@PP0���h�qq�Y��9�ޟ}��4�y*l��#d0��b�boہ F08�cy��t&����-3���'��/���j�:<�L��739�����3��9/�/̛~�E-`���__���e���:h�2c
��x/�I͞ب\)Ϣ�Y|�C���dT	U��}[�0�ɮ��w�H��%Q�=F�[b�)��V��.$2�3wp�~k����&8⑩���T�~�`��I�F>��ێF `���8w9���,{��{�q�gVEB�~Oή�{�[���C��Uif���VF�� u����e�iN�p4emr4;���(fBi�J v�b�TO�_��3�6��&Q3��xD���j�듊Vqq���{�
��6hP���wG���+ƗaM.��a���%c��?�V}H��6��Z�����]���m6�nK��n��/�mC&���T�e���W)(�Qg��WȎtH�	/p���>�Ϫ\�����*�.d?)���'��&fG��g��]C�P�M�UD��	�.���00�;&}R��SO|�]���Y�?�X��(�$3\��\�����n��ڭnǪ���ҳ���ȕ�䵌8Iˇ�!Ku��1�gݯ��k��B�
 �ޭA�I�g���e ��];E�E]Ӥ"�dP�Z���w�nZ�m ���0��_O�b�t;\�	�%���ȍ��~�n�o�����������1��ܽ�y���sZV��[��ß���'�U������7x�uԬ�Ag�b;��\'��M�o� �G�B���f?Rϋ��S["xR���ah��/�a�dNS]Խ_������q'q��a�#�0��A��P����ML�?vw	�.I��K2�{p����W��R�vޓ�$�u�CǯOZ�D�L�x�NƆkh�X,J�T4��6[�>	��#ް���h�;���z��&� N��`���J�]�U��v���+�O+�V@�>>�v�����q�B�!�/�Ӄ,���zȡ�t�n��A]E��@�L��H�!�=)�N�ڙ�3 ���N�r��S������s�L�Jz��� *Ћ���n}�|�_ф偺��|w�U�Zjl���s����/�x���WK�q�R����5���ߟ*��|рo�Cn�L��}+�o�s�,��c�ᣬ�K������n�ԠeS��X� `�Y�Ű��c��v֡e��J����t�m��Z����v���iF�D��@.�N�>��x����^A8t����o��DH�M�r��
��$d�h��z�mھ5�\��ABVD>R�d���y׎�=(4�����xw�;6�{.�������
�LjF���(��( �Q�^�a��k�:��-�U����������M��b���>�ݺ�?��J<Q��-6[ٗ��!����A��#$��E|Vܘ��{�Z�1�;�x�m���@�nwo"�ܛ/�pp�oD�����4n�|�hd�.0����KdP���>y�˿8K�m�c�ݼ
[����/&��D�j	�*Q	�ZG����j��H/�(��?��L3�!"KXGq��(��Odبqr)����&o�F��I�������$�!�OST�I�T�c�
�L����+M��|������i�K�6�,H#���M�r`��^a:wOF9 5�r�>v���t���η;V�cqS/"�i�p�M�, $l�!�ّ��.�8�.vYk�¥�w��\d��.�����bb�v�`����i�Kh�q�/��������<�$�?E�o��;����k%�)y�����ۤP,�InaG�@���V���mS�S��= �Y;��#!U�j�m����.y- �C��l�Bœ��p*+:�Gs���gg&8���=swr[hƌ g��xcCR|6����	�
]z�ݘ�k�^�W�Pc���[*
���XJ��GM W��r��G�,�!F<�Lo�-�+��U��i6�����o1�z/-umUDɩ��ߔ�5������8dc��C�"�j�S����aL
��*]c� �	�OY�o��U�5�)⸛�WBY��!+Ο,�b����	��ˁ���$�^���uk�l5��J��"W
}!�	
F}vG�fj�;��x��kRc�5}Pz���I[� 5,ɔҥП��n���ݺ�_��n�vq��xVʎ�����|x$�1�z��%������ 4�{]�ݡ�>��Gp;[;��������Y�4&f�����J`.�H&���:D���4 ����}���|�m�Xe^�BsuZZ���b�	����\�υ|��|=�Ks]V�"��3�q��/?�3�RkS�+��������ewSt򧛆g�gG">ΐBAU�Ë3�p���������8�uOw��	���H�#�5(���Sr<����W��~��	���k�k����H��㽥W~)�#Ә�Es樵m�9sn3qQ�=�w�w���$:-��	���;~
D�6��_j@'� �[yK�(X���E%�@BN��\j2m�NYO��,�hQ�)Ry����_��|����T�vB���Bi�KpĈ>��5s��볔��L����^ ��0���7��BeBP۷��/K����&���"B�8b8A#&_��������/�P+��_bp�E%�t�v�{f=�F�Z���{?�4�\��u��6kts>Lt�ӱ��MO�_;bt�ڷy|ȠIe-���>0?�N��!_a��!�]��bBŶ��g1�F֭�Q70�gB�K�vO�����?�m��m���ĩ9�N�Ę.� 3�'e�H�|����_E!�yH����ej+�� 6�&��l��!#*��(u�]o��ۍ�NC]q�
�Z63s���h#�i]� ���iň�7s5~��a�-H7����.V�F�#���PB���Q߻����U#�3Y�
��	"����^�/Yҭ���!�U@l�t |�O ��� �>���]���E�h��r#��}{������+Z��ݮ}��3oN��B������V�N�WK}���Dvh�����#�KKa��9P%�[��zDl2&���a*�g��ֈ�#@H��]�����af"6�#��_Nq�d$�3���uO'<�Czj�9���Qx*�z��q�3NA���U'U��B�}\�r�7�keϰ�E�.��qچhۡ�>�K����Y�] [V�^H�n@?�s$��7m֤~��e�ť������U�ƿ�3�}�+�շ,_OV���v���s��0֗Ep�n��DBPL�l܉��!&�sKx�%�E��D�\��f��&�V�ܵ�;&�q�Qe����w<>�e{aHwWao���H��((K�~�&?w�t�^�E�`�)��<��hџ�q7�,8��q�sj��Q���-4xg@��t�b�ǰ����V����2 �P^e7�T��.�1�G"��s�
�a�L�l���%��g��-
i��B;���o�,��� �S���͙�!�n�ꄩ`2$����{�.���4�ix�~����{��v"@Y}/�����1�K�#Z����,�,4[<$��|�0xDچ�*�FPbQ�$���ƽ!���!��D
#��t�oZD�W���4������1�.H,m��s3���_�iF�<�O�j���v��H��/̎&c�>��<��$ˍ,�?Z:	Z�U���`������ 9TuF;���.9�V7��|�z���!��l�V�X�Iqj���odnwL$)*�9:j�E?��=00^4���R�yB�{��	#�n�fla��?'��z�@�t���ե? Ue,up��O`�n,#;��?z���2�]�?k��3���nR�	�v��z�ێ�����qQ�>|?������"p�>�X��4�-���J;��_�N�	3�U�
}O5��>|�F�|�g��q�	Bt����}�w�߰�Ņ�T	(�@%C+�Y�	O�> ��V�9��mEŹ)�kwfr�H�s����T�Q::gӑ��l���ێ�\{�{�i�B�FL�%��5G��"ou��»���VW���ѕ���~L�|���4���÷<4���g��o�17��v�Wn�f
��Z�R����ȏKAB`�3'��Z�n,g��bw����Dk��F�o(�ޮX+Ȕ�$v�W�e+5�g}
Ӻ@�[_�4�Z��ւ??�;���/7�v<�񶾴""L暷sN���O<�x�6P��<:z�"���9�
1���J���� pJ��B�G��o�f
ŕN��8z)�+k��]�b��8�`R������>��֊�(#�
V^�? �_���8ʣ�@u�����D�$V3�~��o�w�{��R���4���g��-��2�ψ�>�>*�� B!y5��P�������^`�N� A�W�Ԗ�����^�4�'��U"J'�Q_V(�����l��^��i�U�^�m�7�ۜ��'o{{|U3���N��Uuq�+�j�~<����;��&�Df:�͊쐐��o�U70[��b����#� 4cu\M"t(r��:(^��{&!�fPj�5IK���^;��#�{��a�"(�&��]&=�������ak,r|jg�U��f��.]{��mr2��uA�W�T���kS���|9	�r�#�*���%3Oɕ#��$�z�z�1?*��4�*w��o��^�eO��C�-���?f�ܟ�P!ON�E�t)��cynt�@�"7��m֞JU�F��Cޅ�����O�wG���t�������l�U��	�A�% 8*�Pi=�"�2
�NJ.1�	�j)��f�y]�|�L��6����B�l�tfl`C�w.�]��`��YO�����4���b	聲~��)�X��H(��)���KX]_�H �(�B������=���zd�����ۜ#�K�M{T�~���C��OF�߂ڿ��֒T��-�����$���;f.�!
�QC��� IٙHĲ��n}��~�f��ql��&ڞs��2n�{����|j4�dŬ��(=��u��U�)�31������ҰV,�9 I"� -�l_(�/����֪��nrX�ǳb?�t�*�D���'2#�CI��q��#Y�n�L�f�ǔ٢��iϢ����[�܃٠��{���,]��N��������9�ڪZO��tD��IH�O�j�Wx(3��������^�܀]
��C�!x<��s��ȯ���f��^п�"F�q
���^���nYpr]�����h�"1���0��&���F�u#�K8�����!H�<c�,�V�kIv��13���eZ��!6��5�9�|��wL8o�P���3g��_Gރ�ޏ����%�
�+��K���D�j��S]/�o+�'��0ȟ���?�z�ߕ!���{����/���xˋ��;1��`�2�J�2tQ+�X��&Jf��	j���NN�F��f�6�[:�,�"JX,O��e�[����ХJ=��	����`2[%0�bD5A-@ϖu�É油:d��ޚ�
��49�7/����jo+�=uz%�T�ݎ�d^��K`���柬�UVwOѷ:�ݫ�T���~�;<I4`��HQ��+	=T|��|�4j�ޮ�a3N.lz�{sn(�:u�i��~���Y
�#93�x�T
�F�N��+�!z
�|���uR�ְ����ʘ�K,�ZN��˹H�o/�;Z��+˔�L%�r!4��RZH/�44⎘��5:�z�����ۤ�I��|Zֶ���SK�*I�$TOn%�0˟t ��8@����b&'4�؉k�V1�0�>vŽwS����͝�tt�d�<�w���j�_��!���&x�(�Z.p��3�҅�B�pc� V�;j��# Kd�:��E
<wg�aφ�/q�؅/r�5��蝲��}��)⥷�d);RX{�`ʧ�H"�m4�%��=�S{�@o:�����lo����*��-K�>JS�$w��/�# �����4�R�����L���=�Ӭ��i��٨�fڝ/K��>���I����\[�7t�ν �	�sh%iB����taj9uK��i�%mmo/@�~��� ��HWj�q��L}��d3���-��!"��"���m�[?�tKp�Cz�{1W�vQ%��P��'X�&�S[1���4%����O2��>
�6(��I�1gt����U��Č0�1�Qc k�*��aE3���5r���p��f�1�_Z��l�@ϧYÓ��'�P�įĬz���p�������_a�*�jza^&��18\��91�&�����kk���0��n��k��	7u���y�n�MШRI���h��@x��X�(��h#M�6YD㇏���	��;����kstl6&GL��{���"Pgp����p�K�����ô;)�U�<�e���A8K#����p�&J���
|��磷#	��-������h\R'yHl�l�����QR���"��]�Kw��SY��&�Nq����Dg�U����t:�;��S�`�q5k� �`�^��q�z_x�K�O<�ʩ+'	�Z?�k6및�`7K��֑�,M=.�O�,(���Q��z��_o���/�)e���AŢY�܁�cX���G-1T"��sq��C@��������a�Z�#u�&�v!�)�'C��t��6�.ߗhC������
ʴ����� ����&ِ�T�|�ٛEҽ-��� ]����w����J-�^?1�x}�^�:�7�	e~L����Q�1�!�D�x����˄d�ʯ�w�h��|L�����ͣ�H��j�)8v�`C�$^[��V
{�ʿ	I�{:\ڇ�yM�]��&�T�X�JH�K���Pa��(��]�o>s2�+t����;�n��z���PvD�������({�������\��6X��_��g���lĵ,J�f'UG�/'�LP�c���K�z1:�ø��V�E��߀'Ơ>5e�/v]s��'z��G��:1���K!n�4���C�SҶ;�,��h��N}?r����?��މ+jQ��1o���a4֎_��N����#C�u���/r�L�T^�4��}�4�@ �������*Q"��wsM�)K_C�e��5
K6��&T ?�Q)�/��c�R���u���$T���f]w�v(�l�������y\7\is����hۘ����v�8��2���+�gP%�2���1 �!m�ja�➩�Xơ�U�Ѫ^wvl~XҮ�k�-��{�����Z���q��9	q��l�'Z�zt(
Ob��s#�$��452��o;�i��4<TjB�M��~�즱�W`L�o��~�6�C�����=��j�O����ԓYВ�D�'���inz��y��9!����h\*�F��M?��t짽+5�&`o`=��!�;η�3R02Q��,�jH%&؍+���0�@�@+�`Z�c�uѭ����R���$1�����p@--B�Y#���EX���Vt!��U�W��\��(?���6�6��Kq�N�o�Z�撧�#0<��?����q���w�ړ$�Z7���� �%��+C���,��醾_�K�<#B=la=�J�&}x��=��`��,����J�V���r\����˛��TJ��M.��U�Z����օ����3ʚ�(�����/�Z�Υʰ�4�c�8*P������C�VՀN�o,�/	r�Y]�l+޽ns�h��-s~�܁|J���*�z�8� �߅`"�x�1bA�����V�ϋD����iGmI���.���
~�4��ނR��N���v�[����D�@�K����m��c'I"�����4FT���׭b���T�s�d�P���e v��dȈ�/F
����^xOƨ�3�

&/�A��>��Ŏ=���� ��{�{�5|]���Z���OW<��I$����ق�4�]XL	���d�};wD�'.8�������.��$-_.����E	I�������X��#�dوOrp���gÑ�|%l*8i��j{��	A�����Mӱ:�!L�U�^6�.��ց��8�f��8w�d��{�ĕsB�x��W�g�?PY��Og��>��.C��k��9;��y�4��!eF��}I�צ#���ID[���	8���y����Q}�k4j����l��[=u`P|_���1<B>����(�;�tE��yRB��\J����ԥ��,����H�#�����N�Z=�xF��|#��P��s��C�m5EҰ*���8ǩ����l��q?Oh��l��Mb+]Z&Cz�Mzd��Ii�5���}����ԝ\/�O�K8�=�|��d}�r�Jp����44��5�Sl��n�@�����MT2~�)��d���G_���^+cJQ;m�������g%07�6^�b굪>����뤎��z�re%ن�%��:ZՍ�o�2�ʺ$PYy��B��7��̗��ϲ�|
�T����A����~��lɦ�˩,�C9��}��IV��vmf����{\E�Yv�IP�'=]q�I����Kp��v�g�,�~{��i\Ȱ)���f�8���$]̃�}Y�~E��S�+�%.9j�r��W�>6̠�=�Yj������4	\*Qo"�&!U& mv���cO�A~9�KnC.��4F�)�k00d`��SjA��g��W�´e�tO
�G�nY�R��p����E.�����d>�}���%?����' m��s��sͧ~#(�/�h͒�S��V\6t&T|�sX�#� �3,�}",�Ⱥ�_w���kItM���/���Y�=O��Aߖ�N��F��N��xd ��٤����w�����ct���)��͍I
/8��EU;�	v�gǽ�k����Z����w�_g�%�G��� ��7�:���t����ַ����(�Iک����(aH�E��HG4ڻR+5�o� 	t���"���_OL�S,Q.��|�.)Ȕԩ�G6=�݆��X畝�h�7���CX�}�iP�<�J=��.5;��ևF��TyR�&X����F�LRA5,�9���X�*��O�xiysA��۷�s�B�E���"�� �\�s7box&���]'T*@��</;��`��}�w�aN䵵e���+ږ!I+s�е+�|(P�1�a��������^�Z�X�nD��x�����F��CD�m��#�0Z�]�"��)�W]��^�xG�l`9�~Ь���3 ��w��?8vс�,��2��L[�u,���a�4���]h�����}�Q�#oX�N�N�9���ܤ�ݘ���?f渓\��*���dO�i�X��D{�?hlsEQ�և�5̥"ʴ|m�k#ɕ�QS��g��U">�n7���B*r>��ʽ$
�����>�"{भ"��d0q2)/�&Z�
쒯aJ_3 �kŸ����#�ٙy�j�Mmk��?��Xz�F�.&�˭ˣ��a���~��<�qF�T�hK���<]q8�vw�{B�q����jK�:�e�H�[�>�/t���ݗ'��ӧ��ｕ��h�(�p��'��|#G4�l�o:n,7ۺmX��ݹ�HF��1��{�=Yf)v�� �g#rJ�t5K�\#X����������S�}A[��Z�K,{]�����<���=h�0w�OwЀg8�OہFb�z�7Dz?���φ�Dk��Rvw��9)�I�Q����c2~��|��qE~��z�0�l�J8�f2~�>/>��":�}n9�>����x�}�S���`Y�������R~1��7xѾA�%i�lK���>e��C�B�!�^�q�ȫ4ɾ���K2��ϣH�g���������љީ�[1�(�V�U 38�$ׇ�D��(7U?�� _@��n���0 ����e��5�7��� Ԑ����F��
���<����N�L��* �e<�ê�QlF�%꺜�B�8hV�����]˱�����1�.�Ȃ��]�P"m�����x��%NΙ��"�B(	N�P�h'Lל2�&ZI�#��E0�A�?�6��w�c�x&N��g;�٨L�HahvF
WM���'d}V���mCK�9��Y�w�uc�=:��J��}ֆ�E�}�;�ȋݡ�@�o}g��5� }�۴9�Ӭ)��}���)-��~��>��Nɯ௝>���>��-ڡ�]l3�EO�Y��V�3�`8��0d�zz5��tR���9�>l��
Q�����r���Z��9�= *2ƖdH���H=�B�k�������1�C.��&��>_Rգ�z&�[% �{�IXKw^	����'�U�T��/umu��P�k��]K	����,����?e둅�~8���R�k)�p Fx��C�t�2Yv�-o�}�ו��vZ�� _rCc�X��wh���c��ċЗ�S�Ae��X���%�X_��y�k�ͫ�+c��Bc}�����^g�����JNU�E�a� ��%:AG!9>��_��:��Y��u@3/��`�\�PЁ@�:~B3C���i���1�O
�y:#k��a�sVHq<�7�"��ٮ{9>�����>���	͚��W$�<��U��܃w'7r !��o�PX)ǌ��9��LN�0�>|kj?>�3	�~��Y>a;@;����e���!��N�sL׎���un�������_���\��\��uad�kjKȂj�
�~��Go*�	@f�o0�i��2?\ ��B>kIco�]Jڡg��_��n�뿽[�����7���n��^�=_���֮}IZ,mO�!a���ae'9��<@�� �A0*�g�/�h�3�x�?���"��f�Z���Զ}6l ��3ʼ�S D�ʅ03W *��� 4�����ʞH�K�xfI�RttQ�����
H��8��y���s���Og�D��y(��:�[�o�P�a�s������s��?]d�q~Y���S$N8��4�F�v�=��2�ʕt��	�Z`H_�5O��9��\���t�D�FQ��P'$��p��Q�|L:`���yM�I���!���OL1�Q%~cK���/&<�W�ک0���ڗ&bj�gc��:+hᰳr�_�yj6�$*Z�8t���`��
}1��)pV����O	�Y�@��;w�W��9�>��k�Hwh�&L)��ʦTL0A1�\{����� JršC��~A�{���nG3R��Hgw���n)����pj��$�n,h�f�''�s�J2�LT�"�e���H�D��x;�R�?"䓙c+�RQ�}�x{	T��={Z��NWY{�{�[�᥋��N�f����v�^� �S�Ӭ�!�}ү������
7H��G���������n�XU�>`3nU��ҿ��U�����&�b�@�Xh���Ʉ�8���9ڑgG���S���#�i��_����R\�I�s��Ŭ^ ��)�rsdmS]o�l'��������~!<�w\#���}�O�����3X�<�`r��v��b����f�c�v���&ʅ2]+Y���=[�Y���Z7�Xۆ̎&;���_'���X�X���䁬ȥ����CЌ�Z�]�����ȱ�kA�����V�.@\�ɞ<e����Xa&H�>'UT�g,�r6c
�+�C�e�������}4k�3e�����~�'�b�� SE�Hd�h�ʫ��5m�����l�[�(�1��!F&)�C�h�S!���[ۚ�q:��c7����I�xuz;q�z2�`��+����w����U1Z�fc�.��䖲��f`�a�؇xq+;���(��uu �f�6NkܤS��YE<�z�:��d8>;6�3�<�T~!6�@րhF���"C��d�-�e��q�t@�ܨ�e�l��t����?,�AI�"�"��p&,�R�?�����������@(|�ٻ��ؠs��v'
����.�cCyE6���y�_�ږ�L�b�|3���H'¨���w=`��(V��5N0�`qx�*}�8�6�^�Pw���a�?& ��]Rc�>`N#��A�Չ3��7�׼ ���3�Ǆ
�jm ��b�YBZ��ń���V�����@"k���5qg$�4 c�
7����NA�Ih
������(Ь1�~b���e��9��S������nO� ���;L͑W��MV����Z�5Az1^��΀-�5�?pg�MAg�Z��3��q�fbQ�i�
�	�T�j�0� ���*���9�/�� �x�?��Y�1�����w	��	�h�󱏃��G��� ^W̑~pMԬ���<Ui�cMG驄3��@����9k,�iG`�%B]BEn�Q3v$uA�p���X�]Q���
�d�3��W�G5pU:m����KM���,s���jO��4�ω*k���{�[\�Б�X8~�Y��=�j��M���fc�̶%VM ��]�2��+�!����Jw燿�|�WܮA�Y�Rݧ�K��|k7R��$�m"S�L�r���p�>>� �=���f��`s
�`��׫g�r�fX��k�O�L�-w��Z�� ��q���6)ӥ3�I�R�ƅ<�^�G���P]W�c]��a�<����\7�� q�$Pf;�#���X��紋 ��T�(� ^أnZ�d�>�=�o�N��X��$pn�$e�ES=z�&��#�)j�M�p���j1f<w�BwWi��cL ���1�&]�R��C����'�d�P�
�}^�].���U`QGQ��:Sh �L]��GGǗ��ѐv�)�>�U�j�A���� ���y�FcD���?B��PMw4����Ƭ�"���5Z���#��N�Y/!��Ҏ9��w��w('l�I��jPif�F��m�>�q�$~�.���\l0]K	�%�\~�l��;���i��ؖ����=ԛ��������§�a�Ijw�
�#_P8���l���Z��p���\ -����Y���$՝_�e�ahڪ�Mr�:��#o�fۗt>�G�e8��A��, A8�n�P����>dv|ZvMB��PY�����׺�?��ľ��eci��K���Bz��@Z3����FZ�-���u �
��t���Z=��l�_:}�S6.O�Br.?��}�Fp�򬹯�'LL��;�%��ш�RZ`)�S�H�j�4�'}NZ��1ш�؏��I�ɵl��Ih�؏�n_'_�� �@!I�mWM-G�I/�G�s@#,���T^k��=�b�p�<�~��)3I<��ח�n9�<Yiw:�;qc0�C�u�wR �B�/ڲ,հW1/(?-F�=Ux�}���M�7����Xt$���.��!��M���}���m	�O�=���ۻ�T�\�"��3��:6�\Vv�'tG�k��<���.zR@;�z||�n����X����s�_љ���N��j@/���:���b~��0�af3�4��3֭�r ?��jt�c��b��)��J>������;I{A��X|��ړ������La1�R��0��<#�{�1K7{%��_���z�<�]	:��B m���0��G�NZ虢b:VBb.�kTt��I��֧��֧�,F{M�
����{�����b#�DU�|ǻ���%�F�px�F��j?E��߶�Y���Ǥk2P�áP��R��槵}	f��H����oꆿ���EU�UuaTW�Ar��tŴ����p��tU�n�ﰮ�X��e �9�dV&��!L�R��#����	H,
�Y��+vp�ӳ�,[ ������3䕠�}�k�FF#W�ƳA��?�a=M0��1(�d7�� ]������sb�S�`���f+I�R9�' S@ϵ���J[��y�k�3U#��3E�>e�Y�֥�0�$k���*uq�"�_Tx��D���:�S*[`C�~S�B���(��5e̩��/,�'���,�^��գs�A=2mW��:kh �]�y�G�G;f?��4�0�T�j��H�,zH���ߥbRQ�Ƞ��D��a1ƪg�yƩ�n~hv�J��|�`b��N���G�0B4�j���'�(7'}ǯ��L�zfg-��\%�>p4�_�6��ᥓ�僙�x��3��V܏+=�鲫�*��*~e��􊐕-'(0Ǖ��e˥�7��{�;���t[b�RXѷf���;��Ko"��bv��;���.�lq���<FBoc��!� �G��P7��Ǆ�tm՞c1��6ԉ~�����Ь~�;�"ِ�*�!�XY�l��K��I6����Ǖ��W)L���ٗ�8�D��CfT�B;c#����:�P$����u_��C���8�\��gQq�8�y�t����ߏ�j��fZ�l�#*F������d'p���y==3	�l����=���~	�9ą}��ӓ�� x
s��fI�&�,ƶ���`�1�9�nG��l���9M~(�)�b����m�8�4|�X�
ny_���>�B��a������E5o�t��l����:;o:;����(r��M`� /����Π�߼/mP1B��*^V1�.�4������Gl%XD;DH�W���H3�	�g7pdp\���ɢ"�E)&��+�ƺ�}��$'��S}��M�;x���]e%��G�RdFO
O�<9��Wߧ ��`.� �iM8�L���L�,FKY��b��wU�.G��8A +g"�eM,��C��-?�qEOt�tvS㑀��w~�R�ewN�+�R�lh�2�;^U�.���<e�d�(FIX�m�P�h}�����O�h7|�K�rt3�/k�#������w"͆������P0���Pg����bo�2ا����!SrUey
�m�U�k���`�{(Y*�c�P����$�A�@�(��W����k�����5FO���^����0�VT����XZ"{ՙi�����܃mR��]�o2Tq�f�qPq�m� ��/iW0>��[���A�e�3�8�}�n8n����8���@�k/��G<� �(�,O���w�Æ ���*�v��u�]���L�6d��>$h<��Ӏ�s���ޜ4tf.�+<Qu�``�/���Yve�1�T F��̲X�}����Ɲ���(g���y3��x!���+��:���݀r1<v
(+eG�[YQ�b~��&�������T9<浣��E�lS��Rv�3R�b�F���=IPe �E9;c���̞
-S��`�0�<��PTjZ�����`F���젻�s��[���4:?i�\��7u�W�jya\��j�����c���])Gn}J(�`��w/�L!������$��UڐK����է,���V�����]�[���;
͡5��S2�#lԇ��(=�)��g��>�I��d�{�	�5:��G�K��)94z[+��<��pCD8(D��	�/F����z�e����l�d����,�����/z8���n3�s
:�S��~�ιmLSBa�8�,@�	DunǑ�&�N	�eML�����t��I�GO�������c��+���b��� M������T�.��|���՞	��^�R��k�i�`{�5L�`�y>x�af��BOEy��q����d�q��VU���Vl(�ɛ�ԥ���u�,�@�Y�گ�\o޸�0������U���R�ড়3,~�������U茞>lgM��j{����=~ +�tJ���BFZ9Ϙ���r�KP�����2��Y�M�l��P��_R���\	������GSI��t��	m�h2��'h��t��b�Ʒ�Cl��PR�x�q����{v���߳���iX�J(��B�I�3~����M7� |K�6=>PK��nGl��RM)��E��h4������tz|a�e�脧C�@bu!_C�C��ĩ��T���'�+T�Z!9���w/w�o��n�����u.	.�Z���ܿ=(�s�A�pia,셽�h�S�Mo���1Yك-C�ҷ�E��0�/��?ж~#��d��"��}��y�ڠd�`]����	#�<l�eA{�T���G-#���ZO��� K@����<�����8N���6Q���T؆�����[D+���R�D�<�`{i�j^���5�<
 m�Ѧ?��p'� 7?�=ȩ0�j��
wzX��P��`\��f��%➭p=!�
�39�Z2F1Q�%�X��X���3p�_�S�`���ꩧ��c� �s
5��Ԭ���W!�g6WT5 �B^Bc��2���i�N�y&�����o�3{�ɎhةAr[����x�����ZZ��L-�՜�KK�쁦�O���tή�@29kf�	���8���YD�Tع�Y��d~x���D�"qdU�U�E�9��3�:�r
�;��u$loZ�"�����7MLЦ6w���f��s���@�}~����=��zU���'�@n�6#�b�:��#2��0� �T{nH�9�/g8	���?���8r�҉���k�
_�����-����1��`� X�3��/���8�]���c�5O���+�0��Yde��p�3͡���s1V�q����v�z[��cuM�,�;��G��*K����D��@ϔ�\ A2;p*r�60 6�ܓ��P���V�.�du-�����B���&&���+��'�M�����xBU<s�״���sg=��t��yeN<I�~�	.}a���wb`��N���!{� ��)�g�&�肪��*�C�����3`����E~5N���`�z�AOJt�a�ŀR�3�Q_�C�Q��Y��*�Ј�(����|д����)�\���N3}�J�	�� %Үjzq��G��C�g�!m(�����3�C�i��1���NN�)�/9�>����>��t�DC*ɐ���c�u �_G̲�������O���8�r�:��j𸛷���ɖ�b�����hw���E��p��[\���[�]�r}����08䒡�މs���u)�Lҵ��8�l/Ba���E}1l�ן�wn���jF��ԄR8m�����}�u$�8eښ>ܒ@���Z�����]\��+��g���g:� ��P
�_�*��á��'��	P��\�������Y%zH�2}=�5��!�=��ͳ_3�:VݧFr3��+؞ ��tq:��A��5�>4��3��:EBf�C�����t���Ds�xnN Y����h�gu�k�E�n��̣+�~vw�֒�����U����� ;�U���gBVZE�.��g�p�!�n&`�M
��6��Θ:c�垮�=�0=%p&���44��HY1;������2EO{ ��l���SQ�a�7)��S%h]��Ϻ��igBcj��iJ��
�Z����䌾v�\w�@�`���Pv҉��H1�B�#�qq��!B��BNҿ+���p�ꨐV��!:c����u0=�[/����0������$�᳡<Z ����	;�l�,�Ɇ��*K�y�Z=���R�X�v����P�pw�v��ou��\ǡ�R��.w������{ji1��&��m��t( @��!$��	�{_� 024U^����FQ?i�Z/����~��n��/u�¡wt��)m�{��+o�N��A=��N/a� }�Q�%�p#hQj��z�C�[�m��5��p��a���'��.�g(Ă�������;<e��p�3Y�b����c��$�tS��b�f^X)��l�*��9 �\�w/�;�X�<�L���R�m���d>��!��}�p3tK~`���¶c�P�ZAN��T8WlM���"���Ȫ׃��	�ݺ�P�ْ��P'���/����n�J��T���\��
��f]':�M��y�P$���u�����U�p.w��7�1�%��P�#i�t���N�W�%#CT�MZ�h[�l�:[��e��f[��*��D���[d�bu�U�F��Q��UCfm0GU/��Th@Ru�g�
S�^�:�T~�0����3��Æ~Lz���U�Zl�UuM�K{d�$�ɡ��gh��'�pb.��`@�yJ�Wv2M�
'��#��ʻV�;�H
r��x8!�Tde9\��,F:{33y�8�`�R1#��.������7��O�u��RE��h��n|^t/)����X��������c
Q�HQ-��D�Vi�@�	c� ?�h�e@<���h!���9 ���\#:�?�l�.[SM�����~�n�����%m���B6mj`��CR AY��r�ކ�0���l�2�K����%ȟ� J�R:*�¦8~�D�C�$ ~���H�%��Y$X#��"��ږ�:�d
]�'��sb[	�h�,�]�*�b{ݷ 3��H�ɩ�J���W0����zUb�k]��в@��k��7��d�*�森01�
������,7��.ա�*���|�Z��8e,�V���1J��QwHal�9��G_�
�W2Ǳk��ވW�B<莎��^z��_�h ���_�3T��25j0��aEI3� n��G2����qyw�7S"���[��:.x�)_Q�0IsW�e"Ϭ�yI�q�m��1�~�Dm��4�;b�w��*�@y|4�64cšL*k�krƼ֨[Ì5��,m[�d�T�1��*ra�0>����+�=0��pX�b[ןI�杤C��ܼ2��zQu,��|����
���vȪμ3W���L���G|^���nx�!u�|s�����{a�p��t�5��0��N��1�3�]�(�a��h|k@��+�*�C�+���k�k?=�X�*�r~e���1�5�I����|����')��/��;�_�Lٶ��C5a�^ST�_�L�e[N���6��k1�0C����Sv�� \j��w�X��
�`�A15|�zb�d�������s�$���x�R�o�L-!m�����Hf�3kx�jt���5�33���|0�'�d!
wH3Ͼ,@��ަ�
���m��W�/�1��tAU^㈂�0��3��CF� N��;���9�^�t(�������6ce�8+o:+W����M��.Lv}f%"+��?
cm ��lEW����A�fu�E͊-*�Q1NN��)����>C5x�7% b���=���Q�yE hC��q
�l9~�0Z����ZqLGkB��vP?�и�] �I�	���}<+�4�U�i��U��D�Je�J���દ
�3K�L���69�͋p�`��3]3�F�@���֑8��[ݽ��`���畺��l
[+�6|�ۺ�����>�����B�3�;"Vf�ιR+�Z���5��o;vل�
0D�	M.]��;������C9|�x�r�nn6����`�l�^`V�ҪJ�A#S)�.��>Y��,_j��"#ZV��u���`&���ʬ��{��O�}sf����וO���z|�X`�����F���Dn]��� <�"aS�ma3�»������6�ƹ�rI	��Q��p��(��"�f� ? �|n��yt�:Z!7���S���ޮt@
e���oP�#�����$1.���'*;�CAժK�{++�W�F�8�u�U��nm/�>��LY���3u�_�ɪ��)�U��ZeV0@�f0�k������jp�L=�? ~��3H�=����5#�E�� -
�Y��l�?P3�p���}B�A.Ɇz@���C���W��H:��؞��&l��I�u��B�:����70v|f�-� �N4@a�(8g&���b��[U�6�Y	���� !h홉r��@\�b D��gg��]����j������v���?���\����-釖ݾD���u���t�?�;b��7�w��&ˤA�	�u��T��@��a�b
Y�o�i��Jl]�<ܭ)�zbp#'��p��^���u���*���?}Ʉ���C~�2x��Ff��陙�{�4Vv�\k48l���!��^�?E�,&�zd�U�7taC�q]�@2Ó��>©\3@��^⳼2��7�y#�@����<@�g� R������ǹ�#�L��Ty���!]BU�.a=��Me���٨�`'�,�3E���)v(���oH�s�܅���n_�?@PTEGȫ�Vv|�f����:n��W��tl�m0��vY���vZ��E�ګ���v�_��~�����*7���A���X�;�>���Jge�h��Ne�%� �vn�Tj�C���:��p��p0���`�cdd�����pQ|Nޙ��w��nli�K���f�Im{ � /绮� �|C�����,�8y �����eN���~�`��!Ddw���)2��w �~ g� B�@��a2�lcу��d1r=���ɺ�+ٟߐ:��b�5�-J��]P!���C����D79PhB�dM�g:��N���n�/�G��[�����;�;J�_8�J?6��Ѓ�Bp�����쐴Dӵ���ƅ���c�R��� ��O��+f'KU�1:(�<�H�HҠ��+������>����U�?r}	���B�W?�dd�*k��� ���`X�
CpO�g�/\ =_k�4����,g_}�|�+4���f&�`��A�a���򰭥+�����6�W�`Ϭ�XX�[�U��D����E��ݢ�e����9q��A�>t�/4P��貘�/ PB�mMx`���,Mƒ��]�=���&�&2��9��?h}.]��2HQ\�WU�.֧�r�R?�U����KJ���Y�@Ag튿��� �V�5��<�HUieV3���D�����`b9>DE} ؙ��C��]�D�9#���0�&/P7�Q� ���91����P�&k
s��p�m��j� �`��%��D�ǚEg��b��ثk�m� gT�6����-��0��>d�Fاc��!,���P�*[agZlX̴˱��LC�S3g3A�3�2��hbv���0V�k�n��v�o�;j/��j�/��޷�������n���2�T�W�[��Y��p���2��񴻏�[U�l��x�|�7v��]�ؐvCm;(�7�>F�gM��d��k�Cwbڏb�X`���'�f�q>��-�˯�1�d���cG:�Lg�g`(��'� a����m� 92�"<����I06�+�n2wQ�ۀ�Ϗ�Y�����}�.*C����<ar2�eM)��V�Ɗ�$������UU8�r�-�wls� ��D�]�1�S��N��d,�v�����W����qا^Tt��
���������ᵯkׯy���&]P/0�{Q,1�g�hU1��
U�D&pZ&i�4p�u&,�@Й�̯�$��` �n�� r���3�	wU��^x���5cc�9�+*�b��輸�Hi��T$���{���"���A$��Lq��q����GR�h $6��p��k��	�,�{^lИ��.�5]��X�,wU�ijT�E'�U�dYHh"U��M�L��� �����I��&5��0@m���)����!��X��W\�>�e��b�mg�Z�L����C!��(@�u���vk=D��P��=郎~��w�O�r�~|׶�mw���gik_������N��ۻ����_���!slA6�B��S���&����G������C��m}�wv[o{�S�J�;p'r���f����E��E���6����`�0���m��Ҝ��{TZ�0?ԁb<]������1�C�"�
��T;��؞�Gl+��`�D
����"4��6�g��hR�ߙA�{X�O,��uN^>æ���lw � <��'�l��Po��<�����+�}� j�Ӭ���g'�{N5x	u�ᬖ#�Laf�63d��Dɜ���8=]�@�466׺�bqx�&��D�,&L��>\��	֘LQ����<��ڋ��.M�R�Q�Z�Cj�}��	���b2_L�n޼�}�M>��_ml��st�7�{.�+=E�ѻ�#��u�=
���{w��`*�E�f�N�=���cd,C��ʕ+P���S��n߹�d5PޣN��Ck���D��1��n(g��@\Ҋ��NM�&�U��R�)�6S�kCNz�A|MN
���Z�� [c�ws阉��3kf�T�(��&�9e]eA٩�<�w�'"l%�������Ph�����2�
������q���^#Y�Z����zV@ۢ^�C*�� �8|�wz�>����_>ӭ�s=��z�@q���@�����ζ�"
7����>ӽ(�j�P�h�����;�����w�O����wGT����S�m�1q�U�-��:,?���l\�3!�����8�E��$��X�^`c%��h5�eQ����C�	v�~it:���91\QXҌ�	A.��(� x��M�
����H��L�a[@V��2���*���I*+�U�r���(��Z"�dogE8o�%�ǫp?��
�/���� w��k1�����i�:R��Ne@�6��|Dգ�Yg�-�v��-1�I�РO0F�b���2"���*�nz�ݥ�yb���K��Ζ���:���檛=G�7�
��ϧ�
�ZC$}� ��S�����H<�8��:h �L\�Wv�|�����J1<ffȞ�hl��@5S�/�$@W��|vO�enG����}�.*$v�����1F��q��@bf��h>���wk�6Ў��rL�>7�L�4^����U6kZ��0��8F=��@WQ� ���`fkg�?f#<��q�>	��"��n��ty>��g��f��tp|��9�+f�f����M`�xqV��$�.� e�&��n ���^��mH����}��}�fw���o}o�����-/�AIe��t���tC�W�x�����uǟ���ەn��QQK���-�Z��)��H�@��8	�
�Mgrx�F�rr��w7?��݆2�\������`�d�|��&uR�$���k�(m���Q�kk�m�nc�.���nB�KZ��-�Q��H���	0�%	��������S��@@����J�rεe�q-]�kI����l���QȽe�Bc7 N��q��&�C���_�vךh�=:���$� �oغu� p����-s�� �]�B!�V1L�zz��z�]�h~�;�}Wߍ
s�a�ϱ��@vMĞ�y��G H�����=�D��zB�/!�-M�s`��}�A�j��Rv�S��x[������}�NM��=fJ��G��R՝ͥ���xb	��e1���q�B�4Pk`�x�]��'E�Y2����>-N�Jx !%QB����������6�g���D���)�s�er�Y�0L}N�� ��r��)�O}N�T��,�v�u��{��%�EQ9�yN'��J�k��<����$�ϡ�U^��&k
��Ā��؟_�w��=�;� �x��
8�1q��QM%9��׻�_�hwC/|��u�oz��9�]���G����@������ kV=���j��C��*ϵ���BJ㡊�!H�hؿ����n���)��
C�a%�ͻU	L�J��t�y��婛?C3�go�����x�	ѢX'�F=�O1�P�I��;I��fP�Q7���)���e\� ����*s��
���\П�����ye?	@���{%��m�k/���-���]�uu���"��z?4�d9����Ys�>���1�����K�����Ԉ�Y�0�D�[��l�k��w���N�9T���doTG�2� <n�#pͺ�Q���6?��s}=��\���-���Īp?�q0f�6���c�RP�����o��^�����؜K̲��0P��0p�zPsG,N�����q(^�H��V��U[�L��}�k���Q��������;7o{0��`}�^�8�R��Y(�xK��"�T�Eő��>6���.Х0Κ4A���~L5;@�.+����Ax��Y���2}3@v09��S��0�B=x�5k ����k�O��H᠅��r�ڣ0�j���ej6]0���7K�N�b��&%��Q�/��ZU�bq� ��r���Nv�����G>�M��b���m+��mn+ܸ��FU�搸�\gdvm�X �b���.〣%)غ7�:�<ߝ|�����c�މª&c�z"�.X�@�����F��]e�	�N�n�aWV�;�N=����(Q��`��	�#�3 .tO�	;Q�k�b�ٹ�RuS`�B���m4������P�.Dȟu�zօ��!Y�"��kZ(�{�������
�e�/�$,;��ܳ��*+aӞ��� �Q�qP�'��8�`����X0�~va��E�=������r�Zo. ����M71���a��c�D-:�U�T;��*�j�����{�,Gu�g\�m�S7��:�����޼�-�@������ q�ъA�A��G�E��\�v�[���T�!�R���q��?�#d�����>޿��f��_��gz,�Jk��zC�#--�,B 婢ڍ9��\���i�:��ӣH������3��c:_i�s�vaFB��ԉ8�:	;1�Ff�x_��9�>|���o㜨H�6
���T:'1Fvl?��H���s�!�ܶ���}�"� Ω���,Img%�NTۣ�]R�/�ݵp�I� ��BD���;�Q��K���ǻ�[�խ]y���T��A'�(�:�tk��n�l0�h�����f��q�;�������F�}��;�e�� � 0Q�3TyN�pQǋ�����a�|qM�ĥ.`	QTH�gг8��X��$��=9��P����n~S��\G'�^��(�0D��7�
���E�d�q���ר��U�]<3����Y��+(^��{&G�V*3�zPN���K�)��d�ԫn�:��F�&q�q���2��"�F]��P[���<�4���[cX�|��sa��3(a���{?3}�ɔ�BU���.�eS�&^;�[i�5��s�u.�T5�
Ÿ%9FhѴ�-7<���^1�u�,�@�Y��/�\5hl;������
{c�ŷ(���VdP�	��r`5#,���v_z�Ie����6#���9���fr˃;��8�ca��X�?�S�F����N�M��s)z'BS4����p׈P�����8F�� !g^:��m^Qd�f�Nf����r
P` ,Ltٶbbs�k&�:�׈Y���*�cTULSfw����1[�~�~�o\i�`�����o���S a<X "�j%�R�����8gg��Z��g���g��Y�GaE	���|�Mݡ�˗�5�ll;��6�w���ԓ���4��ϡ���\-В��A��:�V"�)mӋ�W�벛qF�h�I+������l�62��g���G�<�M�؟�aJ@,���T�U4_<��nv����_Թ(,�gs��k�;-���s��h�ʽB�XA
��&�2����T67#-.,�7�2�O
�ש�b^�@��8�;[��e-x�R���,�Y� j�ɨrB���R������C�����V����ΐ}X��y���� ��7�ҖI�=��g.&�������x��S=)^�+ܒV���{��ǿ�:_�su�gۻ;~�wf���^Z�Y��D�ַ�ڻpʎ���p{�%4t����<W5ܶ&H��?�y������](cWZ/fZ��X���pf��y�.�����)^�6h���޶đ@ �1t=���쏻ì8ͬ-�4F����4��'������Tځ@���R�� E�6R�Y�4l떘����6�Yc�e؞��0�����E�Wa��Tٯ��)�S����e�����+�D��;9ͅf��5R��E]�4�"x���N�.�P��$�h~+!��Q�2�gF
 �0�#�s`���T�̝>�����'ۖ���I-�.�f	lN ��ȁ��������[�$%M����Y ;�#�|���IA&�NQ�z$V�}�503ʨ32���&{�y��;�+=T�u��� U@�����3�Ճ��[��|�6D���+�6 �Q@fj	���:��<ZW���M1�-�ͫʢ������սG��eӻ׻�>�>�%�{���)�s�%�%R�pB�l2�d�!!(��L��}'���r��t��[q�:~:�s�c�ԛ ̿�-(a�"�=Pz`�sB�
v�`��}���C��{���r8��\���qN<;<x�	y<�T�ޝ�)y���g���#=�=�}��>�{ч�f�0�׮ɮy��)M\�<c�OM��h�\F��*�pv�>w9 �_���TaГ����tF~7tF.�+9���t���5DN�P��3�T�1D��� �����>�hU���w���6��z[�DY#з�7#�L�r�� 0�����0;�	;h�ie�I�c����"՟(Bs"���9�L�"���ݭ�`
]3�Q7���S�6�Lܮ$Ĩ��z��\'(��{�$V�0����O��=�v�y�Ś��7v��מפ���pP3f��ĩ8F9oÑr`��2Lћ�p�3s���\RD�;몘EJ���FvR �9�'h�}�V3h͌Ԩ��@�,T�&�m"{��2�ܲ�{38��40�u\�v I��-;Z>�f�}ȒsŁr�ю"����<V��
u� � ����������̓����i�ހI�̍�Y�P��6b���~����G�6z�[�=��;~�w�X1��{��R��@�g��s�ɗ>ߝ�6��5U,?Ԅ`�&FsC�#�4Q�jJ�f��tF�9�Ub��~ed�t�nX��uϬI��I�p��)� F�z@#�#p��-��XχS�]�����<���t�/���Õ�'�`@����NL�Y3���7�5)+��$�5z�SyV�c?�H���}��!��H�,N49�y�p�+M�Җ����m(�5��6�H.�j6�{UzA1��^/@�6(Ȋ�6�O�����,Y����t�_�j`PK�f�3C��.���HF����_R(���3�+���_����ի��O?mviKb�)��0>n�����U���VD6`g�����db�x�40���C5�Y`KA9c�L� �>���N����;�����r��gÑ�N�;N��D�}ČX���4@+[j��X,3�ٳ7��夔�Ƭ\�97ҕ��C�l���5;��%���� �WZMf��uX ��c�,����I`Pm��p�7��#�/R�٥A�	��d��0��p �b�H��p���m�珽��p�j�>��3>�'���[��ȜJMI27>.BJ���eb{/y�]�6�d�]}u{|\��Y����
q��u��7�$�7���6�v���\PLe���-�F{ʶ�}�gAhG�O�U��U~�@
u�
�
 )�st��m��-]��_���:5'�|��ݾ�[
G�B�HkJ-?޿��C��X���%Mto�<�|�-��a��#��R#�80��a~xV�3�E̵O������ZSW����l�"0����N�����1�~ǀu���1ш�-������?j�PA�BH����M�3Q�2r�0n�㞮��c9�&cU��=2	���^��*�����o���������tnH����l��ꮪ�IA3(1� x�L)(o��{��U��;�X�*�O��w�u�|K�!�TD����R,�K9��WB �Yġ1���cp�(�9���c�o���+�;b!3?�����9���b�
�Ł�)'�z�:ԁ�I`
�f(������|Ȁ�>o>��XbW<� �\�С��p��X%���I	��1e&e���)`�zpù��$����X ��M��S�y��z=�u��}Vb�	���%`�|�6��d�U����1K��!�d�p���bkW1��LO��A2F��u�`�����v0���@l7�	�^�ڬ����u�t*�o����!�}�r��ޯ�v���n. �ܐ0|!`;H:�Z��4:m��L&*�'���a� v�15� R��rG�U���q" 9z�j3I�6��x@���ll!�4�i!�\|�{e���n��s�ֆX�[w>>�n���v[7�ܭ�{^6��@KLgQ�jc�3�Y��φR��a� j )%���J��3��Bߕ��Z.B�u}|M<1i #�{�$^�v41:�wӓ�1k0��xyu\!l3�gU��&��1YҤ����w�Ռ[L��e��+W�������^%��Z�LA��+�U<N�NفBg��0 y�Ҭ��l�l98�x4Ȅ^w13���j^H���(��S��N��'}�0�=�=�Cd�[-�,+��`�`��P�Y�)�6�A����C@8�Vl.���
���Z�sԢl7����0[N���X8�#
�����i�>��S�o���@��>c@��,��Bg�n��&�WQ�'i������י9D�>4O2�u&�d'����m��H�Z�����^��z P�&3=�.�-l?��v	}������c��W^�S��(�V�Nn4�`q~yOYh(* T ���.�_���L*�W�Ҋ=�6q��\H�(ǜ��U��f������_��N�m�{t��n��OuSB5{Ը�n�w�>��n�����$�sqOa"�W�OŎkjE�/=��Tb)�۾��M6�w�Y*$�w(*t,���[Z�݁�󖞯,�4v��
��I�z��O(�ktu,}�l��ww���������n�(�*��JT&&��]e��B`ܙ��K��k\]�ie2`ۆ<���:�A5@���{��BiI����7u�Ҍ��9������(t>��N�t�u���M?�Z�q��I�0�"[�������c�[,��/��{�Y{�4tf.��?ѣ��K��#f�MN5hVh@�Zbh�n��j�aᡀ��4]��ZT���Ug��)�-�y��mh���`��vN%O��_#\�pQ���Z��cs�ibi%�mL�k�dA�q���bkϞa�*�
��6}w�&��d�%!%mW�d�T��X��c�ϬN�>Z6�я��R��zAi������c�w�/=��
P�	/�zp��v $v���Qh�Bn=�d��U@�K�*W�6 ��8;6~#����&ұͲ���ūBGO+/��"ӽͤ�=�J�
�����b��KI �,T_��9�b��� ̻��b��1'����* ��(Vi�*C{Q#��Ba� �u�n��
���$�P �e)�o|�f�}�K��}䧺���j
��g���9�YW�+݉�h��X��C+匥���D���;cM)����h#�0���j=2�i�3��
�0��j�_�
++�6�\薻ʬb]�н��ҶUMԜi�$�m�ף�%����s�j��y>]�j�y��雰:k��2��ki�4�D��R�_P���
���Q+�
�3�`\�O�-����*�*0t�|�n�k^�3m���"ݞI[Mx�܌cU��t[L3�%Y����o �'���GA��k���P ��R�̹�2����`�`B63��@�E�s�j% ԀW=zx� �߰F|�X�g��)��E�;���%:ՠfF	��j�t��勤\������?�*"EߎV묉ʧ [i��!�6�@�P�W���U~t0��s�5� ���LH�$�M�4�=��0f:�N�C�c��3v���F�sڳl7�#���%�@ٹ˪�,F輜��+GZ?�l93tD�a);�dJ*���_�b�BX}8,�@�GR�K��9$ȇyN5D��l� ���v��rv[1l�-X���@�]��՚>+,M�ۉ�U�
���h[���a�0�<�S6��Hh�����[=�D	Dޤ�㗹���� ��_s�R��{vS��B<�T��֓!����	�Nu�揼�_}�;�#}�{Mr擽]������8�/\(�=4�=��=ҽ��X�3�G�ϲ�"	8Q�Rǹ�}u��(�n�n�#�J��������Jf�x"z.U2%�C��N�2�qnWa5�4��&{�e��{V9�{����`��(#�g�������d�{����6�	�!�h�� '*}Q͘=L�x��xy�Y�!�6�e���������M$2�g-Oșy5tf.��?��x�y����l��|��fL-����D��@�SČZ���Z@�0Kg���,�BN}C|UEMW�?c���˧��
S ��C�D�m�Y_h�a}�{���'��'��F'��1�%	�&B<��Մ��`��
)�7���i J�V녒qr���E�%9EM%��B7RcY@��1ؒ� #T�>p��8'X^����(����E)0Q�A5mR�M��|'���@J�H�w�e���V�-�[3�����@,���,�\��:v�T��*�SG�
�V?�m�7���=U¹����
piV&�f��Ðv�u�Z�&�
aRÈ�D0#����m}(K����.����䄹�
�����g��=��Zo��^�$���o�>����L�ϊ���^|Z2�K��=��u��������/+�I�G���ǤM��� ��sNWz�E4���،�x�sǤ6��gB������{=�>X�8��f��nVp(8<��1��~�>��́�������=	�.>�V���;w��L�:�
p�JC�dʵ�t]*�0b|��8D"F��u�I@K�5�p�,�i���i�3d�����~����f��k/�/BC��0���0�#�4��Qi����! �f^V5p���M�k&'�r|�Gr ��y�;oJj^l�ԉ4�
u���CT����PQ��a~��z��
�)u8���J	��wJ~��~������D�U���UY�.yd;�)�� A �v�ׂɽ8|F-"&�bƴ�P��L��'7ԙ��ҮR�q'�u� ���jq�A�22S�n����+[�IF$AQ�5b̐qZ�����&�� l�,X��92�bh9�� ʽ߲�_��c]�Z��1��&(<z�7	�|��f�����J	2 �w����V�"��ƥ��T&U_����K�u�����q}���'b�`@H���t�.���?�J �0�r` &C� B��{��S�Y.���4ɸ�������;��?�c����z�$�^SF������ݝ�=���:F�a���聒��+O�9zg_�D�=1H�֏u�#�:�}Yl[�s��8\G�?�AgB
�"(vi=' G}G�K4L^�������gɤ�19��Z��jg��
Ƌ;��m�d�����vǅW�	�J�֗ν
���h��b�	��qz����ih=~�7��Xua��ioπ:���������q`���1X�`�@:��2Д.�u��),�A�u<Ёi����3�Aaf����̊U1����Fb&���3�A�3\����(u|���i<t��j���I�sÁ�̠K�����Ҋgb��n�ĿfŮs�Є��Xi�d/-���p��d!���)d��:#T���A��?t���8k  v��JI'���
p��b�(�M�Eb�O|��z�a���);_���r�U�WN�Th�
=c�\B�aa�D��s�%���9��d��7���X�����J&V'gL�W@����K�	@�a)3g�	�Z�����ZH	Q�XW����N��k���L�z"L�j�-�v=��jbi��j	�����:�$:�	��M��F�v�@pѨ w</d�"QF@!��B�\�&��B���rk���hw��_����d�3�i��}��0��Fe��vx�6'�_m[��X7,����7 �� ��e�4p�2�`��Z���Oh��J����,���9S�ٙb[8�%���,h�|���Pz�c��פ��C[B�
R(�P��&��A˴.��,�qQ?h�ބ����W"�T�]u�`w >|^M����S���[��8[T������W:^��_[h �u��*G��jm���"i��Z�ê�Jh˅�4�0Sc�ZNU�nN�'��=�(��'� b�D�-�V�1�c~�/F�KX��&�=;� ��¹L%c�{!��-U@�L(}!ҵ���GT=�zX��O4������z%4f��0l$T����@�@B��<(�.����q�aD�Ε�k�����Q�{<�ʗ��B"K9��孻b���t�۲��&�ǢmQ�0
�%(�"�yv�Ɉ"��`�52`�c=yVX.&�_�V�d}J��2$z��61.(��;�' ��fm�X,_�,Y)��3�g�?�ĝy�x?,���_�~���D��:�����G�ـN=�̊ � ō�N�)J$Pt2�[\/���|D�H�2�y*�/O���q�AL辷��m��Nt���G��8r��Y���8��
�+8��}��2�O����}Ti��N����s̢qL���e��Ϝ=��6F֜��П��#1��r?���ϸ�Zp���4Ռg���J�(v�¹�O'^��X'�*��bdo�י�@Ag�R����v劊�ݸeP�@�ꬊ��j���te�3-�{�V�]��$18-��0`6�J��L��Yu���,O�J���(��W`���1km>��`�i_�,\1���#YO4]U½�o:t���*]�
��CA b'����]#!����\���v�q�� 8<Z^(����  R�a�4�� \���9��hz���
XM������Mp�ؒ㷃J��ЋjdB�5w]��!0�-�e���*�`T�-�PB�5�X8�ˇ�#�#�iO�[�ii���#\��8�t�ގW%�-���
T�Zrx�1N�3�,���_�ln4�O�~*���<}�x8������] ����
�3�a�S��,oU���̇-Y'�/�����CR�n��b��L����Ac{hw�]��{V���ڧ?#��5���,u\Wq�:������|<���:�o�����X����g�� z�"�����uL�؄�ud32Y�8���/��m���1�}�&d���5��f]��)�v*��|��-~&��l�8�v�/�l6�ih�_ �1U!2�c���x;쏖s�^���_Y�`̦)�fA4=��C�hءS��"�hC�Qe���1 �5q�X��!�6�c=Fz�(���9�
�1pj�,�!����#��!k��]��5Q!�����=E�����qb�!�3�l`D8��0��p�����6�0
~���&�t~
II��9JD:{����K����z뛻��{w�j��ͽn>Vwl�d/i�)���+0 �s�����y8�N�[y�����v�����鄊������O��Q�΀Gt#	�p�0��?�NuW;{12�VhxնY��_y��a�S����}�����Ќ��$h���N�����x���� *�[��s�^[[qP��%�eJ���rh��`	;��%��?�'4k\'���>M��j>>�/	ث�RՑ[`�^g��c�p�l��� �&|F�P�m��9o&
�5d��=�#���9~�=3��N�����~�Dj(�6��X(C��c|����}W�`\;Y�Z��y��}@Qݣ�O,_^G|�ITF�,/��]������9�}�W�4�lT�)Z �?08 ����YJd�b���L0dp0�R<�j� ��/̓7$�F;䙙Cb9D��3��� %B�C�\��Yt���ud���\�lv2���R�k�)�1��Q=g���<�yY�m�z��rf��p�c�B��	��	�9k�H�wf�$��fP�gh���.��c}�nk�= �2���׺�g>��i��X������]JN�|.��~R�!�:��l��V-��[+G\�2�iv�B� ���*��;�DҮ��ۨ�/!JǏH
�F8[��q��+�ʁ:��=�W5@}x(�a���H��äqoT�G�k�� ��?A�����y����;e��E�G��CY3��F^��8����!)�''��}�V.�rބm$�ϗ����Y[ ���ui��q�s�{�[��JE�Ȣ��6��=�ʖ޶��,*W���9[�(�Y�o��k�0;�9�$ �1 T%4�q�� <VU���X��3>U����Pf�J�Y,��.�Ʈ�TTm�3d�F�����rNUNCc��1�)|ȠIFO��`�b�����4�x_ݝ)|�����o�5��i��2���3�>x��a�]��GI�'H�4�ь�u�}g�X��� G�N�}�FcQ�N���왁`��.��P��}$��By�|	�K��~�wV	� � ��p,���xf�E
z���:x��S�v���?c� `#1JK��*tM�Ր�>�e���<�xXǫj��_7�z7|��R���b%�?XCX/� *W��ϋ��3�e�q
>*L��x���:�d��=x̻��Y�����"�a���"�d6X19l������\� F�Ǭ�R��&�И	E��8�г�q�� �O͜%(K 覤f�¦�1̖EH�>�Y���m�^�A03����{��߄g9f�, ��L�E�)b�S�f�~L
����`�Q!����:�}�3�\�2@��N���C�i3��A���yZ(�c��d� �f�N��H�C�CSf ���jv*���JШ����'Y�jĺ�ZL�]��Ǥ�Qm���LY�1Ag�r��OV@g��d0 ̀��� {S�t�	�� K|��� �� ��&�1Q��Y� ";-��'��I��5$�մ�p�!]� �@�Wo,��A��N���ۡ:�}f���K�l;}F�D�B	]�<�U�6|B�d�J�q�� �a��e��E͸�N�����S~f0���`J�R�1"���g�N|�VIl羐n�'��/�Rw�����{��n.�:|ﻻ��ce�) ��	��)���۰ƃ�\Ms��H��l�Ey[0ꙙr�e�X�?fHJ���d#&齟�,���;�
���LD�"Ǚ����eJݏ묄��%H1��<O����(K���O��iE��bߕ�U�W07y�����`#N٦��b�	���O&.�]l��y%���	�^�Taͪ'շfI�Ƚ;c���t4p���{E�b5<�d-�����B���L��Ɍ��%@���9=��J3v�y�{`{����Li�Ar2��W%;`���KT�b�iU����q$��l�~-�@���ھ*gF���[����̠Fg�Siw���0�	\0�ÙR��֍�^퍗���@�� �@�9� G� ���"��9���/�I^s�c��� 4�}N21#�s�;n�	�wkZ�Z4�5��f�ݙ*��3l��<�����q�����ճ0Y ��Ƭ�l�,� G�Q��qx+E�ꊰ���m0�3���Q�X�UZ1�р(�X�-��Y���k �$�S�����>�k�����������nz�rw$�ɹ�!C�:�0�%�vO�XPXO�İJ�jm�;z;�rຮ\��U9�𼹞׉�zV-���O�+/��W��C����Cj�Z�򺑥W����D���o��,���ٖW	$,�F���{lV�@mR|����qN��{Rv�60���Q?���%�`�j�z2�M��%��uʒ����>y��*�O@�&�6�B�ֵ�9G8��n\��"ޝޙ��v��	L�,u���,��!�6g�¤���Y��g�Xۘêaj��XW�D����׌�X�D� $cuW��{b��3�C�#��V8�@�¢S	�7U&��
���Zi=	b�m�{F�m8�����G?�+\��:#h�3r�_�i�x��р�<"/�ijY�����������e�%J����A� [eT��]Q�t���������r�J����5�-�A��N�p���lJR"}3.T���>E�h�!��9�f`�qrha&���	q��{F�hb�d�/��Ӏ��$4h|��"=� �;v�l� ?C�����B���Vv̅��Μ	��KFW��j��VC΁�m�$o�Х2Ǝ�7#m�H�~��]ȥ���{Q�m��8��k��P��W�~�>H笓@T_�P�HB'C�\ׇC��t(�k���+׵��[$r�۷���Y`h�ˬ�9����-���tr�}�*��r4�"Se M��-!2a��$y�د�	�[aF׮Ifɀ��\	�&�!^�����\V��0�b�Y�U��͂�h���\�2o�# EA�l;$��С�v�ǘ$�����x��L�GQK˦�>B�K�И3傍�I��ߠ�g@ό+�3�XӺ
Q�TlUcMwN��n�8���9�I���{��G��t[׉����t91�*��������}a��hbe����������ԗM͚��������^g��	:W����_;.M/� p��� �J��+}�2�|�ë���}���:|O��0I%�v�wNh����h�cv�;\��zix�ϩ.���0�����78��ُ�eV�8��H��8 !�?�r����sy�o�)�'	���y1K�!��ؿ�P���̑'��x�c�_ �&���,#��M�:�;���u�D�[o}W7z��r6ʪ�(C�
U ��(�\���RA�e��$�*-r�P]�2�"C!��	���ſ�3c8�V؆�eC�c�UwuC�_��K?/Qt@��:<j�"�[,S��[�<ڹ� #�1z�i]9GݠfjX�gQ��`�Ȯ�s�.]y%�U�襅���Y�����6G�x9�6�匭<la�Z�k�0� aZ���[眡@/�O	�[krH9_a�`x�w�K?��5$$f�K�mD�M��-����o3S�W`�����e�KW��{��ϗ�w����U1�T�*ˁ�	}�ScZ��6 �R�0]
/�L�X�z��K_����>G���l��LF�m�q���c��^?���L4�ڎ��>�j΀Q������Q�3��Xں23�U��5MYG���ڮ�Ȕ��q�+��X���]x��+���1c�K˻�E�(x_bJ���f�ܱx��e�	90������� �3��p���]$1]O�	�� ̬h�*�Ь��Э92 J�� �&v.�����c�^G`h �c]�^�s�~����#�N>�n�����[���/=��/e��99�`O�]ٹ����0�A����
j�z�JC ��
!��1���Oe:�}�*�l0��;hb�>���wz�f��p9�:�#ט���d �LeУM� r>��>��ˡ_���e �V�� �t��Ľf[�c�<@U����*���Y���n���t@���Ii��uR[�u�n�V �|��ay�X�WG��	���k/z� @�+�.�6U��)Ϡ�|̓9J�,�Ny6�H��������x0�΀&`L�`��>�sW������b���J�/c�JĘ�w�E�ߠ�ɟ>�g�]Ag�*��sԀ�΀s��3&�03#��OՅ 11� rx�� ��Q�>g2�cy�c��!!5/f�0!����l)�!��kv���ۆ@�oh����>#��T�~U����"�d����<3�G5`?1؇n�I�̦�	Z�>�V�Y8�}c�1��t��Dȿ��\�fg�� ?�W�">3��}3�G�E�2@�ު��L��$�ԠQ"�1�vh$������_�?��n�����G�&W��<�-儎�:��b� 	ji` ������^2+ڿj��� �����/���5����}�+�� Հ�� Xr�����;���}/�F�� y���Zŵ�^��-���6�iL��F��}���塶L�����i9&��C����	�P,���\�{�����r^>f_?����ˮ5�г�y:�H�74�r�l�j��Q���GFZ�C�К&�
��8�WsT1������h���lj�b�U�}�g������g�Xe�{�`�x���OM�w��j�Ś����-1I�u��ZAq���WAg�2���Ԭh��C�cPa�� d�H�;p�]�4�iЋu�jV� VB���������2(��Nj}��p���Y��ߡ_#^f��O��T��։4
���N����Nc�)�K�̚�>c84k8����+�S�˱�tAhM�U�C33�f g���Y������n�z?K鉖j��� G�#~�"O����H�s(��R��J_�9m���d�#� ��l���&���+/v[ϼ�u��u9	�����e����IƲ��9YC�P�+ә�Yc�	x  �Z3���KŠ������dg�Ι�~e��u��>$f��뙦�4��7�^�N �`���p-��YH�"�`$F�X;;�M�k)"��0cS̓AH��(� ��I�sO Գ< �}�m\s���zV�{��0�6+�}Rؓ�\��7$��e�[E��k6�H	���x \�y�ك��4Aq�3�(���i����z���sm�L@�a�����{�9�Α11nL��]:R����Xøq��U�CT��=�ѲL�`���?�Ðs/um�� @���d��l��:h �L\��8.z�De\>�v�wERh�S��+{����V�>�/
�fpl��̮a{��������c�q߽w7hp}���f_N�:A����s��L� E�鴄�O4��>$�tq�qt8a��U������Q�S��x('|/o�'�'���`(�>�?^��._�M~�h�%���D0D���Y#f�:����%�QWȚ�D̄��u��#]�'?�->��n�纵��n��+����dKY5��"*T�a����q�2�s�#S*�X�t�=Ӑ�'pCr>�Y�����0 J1�T�5Y�Ȱ/�dN��n���:���ՅK'����� �I�J�9�@;��Ó�O*��ŃJ�B^R����¡�F,�ͭ& Z��q��)��n�n1t��X�a����J�%د��N+�{e�I6'��i�O �;�Tv�4v�XLR�j��+�7 �uI��~d�)�e��C�J��U���*�I���g��n�p�����6���<�'�̓FY��-UZ���)��w �>�r��~vi�!��#˗P:N?l�\�4�5&�廌�ܚ-;�5w�~gX�e�8�ꔭ�1��J+�g��'Č������X�֭[� � |pt���*���~d�q��֍n~��Z�{b+F�*��� ]�b��(���`/p��qEc��CU7 1�㰜�"$q�C	DV�Bf��=u-��j��l�o��*��eqD���*N2g�1y����`&�=�+Ғ������<j�pm�JF]��f��5����Q�pb>�%�ͺUd��c�8�nqC��t�7?�M��P7�>߭��k���n|�z7���n�D�q-��w�5jp�Հ�LC:�
5:�Rvg5T7L؜�N'����<3�z� ,��i�=�CX2lf��2p�N��b`����&}�9�<,�XA�>��@����[�Pv�|������[�Į��a�� "l�Kf��s{�<��㾥,�P,�Pu�LJD�}���e���2�@����)�	d�\F�?�
`���uF��%�^�{ә��2�Y�ٔZv,!��;�l�n_�S��]�~�}^T���O?m�Cf��Hk��/�5�!ƖU��y� ,\s,C�|�r�}�q��� ��E��O�]k��;�f��{k �j���;k���u8����T�	਀-16@Ј�a�aY�CQ�n�3 `A[�L���8q�� �*�_���Bd��t����.1[�w��1і��n_Y�����-�L��L���"��mk���$Mw�6�H��`��=,c
��/q�8%�
;��Q6z���#���R�քV���
+Q��5K-��~ՂY�#hX_����J��T#1�P������������'����7M����D��� 7�c�������b���|K5����BF�&q��@NcŚؠ�¢kf! &����Q]�K�J�}��
T��Z8��%`����by���Y�L�:�}g��Z �P`qcY���
X��9���c���+�i�	���z���ůj6�ú�� 8�.�Goii��-����i��x��� �K��=Q��ZUZ���LJ��9�NCׂu�����឴��q�8D�ZY��Bn*jsN	�����<�6낶O�aRA���V"�X��'���i]BB��ώ�2cO�:�sK�)	 `�g���:=�桘�(�z���I�Dz&lP5�(�Jg��2��=�]�&�6'b�T�I�m�ߘ�!�W8����	=����e~�'��aN�~�2 ����{P�,1�I3��A��T�6�A<���,�֬ͱxһ5���Q͗4�������55m��7�s�g�(��� /W�	�����-	�ȀI�1�I�xM���"��$v�Z�B�d"L�Se-���Й-l��K%�P�������tlrD'>ߺ�����+쉝4LN�`��I�Y��S�������(s����8Q%�������Q,r�sGlN-%�c�d�k%SO����I\���'�.u�w~]7{�����Sr�ʮ�$:]�~D�
]�@�h�}���N5���={`PS@'�2�Ȍ�8�4�mT�T��>�@��
��D�2 �?8S�",`�Tx����@�����2CKF��:�4d�	D��I&ɷ�Y�H�0�l�cdԺŸ�7�6% n '�6�(�(��sؿ8�ոЍE!Lg-���sHR-Q<�1�g7	LZ��&��_�Pѽo������Ha�`� Jq���:���ZBJ�t�/�����R�;2ѳ�3*O��K���a��^*Q�j#R�_�f�Ϩ�0X@NU��L2��5ܬ��'N+��*�P;���I��9V;Bp���?:�x���_�g4�z���¹^$f������j�,`�
j]���� �����Tj]�\��Y*:�zO��D�P���B���Ā~t�����Y�����X�����k�o0bM�>7۔a�Hُ���m��(G�	ke�l�3y3<0	�^+��Y�v���g���2��} �$��t��Bb�Gr=�ώ���;G͠��P�x!�R#!L�����?�A��R,���q���}�6}��kم�#"l3V�}��躞�A9y���ݑ�e��Z���'���ݬ�Yw@�Ű�s�ǌC�DX��s�9��'�CZES���ź2*a��c�T�~2��Ռ��U�+כcI݌{ȱ����^ �[.ÀIF#`�@\���*���.�@��1ܯ��[V� +ɔ�y�"���`0��=�!� c��m�6lM]����5ѱ~���kR7k=�3I +Th��Gx}�`��ӱ���K�����5a[�f�������vl�Z��9:�W���
�5���cC�7�	���LO�4�cS%t�����쭦З�zΤ`:k�����¯���U~�L���<3� ��2���4��APͼ*�`c��9H��ގ�2�����_PEcb��
�������Ͽ�,����H����z6ͬ>��k�."ƃ��A ���n+�} �0sOG�ŢfL�`���[C�g��p��9э�A�H���^�8�>3����g�0��{bO���� )�}��qL^"�C��O�t��o8q�^���Y���M�(��֦
��'+���p� l~�)��沢�$IԺ!��1�J��N֘l�H���C7$�V��fT�1s n[�"�R�S�����1%y_q�aUN�c��Y���pM�s�ֈ�a�
��"�z��$ ވcS��
�y�D�z�{��K����3�a��iT�)l�����U g�w!���G�Be��b��j�Yԏ�zU�+*:C�L5
�Z�{]%.X�Bg�S�V
+�n)�!��B�t
���uW tB��؏������D�h�欢 'Pe��t��C&��[7=�0Np��P�M"�%
��!Vڳ�sWy����	Qd�����ǹs�pu6�i�z���4���Ư�5@�1�\UUW�*6� �ƨ����r��m��J�,� 8@ǿ�Š��Y&�o'EM(�2���AtC�x�����LEQ����{�9e-Q�Y�k����l?���Dp��i��tM�G�A&A�E´ǠV��D�4���r���+�F�֭��6�� d�>S���#�Z�e?0�:t1���AT�:�`�\�h�n5 s�`4�'��H���4�gM�Ͼ�#r��$���a�X�������9��X]U�Fp�}9j0B��R�6ى�0��{���݉D���n���T�e��]���d����}�!&j�T+�Y��������E�8d_�
����|�f����9rh*�+�R�aζ��I�.�;�e$�Y�b�{���ǖ�&DV�)��eSlO���=��� �YT �^'�I�<���]atc��8ε,�MX�ZO�1ص"�^؈"�+�e� kB#d��1%X�}����Z۠��IN&z�JsM����+�<t�]l=�,����3T�#M���8#�s.����gG��}�wG`zS$^�ww5)�t�I�Bk�hb\r�3i�����g��XB��h����}�ώ�I4g��<�A/z�֘ [�l�<�j�f��)��� 2U,�B^��D_X�����U��媀b9��Ș���˷�st���Ҡ��pڶ(o��H�� pqrf�U���g���'rވs�..|'�N�4�FH;.�^���8;�L?�m�(�hN�b�o��?��h�y%h�4v9}t9.>�0�0�[b0F��q2���}�Л8�p`@��b`�s"�`ʾ��%�Xpb8Q W ��V�F���hQ�)&X�܆0��kc��k(����m8�����O=Uwh�4�u��j˱��纅
0��
�n=��n;��ƹ�;t� u0Q	`�AI�a�bap��"��g���C3��	zJہ�"<*�LXE`�X��]���7�t���:4Z\Cm��( �t�K�?+�QB1@2\��@�/`��� �଎������A���@���&̰]��	��=``�.�k�
���|L�����g��{: ٸ�X&��y2ӕ?�V��B�d[:��)�::�������m�q�s�I�_���',{]C����|[@��³[Y� &�)�[�u��������l0�UK���4�YC`Lh��Ί:+W�e���/�RJ�2�>̚�i��)�Z,W�
�]!3�����hf�z��{��������*�_u��^�A[ǿ)�iM�v��5�����Б@�CW���$=�,�N@-<�Α��j��Td��j�������p,�B�w�E��ೢP���4�m1ҏ_�\� /gp۩�HU��s��i�K��!� ^����]�	� �(��=�;����=�ȟ�8E�x�e�=�K9-h-��@�P^�X��	�>��n����ڵn��W�ɽ�n���.���q�bd����DK˒����8w�D�[��ԋ4�zo@PK�(�В@�\L���0 "�;Z�zF���5{��� �ϋ�a�|���(7 1�%�v�1!��}�L�$'��)h��a�� ��7aJ0ϐ�.���2sV��A��uۏv�K��b���X�@*�Х �w)�,��'H�a�ŉ�r0J���0B�f8�:��D�98�H�l�LY�Ѻ
L��vp�a0�����p�c+�@o~󛽜'`M�b��dUU�J���`�[�����lĄ�X�J���U���F٪{�7]{�z�@A��+�
�O���Ŭ��g��� �WH��|��������X�,-���
�� �	m	����K�� �a�dk��D#UhoM��9zR �3J���θ"mX?���5M郄S���@���b���3�I��^]N@��B��2����6z��� G�ɪ0�{>!0ř��8��0p�̅�a#�60P�-gI��'
Y��^�3�8����S�L �i5�f҃��~fG��P!��ٜ5��d�$�`�T�i V彺�/U�`�µn�#���'�NG;�:���3/<�
3�3d4q�0�*�p*&N�N�W9&�
 ����\� �1�WO*F�  ���w 8�L1*�*(�q�Y�SK�[,��Þ	�y�LPX�RWL�U�f���d}~V�Y����s�]�<�/6-�m��p�;�<���@�;��n�B��.L����d�1�+ա"��-2tO�^���p��0�#�<�L�l /o��GN�&!�e�}F�<���0S��g6��X��
���^դa��Ga�$O$ S�/�j�mV�R�	�|�4Aq���W������Orwwk��286�v����f��x��?���X�)��H�Y��	oY����|�iƆ�r_q����7︡�L���c�Botwoi|W
��h��L�e0��Y��U���u�BV1 %�+Ѐ+���b�h����w$v9��1� L�V*�{�~Y�Q�.����hGaa4x�agkF1=T�խ!C�~O�e�������X#�4�#ٞ���!ڧpf\��6�I��4S����`�5"�xh� h�Ju��S�3�<` ̤�,0�&i$V�����}�p��,��T[ ��#!�TB�ɮ�읓ӓ���w���������8#��0�l����dqZ8I��`*�`t�b  B�EfaU[� �ʁW��נ�t�ɗ)�	  tͧ�àA	mL��"��Lb]�'�)*'�Vi���k1 ����`|8�Q5|̏D>{և
*��ӎt�8�`wi�ɶ�岁�q	.��9ֽ���R�ݑv�ve��� jW�;�G��15U��]��"`�F�����9�(0z�B�ce��{�窃Ӈn��+��k���c�ˑ��������*պ.3=KA�FV$�_|��&$yO)������B�Q@:�6�׏�L��Q�C'����$�/�߶�Y�@Ag�J���p�w�BQ�Ny-&����Ca6^ !Jۗ]E�X��Y��g[(�:��;��B�Ҏ
�1�W#U��CN ���9�Brv�� �c�'Ǉ>�bj�Y���{8��D���"� b;�2����� 5�GO���"�G#"+�D��0��E!��.W`��j��wy�/-J1IT��eP��������Q,ܘS�u��z,?Oq�ke�-#M�0h8�,����J��o�YI'܀Ux �d/W�v�zv+}�p���$�zNt�מx��5�@~W�6���Da�Е��DݕK�'�t���n��g�D�����긨O��чN��a��*b[�ɫS�5�R��l�d��W��xH�r����c��
 �UM�
k}����;jܴ���Nn�2�9Ķf@�6Q):��Ȩs�+�{��8�̌$4�� ;���T`g�e�Y{<��iۄ�`2}�����(d��dܩqn�-�qZ��XqVք'�k�Z�݉~l��04�]��P�ii��5��/lC�{��VhFݝ�^�f�O`��&k��҇	�H��Q��-}�ܻ�qlwo�v=��"�_g�����JNQ����tk$��L`��` 6r\��`@��1�0h1 ��A�|9��.m)�ה&��Ʀ #�p���-��"��i�C����)�`��D����oUC�}L8�D
�It���t?0����7�?��o@�{u` E���pL#�d`D����,���V�rQD>������'�6�{3?���,��D8��U-�����&�N �Bv޷��*�9a#WN�����J���&Z��6@6�` ���W�*����$2��m��2�Wa��5�ܺ�rP5�s���iw�-T���@:��i��J���F�߯L .dh�"D6P- ����$א��x	���N��h,��diٯ�}�K�����+�'o{�h�
 �p�t����4^��N��&�XUR�����=�P7}�9�B���mU��=K8���6
�3�����HL�m�
�&�n��F*A�X'�َ6u�.g镔���s�4�z�D���h�(�[hd�m
�R����`/�Q���x���X��F
>c��֎'_���Q3�9%���b�b	ϥ�ޕ�S��6ה9��-O�(�� R�ω�l�3c���̥~y'����9��u�
�Ǧ�W��y�`�YbF^|� D���%Uf0��a���`�h�]�~4(H�T��*F"!;m�MEd��j&[��q���ޛ���� ǖ	qꊬ��1�Ѹ�Y"d�@��9�pT��6c�v*��h����T�� @ �`�ȄX�}�&�'��S����\X� �f�T�0���d�,�>�(/���5"R��������X�zl��� ��!�����'"l�k"GSy�H����n��@ġ�dZ�Ea�ؗ558w�o["�C(Rk���r���u|aO�RaL�K[W�
g�#SM}�(􈱎�9Ja-�u���q|�q}��P
L��<�+ S�mW�Iy� ���q8D�=�a.��#�&#���=�|���^�ה���<~�,��� p�?S��ۦ�����X��B�m��S0R�5�Jtž�
#:��!9}D�1:�S�(',�� ���.����j��T}O���]W?j U���C����b�
}���a+��mtt:��m՚���Yv1�Qy�)&Y�7[�7��3�"�K�9�	@Q��XSl�>�7� ~g`��C�WM!�e?4��n��C���|�گ3`����E~%��ַ�u+����2�ՅM��]|ld�����m��'�5L�� 'fp��._��Z�Z@��o\SQ4���`0ӌ6�Jr����[�=���41ꆠٳ\�(\WP��퀽��_X��� lٹ���h�'�,;�S�U����Ύp����5ص�ߎ?��q�2�#��F1;̄�)L�wc0�c���J,��@I`�#�m�&V�:�H�/��!N�N6Bd���mq]�<��D:,X" ۧ�j���x���s�m�@�AZt�{Bi%(&�F(�D�&���~0R���RUS=�г�A��6��U��	�����@�R��b.v.!/�9�&`���>S�U�J��Cm�b��v`�
��"�8�L�A2;}���]��0*&��LS��3�Nl�Bsd�%���D]E"+˫��2����b�ۄ�4AQ��U5�dK��1՞C�� ��T�/�u���x2<�>xl�{��0���/�eZ���18J1yڴ
X�MaM����S	����X�����0��5&�ߠ�ב�ajlD�y3�q=v�p��AT� �|�y<k��N�T6+�=�g���1�<�
��Y�q���W��g�2�����G>|������AZ:���Ϡ���{Ш̱�¨4n��� ���L1� ��G����{�*#_�ꎴ�{�+�����2ZY0�;H��D3H��
(��`��*���#ԒBQ_X"�|s�b�m�XW��83�j����(��$��z;�S3`f��щz;��ωW�g{y�J��5��F�@�Ch&9�!9�c��TqD���	��t�f���x�p�S��Si����X;�����e�Ez_�p̐�`�Hh�J6o�c�&�^�Vv-7�s�A89L�R�Д��:Z����Zw)���'��Spq��4%4r���2�t�T~���8$�G /PgV� ��DFY�l0%�#$@)Ud�m��g(�L(���zD��ԏ��STŎ�����߅�1d;=���J=в�ܬd�K]y�� ����M &�FɄ,��p�{��F�1�(*�2@���g+ l ���i�[z�	w!E�5aG�d�7Lb��!�Ƹ�#�(�qsMj�c�)EK�%aRٟ����׵�%@4E�;�	�d�]�����3}W�U�F�<��w����əki=7^M�P]7vv�5�b�/�/K�"������/�+=5iv�q��Ԋ��ȴ� �oX��D��H��*�|%�{�+�&�E��&������g�`�;�h����_�-1�(��_dOᐭ5H'^(2�4cV8��N�'�i��^�D�;���YI8���:t��<�$���X̀���C3? 
�W��	Tqj��Q��S Ŷ͙�S�m��u��p=)BS�-�(>2���9Sgx�]f�dl�D<^5��/�񘈭���r��1aB���8�*%ן��E��(����m�D��ġ��-�.d`�L82�@��"zW�v_Ku_�+#��|B���Q-|�mH/�u�:��B���"4r����b�� @���a�wu��~��K,Ccf2�e6��. T�O1�|�8� �A��sI���fV|��=:�g�n
�g��Aa���dBO�&�Tf6��9��A�X��o�W�,z_zf	�l�_ �ܷ��LIg@&�p�z�#m��ň�����Ь�+Z��F���2�=��y���������� ̩�;��Zb'|�-W�=�4&��N��C��l4&P�.�sa|A+O�=Nh�&�a�߮{�p�l�3)[�gl��sh)��y���o �5t�~�U�=6i[q��m�1�',�I8h�j4X�C�P� UT��(|�5���vv�����x1�X�Hz��Nc��l"���T�Y���-�A��l�C�A"���*��0�>ld���Ġ9�n�0�C<�I�D��/���S���x�ڟ�E�0x�4��v ��!�BYhB`<40+41R�)؈�	� �\��5Ʋ[��0Uo��P�Λ2�΅Y3l�B8HW��6qp0R|-K؟҈xf|�� 1җ#U���L��p8ݙΙm���1v��+[�L(�e���)��1)�d�D D�hz�=��q�|}�t욉/�l����b�y�]��{|S�2��}�� ���&l�Л����c �WF�L̂�:�P$�f�
�L��%��	�j�'�nR���	�b�<�M��u�Eޛ��G� 9	4 J ^g������s�C�BS�3@�!���:Vh`_~,%seA	@���q�B[�*yl [�g͖�1���0b$}<�x���@�v"�t_�Еq�06�9�����H�	����g)\ݟz��yR\3۩{��	A@_�+��oM��qa*�0	��Y�<7�bn�Ygbô�Sun����R`����yn�)��^g���+�2��Ν�K/����;�-�Q����H����n��IQ�ٕil��ql�
sE8g��j(͝�5�Ll�S�������c��74f����n\&����Lx�c�dM&�h���1��w)$��w�\��D��t��"��L7X ��!��"�ȩ��6����~��S��\��u	�9l`C���
SFU_���a�N @#vB�b���|-��q&�G�-��Z�PV��9�/�(@Q�w-)&����D�K��p���-}�C`���q���

�#��b�`�zPk$[Y�.�'���s�-���}�S0S7U�}�XN�[����!̡���� b�Xr  �T�OG(1��
3�� ��L�"AhÓp'�J�A 5��u����OX��Q��� m0 �� � �����:s+�¬Q�����2��N�B�0���L �l����\�T�_)�7�C�����)���� ,^ ����i;+�u ���$�&���}�R���	�:-~3�=��T�k���Ǚ��2�"Φ�P���]�|��C�CمP�L����2Q�nE�P��y��2�3������q��ݏ�?���������B����+M���_���L���>��坤���z�UŵfY"�r��Z��Uk�!6Ŭ3:�S�g�^hX6T8�ң-�֠����O>�d��3@2�}B:i�e���ĘZsh;z�,8Q�}5s|����؃g�4�t��[�]�C$t?�Ǣ����W��Y)�+��p�� ��?Y"|f��=�̚���<ps��^7�w�i�0�3�t~39��
�ᤃM�p	�!+��*��0�*�ϡC��+5	f	��lP��&�Z��9� &3H7�� ��FQ;�%j5����̬��j퓙)�#ˋЏu'�p����5�2ۧ�{
'H�S���x��>wM%$�M[+�"�.�m� ��HPz���ˑ�P�X�Sc�
�j�k9F�b���w�+�����N�v,���Xb}�HhxR lm�� �L�B?n\K��C�<�Ҕ�6�xb^;s�*��[��;�����9#�fq=�����8u��7��Z?\�&�ǹ������4� �I�A��"y�Uc#v������m�i�Eff<�1ޗ\@p& �=�f'vg��C�K%3Fc�SL&�N����t�bw`��UU�u���'t�Z�1�*F׳�b��@֍q�ܹ˓O|�����=�80.k{�>-�@���*g��������%�3�6:fg=���/��(B��r%��r�J�RB(������Ѻ�"���o��֠����<��n)+d3E�v��s�n d�P�wO�S���Wl�P�@��P��Ԁ>��5NI��T�5?׀�HV  ���~������ ��S��c'�eP:v�v�ϭo8mr�A3���N��-Z�șu;��333Yfv����Yg� �u��0��"|����[�2K�����u��¹���(�({�R�T�L���֕2-`�u���VTrJ��m�.�nL���|��!+�W�D�Gf��9�\�,�D�^	���@�!��D�S_�'�:���:����Ț�w�C�i�奚3��Zh�B�]�CX�a���Qk_fU \4�=�0` K�,l>ӎ�[�#Sz\}�`k,�z���nw��C��{0&���J���8��0
  ��g�@�T�'@+��I
i����1�G߃��b�\"A��`E_��~��{:F]s���y��(Lɂ�>�uFI�
�tu�W�G�޹A0��U�(�h@��@i��UA,$ڹ�h1� \`��fdޅ��g��l���g��Y�s�i?��EF�0�^��5s
�ҎF��g]�h���~5����������\��B� E��H�����5���ktA�� N��0QA�D�8Mfu�h b�	E]������:���X��!ϩ�1�	���V@�����F�|�1�6�i!3'eN������ƎK�0 �-f�U���M���;N$2��Q���3������ը#åc�1�v�G	jGlS�6T��'�q��d��L�@��� �,�Cf8S;�2$LM������2����to��!���К:��!8������iqA<�e�� 
���*n�P�I3 ��LÎ0:Q����Z
�:<j���2c � V
�(�>O���h�2��u)-jĚu�l�C�"�ֵ���Y59����dK�6t��d�����8�>�!*n�*��DQ�1@����0VY�YԕA��!j��ǯm�M��by~|��1�I�ޓ��+Ƕ̘�m���'�J�)܆��݊F0~��Ԉ��q�y�hz 
{�U�ǅ�=!>����=1{�C�G_Eh^eO
d:��a��:��b;"#��Ge�c��T������N�g�uA��C����N�U%F}B�S�a�t0��T�����콹��g��LSc�:'~�TO4��T޺�^�h ��~�_��v�qAD��+�z��̬���g_
}����=��i#�]�Q� H	q0u;T/�绋�Ϋ��D��Z�T�T���#��~H6���ر1�qE�D�5���p��HF!3���2Epz�����`�FӢ�md��#�vl4 G�� rf`}��̖8�"�b�N�܌ɂb�G���O�	[q� ��2��1k���/*��2h���|�2�R0,��RLF m�L56if,�N�[���l^�ې����7��)��s R�p�΋̢�b������� @�LQ�%��\9���8.���)O �М�� H���>7@	f$��#U��.#@�'G����C���;��> �a�oD�e(���E���H�O%ciR|Q)�m
���P{�I��IH0[]�E ���6;�H�� �{9�=���J�,�I�s��~-�f�sܻ�����ٰ����2u�s�=�.��9	��6�6�l��Ϗ��9��T�B� Q!�д��	{?�^���i��c�}�gඒ!�0� �b�d�E��vw��t��R��s��< $�go��Y�&+ �x�J8�ֿ��@,[Y�Ǻ�4�E�@{��-�@�����T��BO?��&^5��s�3���KZ�N������
w1���`��`�x1���icvX�°;��	<C4�����lIΞaHү����D�-73v�����1�2P38WF�+E�#j�8�E���#Ӌ�r���	9��U�a���'���(G�fĤ�� �}[��X���U�.^�l������dj*��z�/ε�fV-k�h>7㔎ƀ	�c�3��������t#�Z�$���̏� *��	Yy22��H��1�CvY l0rv5��	�"tK�;S����k���"^/Kh0�����ԮYv�~7�P����:G!d!���O��%���2�=��`֬Ŭkxf3c�"
		��`X(`l�MpPDR'uWwuwuW��9�;�������=�~��J���z�[_��9�	��g����`��q��{��0U�{�� q���t���7l'GI ��^��W�m��o�����@��=�I��F�U�����H�� 2(xh/������p�nGx 9c `��ԾjXBSC߯q�L�ܺN[�澣�������ަ�x�Yd�yh��CND��n���Z�Qi(�׻x�diV���lrj�������{��>����� �|��	���?ಢ���Y���v��ڱË��p�4����;h�z��ϙ��l2���0I�aM�b�6��^��y^�/�k�@@����Y�!s���� �.��W3�b8;:t�=¸M�!c��Ƅ�h�C+��k��j{@���- u���a=���|� R9��<��c����X4 g�-�y���ڠ:b�7�;��Өw�ԃ�(�����
��(4@��0ߑӆ���i'ܑ���?(!�J@���}h��0c��Z���V��>�
��@�>�@�2{q���㾡w зfW�\�C�[��[$�N48j�_J�-B4.���z
!�-�J���p��r�|�z��0ϴ�/�5�h�d��0�>G�N�*�|��hmj���Q�R�����ʗ��qj9N��@]��_i-@��{���Z�V��)�3�0�.�Î,��/jp�l��唁@�t���"��*��8�j�K#�N)�Q�R�X������ 0/���ȳ�:�/i_��8�S�p^�]eZ#������";&M|vC&�Z�*4����/mL��D��B?5�R�v����#.`�#�J;{��������@�[�
��3�=��&�r�� ��y�1)W�;+��ݎ��kݰ�����nm"`�Rh�&g��v$/��f�ڭw"ϔ���=�צ�z�.6�:`��a��h-o���Z�*:�_r�f�_L��ھ?������ �=�~�E�v�L�k)��w��w&��^��OktWO����g��T�;�b� �6��+�^&J�3������T��h9������a�����rH깫�,�ߡ:��LiC�#.&#�C0轜�N��E�|FP��w6*��L��`1�8l�؁�\-m���a��̯G.NN��~�_Fva�i TN�0V|d�<\���g�	9������X !�[�Ll�EÞ�5�p�D�k��gGv-(����2���-T�w��@��<������c'��=��Gst�Y���. �Z�E�����\�4.��N�r������,P�z*]��b���g��9���|��Mi3��}Ε��[�
u�?Y�%��-@ ���� B� E�w?�Ջi�Č`N���]�> �0�HJ袉�$~�F��#�G�ZՅ�gw������6�#��Ի���3( l.в�(�:�����0U�Y�U��^����VM�.0�DԚ�!�����Q�� 7u�9�5�`�=z�r'�ֵ̇���h���X�]{�\��vM�lw �\���w�f�r��*��N+w�e���Y�S�͎C���ǎ�,��8�~�����da��Þ{�߸T� |Ɇ�S�5|����w�X�<�T��R��k5�s��{f78~�Ɨj���?e�>�Fl�,=��47�����D��&�A�n�Zs�*@�3�<���'qL��J5G��N�K�+`�2��AЫw��kt�L���h&x�l�t�ct8�����2�55�������c�\�~��/=�����0�|t�>R��bR�Ο�8\�9zO183�3;�lL�{@M��#_��4 ���G7�~��=U��d2O����C���s���ț���G�^��<0d��v��C�pM�	�s�������z�9���=���&%ዿ�J.�����7 �1P 8I 4�D�R;�� �ޕ���9x��-���G�jt���:E;2�\\�"B��]^�n�CZ��h�ݤ�f��W������<2 ʸ� ���@Q_h�ڡv�wT���8%wK������Dֽ(l�^�n�>�s�:�,kd���)��W.ڟ��D�a����� ���C����t�TV�
Lx�����QRz�
 �@�����B+��Z@i�Я'�P>DW��z^�sW/�I��ٻhqv!� �ګ<G ����#��H$�~ZDW��v��~�2<7� �Î��\�\`�{K�v�so�ʅҘ���6;D��g�yBs����Qe.�V�c��+G���]�.����Ɓ2
�lThh�3�>�����I��FVm�W>���k�)`X��-��;���J�{���J�z��Q��2�>�����XmB⥓K���O�xN?���x�֊ճ $u*�E�c��r�~@h�Ƽ����|��>A[��]�i����}u�;q��}0�K%�<�0wv����1Q��wL���s����E�o/VF�=�
?�Q~G�����8�bLDq��3f�+�>�Z���n·������Ƈ�}�N��ٍ]�T9C���oY�K�^����fh�F����%k�o�H�N�		ˆ������cο�cc q�'�(�d5�ä��g|^�L���Duq���hSX�� A��-�3�G��O��@$��YG�_�x[��Nf�݄������牘�=畍�='��kS4���c���}�=r����r'���R !��"�0���[�x���;x�ڧ�RC�v�n�� #�dQ������= �vC�4���.|q��8�P����W߃�f!9fT4M8f�s���K��X�v�SO���QG
 Lq�>�j;�1�ak#)�7Vs�C��Vq�����}nd�f<��:z���3Hr�M��|�C_�����9�l��>�H���:^3����
�Z`c?��2Zt)M��� ���%�R��ߵ�U��p{0���¬��5d( ������j���@W����q�#Uj��E��ڠ\��+��܇�����)�rn�T�f}�/ml<�@�[fF�ѨTD��o��Ï�3_)8*��f��P,P�0%|�\d�����F{m���`�_<hl�����Wc���)�Aw����؋��|�cu��!�jz̽!��x��؉�|B[t�4;�'���xx��
���_(Mu�/�D�L�}e��t�q	�BGU���߻񮷽}��C�6>�On��l���n�=� &r���C@�\us�B�� a���󎐨�u�9����,�D�an)�O)�::�FGT-¯���B?7	�0�-��o�N-����� �R�8��M���O@�z��SO�;{X�ڜUma2>�Ȯ����vC[6^�j����(� �n�h�Ցg��<5����_�8e��$]�P�v�ǿЌ�1�-�� �7$-,��5j"]Q����"�~8	7�Z�qG���;vv������r����fxB�e�2N������um_�&�U�U���D�-��+娖Zc}.�-�AF8�`6�h� �4R¦��M5+�,�%�j ,�ݾ@85��+/���i'�V��)��X����U���3T¿M�4O�ۋgZ#ÆgꞾ��媗��hÚ �o�u<D�����N��|���1U�U�'T*��}񥍳O��8���Z�9�ZfR	쩲{�h��A뼧��YL|;7���t��K�
?�ê/{J���Kt�G��y�
����/#Z~�b����Z���v�'7k�2/^*����V���f�����s�t��m''씗Ge�3#S4�:���@�3v��\řbD�d�����ɭ�5Z�
�W�kG���d��/-�q,� �c�WF��N�!�L8������xy� a�C�A���"��.��Z�����rpp�Y��:�L��j�[�?l�s�Ww��S1P���v�O���^�1���m����E㷭�D�4�c��;�Ш`�-�����g����LӀ��]j43>�a�N�%u�u؆}�� 0p��6��uˏ7罹v����,��f�ѽ� �qт�9	3�1�����������C�#�`	���0�Z��V%�	���@~$^;(qt���@�-CD��?�if^߯q�t���N���e��o�����1�;0�u�>]n�8~/�Q��T  �IDAT gh��wX� 	��vH7@�-R<`nm)�,@�uP`q��aA`b���¥�pUh�޾��b��q +�8��_�4v���Vo���Z`�7.9G�a����J|�8�3H��erV�����{�7�J�@x�"��eUq��'>�G��X�Slt��QpC�i�%9"eN���>�c1o�a�\��8�B�d�>s��&��u�S`���)~����143��cj1A
B��`��8S̆�)/U�캸!�΋w���P]�|N:X�O��ٲ4@�	jg��	"Sr����0Z(>8����~��T��G7�C�A��;;��q�$Y�C*QM%8��4>�� gd�F���od�٢G�� @C���j7�>*;�s�  ���pB���Meɲ-oS��(�f��.���x�m�<��<�g�+��.���m��r��5�W�ZA�4�O��͛�y�#�eB�����H��Cs@W���- ���l8�ͅ@����}�*+���Z�a���pGG�/6|�:=O[�0�����Hm0��oW R�-�]�>F�:w�rn���i�m���ȏ�Q\Z?�����Oǉ��A�!K?�����9^�����D�e��,� M������5Ne��AS.�7I�O����>�^�O��}�X� h�����g�6����	ĳ!���i�K
v�p5�-/׆�BE�*MՕ�e�.m�	����L�9\f<6Ul>��ԗ�̰�,��s A��B���;6����(���o����C (���}�3 	MX���k3��ų7\���yv_��v����*���`1p��F&�f`*�pL�c�rLy���{�|;D�r��� �	�P]����{l�V�<�RKWj����P�7��� 
ڿ\��%j��z�ą��G]_�tOEȐh_qy@���Y�L�%�V8�v. |����_�H��媍���'�n{Dr�d�����З��m���4}�� @�M��ְ,��ߗ�^�{6�ȨkQ�t��3dQ��3���W�l�,��n��v��UpA�~::�[xQ:�8Z�G�nl��F�qw	��S��0�u�]d�A����m�33� 6�s;�/����� �����#<�����pa.�Q�C��P�B"^�ռ"�Z��OM	��rѧ�д�e��B���`:���J��K�S�Z 8@ǿ��O	����oM���E;JH8��GDk����	+ڮ�	Ǎ=��,�N�� ���@<�؎j�cd��z=�x;GU]#Y%�#���� �jCPZ(SApO�,X�y��|=�dt-�̐��T=_��Q+g�;�q�4� ��'H��l� ,�Gs:sj>27^jr�
��f�eExU���:�3l�.p�k�ڙ��a��u�L���A��|���A��>ïb|%4��)ߌ}K�(Ζ��Z����>�@�;7vf|���T,��D&#�Q!�G�$��#clE��XN��Uu�Li��@��s�Y��0�ܶ�E�n�{r-��\&'��K�;���R��̉��I�}.��)aB?I��I�b	�������Є�V8`ihr�,��k����Y�������<��:���l�&�����?]������<�h��RXK��h��h������a�^��7�K�#��Χ�B��X��<�zF[\�e�e (F8"��m��$F�$vd]���%N�o5�g������X@	�_��Y� c�c9N�h�
�\-���ͪ��쀅Hև6`�w4L� Z$� ���|8�d@`���@�jcg���T6���G�,���뾓FRo�C @��굊��9�P�I�>	\Z[�Yk��恝g=;
D]$Y$��_9j-笡��\QK} 0�X�֯�{��//��ϒزO�l�Mȳ�!z�zu�k>��Խ�6^$5Ci�\Z�Uf�=�j �1��V����@���9�P����v���l4h�6�#B�̽�>��/|���#����.��Aw�ľ&ú�s��:�5�sϾ��L�}� &��/&���#b��C�����~�r��'�.��Bu/�:\"0�;S��{~���x�+?�s���
)9�a�hz���hL"א�Ț>�����Ju���	�)���J�q�C;C��A����O"�"|R�-L�u���A�n�"��>u�;�\;�`	�K�i��R#�㈿j�@��649CL�W[���8�.��\k���a�{�?^���l�Y�f¥AH���b��tԇ�d���ku�]�:�������2R�A�V=�]�^�fԾ�B���5" ���� uN�֐��'���
h���w���pLtX|x64��/T���h S���6U��/�&2�����pҧg��f��Z�{F6�F�}`*ڧ�K`���>���]��]�k_���0�\-O0�js��2	q�)e�y\��f;�s'��Ⱥ��Ѧ�z1hj���߻�)身��g*zUΕ��Q�� ��R�-�S[�%"��~��N/��H y�|a �z��{v���bmBN�����������X�94a���La�>��h��=~O�|}:!k?R;6sq�3�/a�!3a����T݋�?t�1sϗ��<������.�u���{�~wS`����}U�+����-�3x�ua_�ix
<��� <�|��`���wmU��r�������9uƶ�ہy�,�ҽ��|'����p��?���ƻ?�6͑]�|��Oq�{1�]���B�_�+d[�D�TYɾ�@#�sZ�˗�d�ڟ�ߺ��)H7����>�tϗ2��4��C 7�~��ȵӦ�����J�Ն�5�'�3|A��` 	ܦ���X~iI�� u� ��X�M��:�h�,H�ϻ�����*��6��mյ	������5f����!��@.W�>|�Є H[->���]Y���k�)�� �m+�A���oD~3fk��Gl�@-ȲG�hӂ}Z��>�>��3���R�x����/��>D�l?"��A�*a�b6F;�w r}��_��}�hu�۲q��{�<;N���UgG1�h��cm�&�4<$����@6l�Ғ�׭ ���:G�Yks��]�J뱣R�(-�ZO�JCs�0��J�J4W�{�>�OWT�ҝ���ϕ6��9P	Q9���|��[9�8��'/V6�3j�s��s���\�70�ﬞ�$?��̱C7�x����o!N�$��@U$>���+����*��z�R;������"w����\c���wx/���3t�ȱ�K�?�}��z�xʁ�]i9��|���j
�A�]=��np��ڷ�����RHN���5�;;2 ��N��@ ��	�@aG���&������b��	�nB�I����KU��Tws�L��b~�ю�����l)����{J8T��֬<u�2���|�eZ&��;�o��s����v���Z	�����:[�Bi�j��@�?B���:2����>�l CD\g.�ޑ,��|�����଱������q�?�rM$M��zU6���w3��hc$��pmv�MHQC�(�m7�#[�+�,W�^��a�x,ڡM𳀲�����Օ����U��_,��Ȃ\!�h�J��	�h���N-�Qfh����ʸe���� h�f��'=�a��pI�&�~��h[�M8�������B��z'�`U��QnD�u� �0�b&16̿8ᗩو����TH����I�<k������f�L�)���*S���a�pS���S5Po	���Y4���O�FaǑژ�<����8U���P%`������\9�:Р�����"'&��u��)��W�w N%@�y�y�LWdnF�Ucyϻ�Y`��֨}��K�� �t���� ��=Np(r�����8}�Ri�!���zΉUc�9 �o���^���O6��'�oq���\�w�L�3ö��օ��Ѓ��{��S(�Aw�L��~~����~���W��E[�A�;�>kg����zJ7uBT8�:D�b:vk���08��:�sq�~�b�w�n����C����CՑ/���������su��ʪK���:G���:��v��)ƿ���25�+���W6����o��җ*9�� [��nA�#�r�,��r���\'�}(+f��X�+30 �1�����K�Uiw��Z ��ї���9 �(��~S�h?@�}@�� �����25�$p�\��dD����5E�Ve~`͗u�oC��jx��Р,�e�����0��W�����8�(�w�ڽW*��E���ܽ�i�VחcZG]������W��C�Y��km=_�d���e�� ����u�ƏW���7��P��!�  �ʄ�絯�<ī�	A�u_i�z����W���0D3�G��y[�WGi0��~q�j�^�84A},i$d,�M����@��e�ׇ3�j�/��]�)K���Z�<?=Uէs�+��s�!��uL��g�l����a���S@�@29W�gt2����i�������j�0������� >>A�oKc�g�ԕ�*�rўCU��Ov"�D�>�π�=*
�7E���bIG�{�c7j�l���L�v֮S�_����`- ~ 0���6S��X����a�C��K_F#�x���^����y���;J���8^��tlsQ�?��X���zz_��
�쫿���'�ju�
k?�b��p����� ��,�a<��`֪���f<u;6�Gk�/�N���Qq���4A�F������9�i�^J<Z����ў��Nb���}�ŞL����<J��.�r��I���b�?��7�P�VGK�t�DjKP��P��I���=�4 ��c����tt��{���
Aq�@���j�N�!����ġ�6�p�Ugѧ"�:L�@���\�@D���Tc� >R%?0[��t�����4�f ���[��;�t���^2gOp\�C8����
�u�1��E�u�	�:_��O�����d��l���"&4L?��U��g�ؔ]$������w���c�2�@��}�S4��p�������fNV���9����*Pq�"`����H_P���u��8Zu�:�U�¡1��?N�g��V� ��;v<��`�A�H~�4=�H�S���RsA]hR��߯�8��B�����H�B��v�=ܦ�v���Z�/�IV�6��-?��ڕ5���,�0�UgJ�s��5��t_-m��R[�ڱ� ��>�ss�xk����j�sSG�cD��vn.mO�=tmmm�y�@����/�t��v�d�Ҿ^���s�Ζ��gfW����z��~6�I�D�5&��9dw_�Q V����e;�y�_���Ts�����qձ�u�ȳ'*(��%`�y���3x.z�T D�?_��+�~a���ς!�� Pm�Xk������m_���%6K���a�r�������;���n�.
��O���?����C�d95ڜ0�!��#�y8`����
��BC팠x�监��1����6�A@�P�`bW�Cjg;Ƈd��~50��q�3� ��j�����c����ĉ%����;7�����ڵ�>{j�P�4 R.ո�}�FZ��OË�5�]4�����L�̞-�>�I0��3����?c�EEx>�,�B ��l�pډm������9_�≑���(uN%4QU��k<D� p�� ?��^�3܊�Ǘs��T�1�!��;�ˤ`�����u�4j��C)�/�@"J�����d�I����s��J[p����%�Є�|����䁕��i�-��p^|����Q���e��� Z+�B}�9��mG	J@��C8�=|��\�3 k�]}8�7_g�ўuw��!CG��ٲ���:���o��6���<�M�;I�5��Z�	�a}�Dx�����e8���Q��s������s�:�!��p=S���0��@CR��f_��Z�}lDVƁ��:D�)�h��' O']B�G�a�c|���WT�6�x�|�/k
`R!33���X�<K���|���!�D_�M�}X�6w��<Ѐg��>�\t|{X�l�j|��Ə�)mm.[��\������a��T�74E��Ƭ����y�����̷�bԃct�aх�8��/�|����������]�v��G��&荣����b*�aV����ڙ�(���r�q.�p>0��@��f�Q��Gv��O����S0H�&rj4Qe�+�.��=�X1A �X�J'�|�a�[�)P�ر�g��L1�#G�o��b�8ıv�{�3�^h|�4$i<�)�������?\�����WL��K/=���Cm<S��pՉ_���=������m�v1i�*Ъ5`%��V��p
X	���/)�q�V��j�Sc,���*L}	�h��pou���%�ΗV��E��X ��Վ�V��銬�d�{�q�iȜA�^z���R��p��E�4�j����:x�P�=���;��%�'5�*�k��|?��"Lm�[#q���^La%$�?����o_E�\j'qljd`>_	�Jx����X'5'Uׁc�m:��w��}���ĉO�����O|~��Ͻ����S��}�+sp�{��+�X�=�so��ھ�h� �y�Е0n�4��W�qeE�_i�N��d˹� �`����Ʈ��\ZfT�f���c�Tfb_��b�s�X�龊4z�;�������½��x�h��������^�m_��i5υ4ԁ���9p�����'@�~. ��������NV�i�Y�4��4�uZ��>N�Z�=WZ��*�Ţ��#� �r�K�����:�<K�O�E�R�n�~���tV ���^�/l�<s���3/<ӧ��9Xf�b�����g��j��Z'ˌ��~;�9�v�(����fx@/胦�px�����km��?�9�ud�/�h��Ľ|f�A�Ks�ku}��_��z
�5Aw������O�����?��ezz�g�Y���!�9L�1Df���%V�3y`�\�1��6F\m��#6�=�Y|M��*s��&��y0R�#D8�rÁ�a�9v�v��}�Z�'�}��?Y���FfH}�I�^�S����S̩�ܹ:.sX�ٝ�%������M
�_DY�yg�Ud&�v�A1���N\CC 8"���PU/��1�'�"t�q���U� =) B�D�v;�֎?�D�^�f&h ��'�S���{�&'�� Wk
<��NA��N}0&�:��ڡ���t�������1!�_�C:*�����G�}E�^/6���.��k��c	�{���lՃ���C�ª��_��4@�Ҏ����{���@��T�GA��b�2��L\����K@}<P`��ڽ"��:賵[�� 6c^X�!A�Ҋ9R�`���ߑ��P�%�?q��}�s8����8� �%��X`����5����k�o���3��;��f�	LgDx`^.T�X�Ҡ���>Ʀ�~�G�[B�{�ר��6�3k���[&b~k�n�M4?�/�U��2��O�c^�7�<�<�9W��>w���J��u$�d^�0繁�T����$���g�:k����3�M�|�	�����5i��G��I��w�-Mf�E̼��>?�.Գ�������+���$
�5Aw�l�ƾ��;�௓�h+���C�¹7�q�� U�+���f�m!HP��a@�(��ƙ?�� ;�]ϵ�4��<Df��4iڻ��7�T�J�W�)ߠV�w(��2�<�y��%�`��r���;Xc�Ƌk��C �=gJ�Y0P��w=��t��������C1���F}j���/G���[��A�~�)�>�� ,���~O@	�xq��G�7�d���9����S�(˹I�ZR
s;i�y[��}��_���Ϗֹk�w���tQ �8t����C�9��@�ቍ���:�\�g
 �z�=���'
�<��w�3�8\�~�[�cU7Ω�3vU�\?X���)LV7���sEK��* ���ϖ��x���$ՃF���Lhe�a����}u?48�⅍�������x��|ql>��Ig��~4E����N�Hb��=�q�� đ�c#(�BiW���q�=���L��е�{�_�ٹ�n/pZ��	�A+t�4l��Ϝ�1���oG��Xo�׾3�+�́�{�4��>��q^V}�rmTֳ�s�DH�lP`+� �kNHL
�Ô�|��=��۾q�y��>���5�Z�'�������~��R����/hCك�6���}��Ŝ�κd���L�ћ���.��7�CT�������S�N_,��BKM�hv����_�5 p��#~4}u��Nw 0�W���V��H�h�-f�k�G86d�]��z
�5Aw�������o������D�V�,!��p2"�dd|�A�� ���Cu+C��Z�>�;B���ެ�26��Ώ�ӇI�ς�3�<��FlD��b�k��bz��?�?Pթ�}���x�De��������� �1 jQ���G��/�C5&"�0Wi�B�2Bq9���+����7�$h.:O���8�'cEà�j~�=�� 4 V܏� 0��qC��� :��GMm���`�ȫ�ŋ/ֱ(h�Z�V��A�	ta�m�~R��2�l*���[2Nh��c�v}�.D�����������  :�SQYП����Bѹ3�֮��>�G6NT����� �k��t �`��:4��l8��z���m��T��⥢�!�{���)���Ρ��������K}�s��g� B?=؂��֡Hk^qL���r�h�yǷA�$c�{�̝��Y'��xFI�X��15ѷ�5dz?Q�m������G<�5k�qu8<f���E��7�;��e�c�K�d�`�z��Z4|��������-�g�G
�s/�[{�h�j|�����&�?�L���*uTf�O�]���Z�3'�Ͻi)~��T4�$�ߞg����\�ɿ2�qGݵAw�tݾ�����W~�O��O�u|����F�M+�L��0$^�.���! P�.��`���,樷U8�%�^�?�^�Z/ڂI��L���&
ã0B�&�p�y j���G1�!,*j�48�v�I9�g�kMM��G��H,�"�U��\�C�?�3����g���R¥5��<FF���3�8�vh0� |z���Y�Ё�TuP�ѧ����G~�Ƴ�=���yA���y�K�a`�8a. ^�,�<P�oG�js�}�hA�ɏ:p\�N��Zab����ȼ�B�� ��p�3O?��w��#l𛹷������|�\�&�
�c@%�i�2ƷW�r;�Z��5�g�����p���p>n3_�g�P�@��"�d�S�Z�(d���@4�5Ⱥa�<��CmVBx��v��:anT�?��':m�;����m�3;���^^,�Մ^�B��ڬhN�Q5M�Ǹд2�΢�u�:�l04nm&j`�e^f=4��U��^L�<S�:Q7m,XoD�8Rz~���c�C[;���M��S�PH9u�HêKЈ��M��;��F_�=}�xP_Gw���ȖY��9Z}Bk;��P���6������
��O��y�^�'��9f�
��r����[#K�r2_�m�}���a�O�a-ez�7���|(F��v*$�2>7�2/;���.;Y��qz�VL��"���0W�{�b6Bx6SG��~����?����<�x	��Z��<�������>��T�+g�/n|��O5�������M���`�A8�{��V{�Q��μ%�x�ɔ\-�1IԸ��~P ������=%��:]�#�����i>���'�TD�<��/w��Q�\�k��t_1�/S��v��L؝��~��OI�h2��Gr�@�>��]���Z��o�E���er8X�r�`��]�p�)��h4*����t �f���{�N��^*p����*	&��|!����ʗ�m�G>��]�.P��#�h�J��!ô�裏5]�+�p�ʿ�=��1�S�
�Y�M0�A��CxjƠ�/V�4?Q�_��t�����@!���N���+�Bg��R��O���W`�rVD���S���SE�
������Co�ul�S���E;6"�������~��MǺ��x����\�f�>�.��B ��j�3)�����ƫ"�jh�|�X� L44hj�󭎗I:J������j�g����h�<������5�y}�;�TG�ѐ4�����qm�3q�D3�M��3��mPa���4	��W���y�� �J�\|�x&�?�����˱�uH�?�Ac�C�X�7��&�~P7��v�:&�� mМWյ�'~�'F2��뮦�ZtWO�+ܟ���?�ħ~�����@1�h` @��ۧ�m�;Xt�X1w[0�����^����}�cݱ�2�fg'p�y�=1*�6�� �Y��ns�f�& ���{�͈��Y�|�����49�`��Cg'#$gZ��g�d�7�F���W�*f-E�^hs֜�j��Ѧ�*~�^�v�as��� �����R�l�a:S�%*j ���h��S-0|h��%�=�����'j�v�`i#�e�}G��G�����K��y�.mz@��K���z��gJt�����y�W��qa�#���ja��¡�ϼ��7�W����C����аP?���K����2��Js}іjq4D+L�sj�M����e�O��h���s���H4T�4;�_���go�&Z ���)Qi��/�<�/�R���^X}|L��Zd=1��Es@�a̯�*�_��Ӈ���굃~���v
�>��CMO�����i��i�K;o��?���������pO<Q�mK=� ˞���-V��&m�C��]�s����g�6�%`L�c�����|���3L�l\<ڂg�y�Y��P���[�a�A���=��$_�� ������>���s��x��ʛE�u�c;�m>�6�V$%/�ۮ%�� �7�<�����ݿ��/�忼v>���L��&�n��W1��a���&L����+���T�`j�2Q�b	�}�ѷ7��Ri(`�^vn���Q�R��N��R_�f
c�A*��?^0�O}�S�P۔���U�S�	�`�#���OB��߂�R)�K�@�h���y����������	ƌ�/u2vs��+!c@�܇	���TY���%4�ဋ#��\��@G��g%P���mA��8��������FH Hp�e� |���Wt'O.�_������ =^�'x�v��8�>Ru^�xi�2?X�%��
�k�tЊrN��v����i�4\��Ą�g9I���G_�U���V������q�&�g��s�q��Y����)#�bG\������x�`���/F��"������U��Zh��R����� 蓀���|���}챮���?;���-���ʵf�悲�m���W�#�f�����w)p�@. 7sw��	)� k:��l0�ñ}����o�7 ,�IB�G����9b���ڒ�x�̢�/��/,�H��) ��k�l���uj���mޫk�	��z(��7Ľ��#5産^��Ǌ�����5�_���]�zW��g�ߡ@�>c��s��~�|֨�vX�h��/�����G�N�]6,��:��_7':xg�2�YvU�#���uWS`�	������{�����?��O�����$�����H�:P�ل�0��U-;T�v;�Z���Na�U�����#j�s�W$J]�ɘh�Uer'G~arf~���嚪y�7�!��(�����#�A�tDM��ЭOB��J�F��4�V��zk��1#� b�C�)�N���`�A�5ڣ��S}�܏@��A# 9\�E���I� �?F�u�$�9�t�E`�П�|+hk�ۥ�����Ec������� p2�
`�_�����>���'����d�y:Yڐ~�O�Sh������27���2g����{�q�SGV�q.���D%�$���y9^�% ��Z���/����vW�;�\���}��8�̍��4���K�!��N`�����5:ֳ�;�氣�J��6�1����P|�������v���@KFۘ�Xk	*�*R��
����}���hI�ֆ�/m�h�w@�=�J� �C2m�'5��s;c���Om����hh
� 8��WsD_�+��z����1������LR�g��Y3�wn��g۠m���Zkhd��Ѡ�i�\���Y2��3��O�AO�s�o�fD6��)7>A�y��N�;I)Q������������W���q�~ݵX��ߵS��v�̹c�a�BC#�������4���vw�ȷBh��ʗr�s��(�����@�R&��)������>Q�n����,�Dr7�{?���n�<ڇvl.p�Μ��\p��]�*M�;˷��m��]�q ��\�L@��`���x��T��ɣE�2)3���!�d�&^ N�
�:��?�&�>c�N�.��D�K[�YI��@y�4i�_����B�\"�|�mչ��q�S��ǎ�Ke�����)��Ea�_.��n��6���lC���U'�֬����ϖ���_z�i�� �&�~�Cx�l�t���e(� �]` d�a��4E�j�nHH�o&�q��[�Y#�� 8h����z�V�� =5����u�8�XT�y���F���j�N���ꝺ� �f����,|���?_�l�K�lhg/} �ՠ
ZX��T�Fspk3ѲY h�y�^ BA3��D��H����@(@$��5?��e��q#E@=�=̖�녊@�Tˆ������e�<��q�8�@/ �4�_�l;�37<�hO�X^,�"�3:sC
�/�f�}�x����Kn�3�+r�|���dNި���i��~\����c�1%^;5�X��M�E4��r�.��g�M��A�N����^k���S��t���G��_����|;N���qR�d�� �!ㆱt����L�aȪ�����1-�����|�wј%�(���,��o�M�0l�Ծ���N�pjU�:\��T0a�U��Β<�ˬ�g����s�n���>}�ĉ�o�>#Ѐ6:�;�E�O��N��yS��@�ߠ�;m&u�G�}}~j}����@H�!�.��UX�� E��^�w\S�@�E'�+���ݬ��>A#�!�aN��s�>I5�6�-�;�g���#�Mhl(�iBS)����u�� ��*��w4^�����D�ڢ/h�>�O�:u����w��>�&@(t��Ɨ�#������:ҫ�Ϛ{�Z��jL:��Bs�65���hCm��Ua�Б2�c��3&~gx������R�� ݌�1x�1wB�><� +MS���+���,`V_$��MMтgٍ��/���R�)��c��ɒ�dD�l:�b�[���~��"1��/4� J6�;�&���$���5�6{c���Zg��0��9l?����I�p��������7�o��Á׭�.
�A���������?��'���N�׻�� ͐S�C�{� �I�Td�(ۧ��tq�F(aʠN���Q�����:t���s~�H� Ӈ�R7}�eFXmw��e��Ŝ#����0a����j�]/s��j��J[��hu H.U��ǜ)|�h8
ׁ�%�� |;|�����h7l�!���>Q�(��4�=����X5h���6G�ͅB��)�	uJ�G'1\~�Ff3f|�IGw }�AC� PѦ`U�`�J�8 0�]����-�f,��p��xD`�h	@����q$�!c�hM�Y��:"dW����m�����I�q��"P3"I8�=t`�N�cdͪ��f�4;w�W�(�rc!m���2�uC�?k���#�xo߶z)F�p�#�_]Rנs�x̷���7�Y6/�	�jV�:t����g���̧?�s�I�9ħ���g�v����y{�> L_'�Ꮧf-e��J�CT�fn"�p�h�׉W������p�ZX���Qиwώ������/��o�?}���uw_&֎�/�`o��%@����Yj?�(`�����f�����HLȂ ����wv����a
)��B�
8`�0Xځy�$'^�Qm�X�X���P��������%��m�Z���i�@�܋���S7����?��ʼA��c�V�D8ir$a���(%��qVuc.A`P�B��i�{�O&?��}0k}k:Zm�FP�_�ݡ/�)�����w ��#t֙acس�.�N��p��a��(4��D�@1s/����8 <�'�Ŭ���^�4`��-'fhGt�oSM͍Ñ�Ħ���Є�S]L"I��A'��_�����������i���Ӯ�[ԉ�g�A���-ְ�p�M����7�O�_L��\�5"��a��5b���<�gh�Fƺ�'����n���@mSkf\_ h�3�ڹ�Y��v;�yх� �{˿��V�O�[�f�k��w5XБ��m����e��Klu�ya]c��h���Jw���>�)�_w9�>Aw����� `��<AP���L�#Q`鐪p0��G�v�����o_x�����MG�]��5��LP�F� ���&A�N���*�`p#�`�0d8f8��(0Q/B
f�X4Sp�#((���#�t��{��������;GѾ:��\�ê(�&u"�q T ��N��LG���;������/ƅ�ĨI����41�I/�	a��C �m�g?B����F�e���3�F�p�g�F�p�Z0\�g#t L��R)O?)����}�=Ƿ�����߃0ȕ������kGY�a�x��W��-T�>�3�	����F= Bʘ���D��z��h�z�G��Y�40wj��:��1:����s����ye�Y��@��3�)Hr0�>'���}�whB֩��2�P��I�3�q�k�`�M=� 5��_���1S��A�D�6/�?����;�~�[��式I�%x��	> �0��X�5>J|��_���%с$��C��Nx�YD�Q��L7`:��~�Hmr�����}w��;g�nkO�����~�Bp��Dp$��N�w4���Ɔ�0W�?�D��5��9�4ID��T��d�ũ�Ih0��NMj��Й����O��a!�.
��:���~F0<C��qcGȁ� ��=��4��5Ri� �"Z�ˍ�H��6�T���D����Qq��?�s��uM(-$��@�.�%ҁ��,��t��>7}�]���5o�Y�����P��(=h�}���Ob\�O;ԯ6�q�;�LAK�e����M��� �@5Jj�o�}�JȦ?��-��$BD/Ɵ�4�Ͻ�q���B��u�`�s�J�m�we}:s����2#�N��0�9���G�;m��p�?�}d�0MX{�Aw��Q<���5����Y6���<j� ��N�-� 5��7A�fg�a �&M� 3��)�j�N����a���c��Es��
��\����4F�$�d��PDy��`�+x��07�Ws;�v�̉�_��������}�2�uc��kM�m'���`���;x�`�^�����V
c��
�`�hP�#,�ӡ�GB�9
�a��˿r���c��ɇ���e#�F�����S���Q,��)̟��w�0`-B������Q#`5�1�2n��j��8KH�}��GT
|P�W�����#uCa�0^=H)��!�:���	4�i���zhvd� �= 	::?����iD���k��1
n��������q��	Wv�c�τv�G�Вy������A��:����OSΰjJz,� �u�0��-l1�U���ڤ^�I�o��}X����k-�����qP'��G�i��i)��6(C���'��3��8����p/k�q��4��d��`�P������8�4�����a.X'2��åz�C|�ӵ��_����HN_t��-��5��<���6��Θ�
#��#Տ�ʬ~�@ߋu��~f���_�������,��[�t)
͉�]N���hJo�Z'2�♡=���t;r���C�"h�1��W���k���w��\�u/���?�;�m1,,�A! ��?A'S��P�6��!�T7���a�0c�~w�0z�&�;�U!�=j`�q2�}��&�a�K��qx9���4b0E�4�A�L�]�^�35^ ��iaX��z�O_%�c�0��ݫ���0�a��o��q1�_us������3�ZA��t�(����ۡ^��͝2u��,���@�8��Oڢ��APD9�1"	A�p�;�:��� ���$�� �df��^QA�U�3�N�П,���1:>���I��_M�ϚM���w�B��z�~�"@C�J�\*��iBu-�Z��X&�n#�t����ԆaB��j9�����`�
��T�dMp�!����t�yc�	�߹si�f���U�)kG�%M{:ĳ����H�Z_�=��0�U�+��'>�D����~�4Q���؏�s�s�&��U���5A REB��}1w<��������d���t"���?��֯��ks�]=��|p����?=Ua>��~��(�_���d8�N��0W7Lf�y�����h2�i��5+Kb4�I!��.��̦���w@�3`�2�`���Q��5v��D\������ P���$��;�����4�!����#���z��n���p"��{t>֯�~ ,yir�	M\0kÖ)���H�å���{��an��{t����H-��B�x����� �ԁ�a<��4,���m��8����U�����:�7������ҕy8R�3�j��6�����$K#���8X?F;I���1\��I9���!�>X}$]���:�L9�H���J��y�A�u��ξ�����'� ���Q�z��cd�?ƨFSm ��+��eMm̓�ej<Xs�	h�6�.ڀ��ߡ�Q`Ҟg��xq�� 6:�3��	���,��kG0"]�^���I0�S<�S��'}!���!f|h�g�,�їw�9t��]��AU�薍4��7FFo�K�.m_^6x����{7}�#������?�ʹ���;���;a�ހ>֮z_����r%!�1|`F��,�eǊ�s����Le&��;O��Bƥ�\�SX3O21��(�#�(��3�s�� q@����B�z
`�y;xW߭C��}�������P�L!b�8� �i�\���#fM{��?����.w��J=�{v:��5B�r�ܡ]ƉfC����������d�=�
ho��>A�9i�ߨ�F�#'�3����kS�y����3:��/�}j����1My�i�c��]��	$�}��]�} �[��i�p�/֩���� �iM68��}�;�FG��d���T]�k���a�q1_�I���xb"n�Uc���z�<
��<��[C���.���VR��#/�-Qg�7cƴĚ`2�j�|���iF����h�?~g���<��E(�P�nM��������.�������35�hui�w"�\���0:Σ��ߋ��Y���t�q��n̘OhD�`Y��Y� u���a��q���uWS`�	�����������uz�>2��(�2�W�m�q`<��K2LBAcw������h0O5�̱#H��H�ȻB�ߛ�-a�0g�+����~ H���4$�!&�#�ݐy ����|�		㿿�͂IbJa<���0�s7�����`� ���O��
���$|��#��:\ٰ��CC^�ES��;�d��?:�R��WH ��*5Y�}0v���N�i����y�et��3�g^ ��B�k�����.Ήb}@#}��V��Mr�e<��?4�8�}�9���A���Ժy�N�G�7x�}�ɚlg�2��gַ�u�g�y�����Wӹ�eT��� X�O��sE_���?�O�s�}�#߹�>����3ZB����dk�����������KS�e-�Cjp�3��H��k�k>G�ue��2eq�q�CߠZ(�Y;&,em���S���͘y�d<��}���v5]7-�c2�
�񹷞��K�D=�a�j��0r�5��d=b�?�����w�r.���N���	�t������������K�SڟR��ܹ�}.8�;#v��ڄ�ǀ��H�֡�LV#�`L0)st0<$�_P�o��M�f�:̻��l�]wr
f}3�Ti��j���՜�	���R��F�ٌ��J�[��z�3��ӧ���ٟ��
vâi�?��P�vt]i.z&+�_�Q�Z�_�|�3.�޸A͠q��J3A}��>ԅ@�����Am��D�d��@�9~ڣ^�v���Q|�K]�G�~�t�5���t��<賝�k�!�Rh���{4�!Z��c��p&7�4^�)��Y3���-�±�콽L���+��&��C��3c�oB��Th��0��C������ys�1�k��2ߑ`^�	")��*�2� �~����d�6�t�����thZ�k�ܲ^{FZ���fN;��~6<ܛ �瀗��-��z+-ԧ>����C����	�t��I��u��g�ĳ&}�b��^�}��<C��c���r@��Z����TG+��@����x�{����g�����w��m���f��	�����;����ZaaD�&����3�b]��)��aަ��I��00f3'7� $� �e�
̆�~#0%��\��2j�����4��Om��Ӯ��0\^'��"��ݫ�4�J�cF�S�h�A��?���#��
�U����Ԫ�u(���Ι�EV;YM,�oZ�f)#�H)����zp���hZޘO���j^�Db �<�2為��}�A�v ��� �i�5U5ƞ�/����65Z��:���!"�JXq����+�Yc�)c�)�L�;'�_:p�]b���v��N���ip�Ƅ։~9��]Ƹ p����T#"@��-#����B�j�n� uj�e��S�b�#�܈l���~�/�z����n5' I ����lD?j`���f� �h`h�{��[@�6��6��_ټ�����̥���%��'|׬̽�����j���t Ci��|��Z���3=��������r��?Qs�Ϛ;�����_���G������G��;�g����)�A��vw������������>P ��5
"`8�&i"<�y�*tB]� s��#��i�QK�C��0j��yX}� �2�fȸ�P��d��m����0E����0GM>-T�ѪE�d���z��	-�ע� ������x��/T���B4�˧t�Ѩ[�]�*X��@h���e��VH�&h��A-�k M'�����ň�}���As�n��rF�YeW.e��Ք�]1%�ˣφN�m@y��r�A�tMW�#���C[�`�a#R�uz�2:�7�4E�S�yyv�`U?���\�9�p�^�,�&�\���'���@3*cՏ��45�p�/���0���l��@?�F1���K�#��U��s�si�$k\`M;�� ��I�����0y�ɡ�a����B`G{�o�냗@�7Uh?KK+����=�+"U�A��8�g�p��>�B���}�7M�m_��kW+������{~�]���<wM�5f
;�W�s*7�(�TX;���;L�c)�:�9!`>0#?`�0=~�OB�w��"0Uc)ý�|�8�t��w���rM�^ꗡz�0�T ��x�����p���y�o��M�st��K�D�0p�H�C@�f���Vԣ6�pP�?� >Ͻ��f�H��t�P� �=Q�C��#\h���ӹ�v�����F�%4���9F!�Mȧ&���x{i�>�Z���m ����.�R&�C�`��3���KMe0�i�jS���^� rh�a��ݩ
@�T�� =Y��
�Y��:�����M��Cu������?���w�g�<�_���'�A�b$Z/42�}`|�ꠙy�x�|�XC�F_�����0.�mRF�L�� ��_P���nht �?��5��g�VhT��5�9�C�O0'�l�Y�ƒ��A[njXk<ǚØ�#ڦ���u
mReo���ô�������d���uB�K��߀��F�@��k�p�S`�	����e��������������
��8��bWGT<ZK�������?(S�X�&#��}���]ޅ�\H����H����	L�A0GsQN��b.�;i�!�Iۿ�h���Q�E$�?S�� *���:�&�!F^�D����h��D�[r��j}��f��&Z�;m	~�p��A9��lƧ#)4�}r������H0ʵ6��,Pd|8�Y��Q�$}��S�c�7F�	�Dg�5��B�W���q��I|�*�u���6V�1N���+m���|���9Xk^�wƧ�͐o׬���R�jR/}�b}�g���ɥi0�68�̀G�Ў� س�v��-ߡ'����Ǳd)f����8"�M��<a�a����N�<�]�+����s!5@�}�~�̜Vj�x>�'t��Љ����3��:tt�7��3kz��Nhr ��y�B�y.;If���d�5�~�;�"��衳5�9�i<{�E��TC�Z0��c��� -`������"���r���~��~{�G>�kL��/}���\�.�-	\��/\���?�u/���o��(�Aw�tݞ�~�~�o�����Q-���2O�/M1���/�b؜���P �9F�Dv`x���p�}{�n�fE����:�JP�����-N�G5����	C}����Sg]��;?L��[3�N�0L�����J���0��Z����.s�A!�`,��P��Aϗ����t���c�������D_=��Pb� ��P�t}����,ě&��Н����C_���H�g�g�uj������)�}F�3@�Ƥ�@�%BZ3\��Q���A݌�$�>��a?��5��y�2��c-�Os����1�q�;��H�!�-�# ����Й�4��P��J^)@6���4w�S� �)����>�8=μ���~?��[���
񇶞g 3r�"��K��4%r4Z!}�x��|0����������G>� Em��q��z [����i�x	��5]�:�&B'�o���0'F����^�g�y�~}������%���~ �r�B�*Aڠ��0�Ƃ}#���Lϛ�>6��iZt,�zb}Fϟ����L�9$�yd���@|�&O��Ђ?�`=�J g|�!���E_����ڵ������ŷ��[y�(�Ao������?�=���~������Y����9t��5��@�RL!���;L����� M&�=��52ɮ=#2�K���-`8 �3��L�J`�<4*0d��/*��N����M�0e����(�du�4��`	�ɟ����|�3�A��+��`4��h#���pk���±�ZiSN���Ѵ� �4F{�Y3��ʤMxONIV�_z��5�hs�O� r���r�F� C+w�#a��9RL�D��PZB�4�7%x[X՘I7���_.3Ngg޹��s�Ƨ^��������/�9&�Ў�U��8}G��)�~���) }��ǽ�ϩh��B������%Sp��8@oN%G�1�C���X��,ڦ�귙����Ǐl\���h1�0Nʞ�>�~��\'g��S�;Q�|w8 �fah��}�yo��'Z�t?�'d�.:�!�2��}�����jm8bw�+uN��X;�%� �_(M&ZW�}=Z`z�. ���-����]��=U��re�N�p��ù��w>� �좹d}���᥌���k��a����'��>�/�~�:s�&�t	��O�G��_����6F�c1#����<(�u��g�2��Z2'�Xh�}�>��U�=��'��3~��u�^
�A�k@Ļ��?�g�ķ����_�����7,��@9�����fV8.��o(ƹ��>�r�Y�����])'|.c=SB�5��ђ��I�����L��C����RB��ei�~��)���� 0�:�l3.u��R�r�Tg�v�r�R	E�{�T��D��
cNۀ�ϑ��q�։�o�H@��W=:��>?�G��i����"+� ��a��5<������8:"Y\ڪw�O��*���e�)gq�&�Ӳ�߮Ґ�S �̾$�C����B(t����d���hJ8���`�L�<�RшP�{[@�栄-���% '��T����^�1��ʷM8��G�[�\���s���m�"�=V���T���}w,�� ��^x�����(8��8��� A��] ��E_�@�̩�콿�X��U���=��5o���q�-G))p�e}������Áv�W�M�� �ѐR_��8�I=�s^tA��� ���hۆ�?��zY�GJ;��3#}��<k�a��=}z8���A�:�~ ��ځ� ;斶Xy��ָܱ�<۬;���}����$�����Y}���? ��#�~��L�y���a����W{��GL��������B?�x��g��ȋq]��l�E�BM�1x2k��`��C��N�t�گ��*��ٍ/|����K?�>x����x����W�WP�O��?���'����Ї�z��bVhu�x�-���؟����F*x���`&��Ȟ�|��8��5�8�Y�z(GR4/�0$�9�J� Pt�ԼAY���2x#t:��" ��}j�� &�%Y"�	t��g^�	 ͨ  Ǖ%���}�9# h�s<D�,������Ƒ�7Lq#= ehD=�/J�E��vqj���4΂�f��Uޗ�#y#��M*m�*�e��`S�G�<�ù��i��/�$:�� 	� �u0�ٳ�Y����47,n��0�%�A;b�W�b�I�9��px�/h��V�[-ڌ�kb��kM�%����O��- ����A�2�k��qUϕ<n�֑r`�	,��Z�������ؔO��;r�P���ʈ>�ޡ�K�ڠ�O��8�e��Ǵ����_�9U�I�f�=@s�|�.��Hp��Z/6��̓X��@�ZL�mfj���MG���[��cݒ]�~�I�5�Q��ރ}؋�L��,��8E�-@8fܼX_>����n��g~U��3���8����i^a�ct`󎪯۪u��<N��_���/�YAc��О�&����ko/�c�������.�~ݵX���vj_�������o��������+s����GSZ�!�n|����$p�Tt`3T&t⥓��/���ǳ�����j�g�/�2��
Ԏ������a��a�|7��F�C@_�d���I��ڗ��P��U&k��  (��q>y~�-�ܲ�A��a�ԏ��o�}4�..9��P3s����C9{L�7"�T���%��X����ƀ]��� 4؍�]/��MF].�H�6R��=�_x�Km�$l�{;�z���\��������)���W��v2G�])�	��
�;K_5Ov(�"�lZ��_
4�EC� �Vg� ���D��Mt=�i�	���V�����ɋ�J8��Ti�Xg��]/����^Ύ��O�]i�罾Ǹ�����P��%9�>9�R�g��-086G��N�Pu0��?M���{��>k �����3��ʯ �ڐD�뚣4C�G�4_�x�Y�K+��`�!/��֔uF��ƌL��wKp�Xi�g���;s4�th�.�Y��������l�>������K�G���H����ѯM����9����i8�ď�ȏ�ks��w%� 讜�W7�����������g�o���3_�8T�d��N��0i��Q����!�PY뼼o���� p�q�n�{;8�X#���>���aRԯT`>���H���Sw�� �Wt����&����?��1�� T�aJ̴�awZ��f�.�����K���Q7��i� �>�9`n8�R�6��`�܃�hZ���SŨ��w����=�B] H�M�`�,i���ü�1FC��s��7�tZ��e��G��������#n��-cp���'�]¹i�&�hZ����.�U·�A���i�Ԣ����5�X����z. �C�<Ln
`.`��h�c|���F���-ڇ��C3�Әkמ�8kp��;4L�< Y�90s-�� ���f���������	Z��gw���Aa��.��l��u��3��0^kMK��Xk��>�?�5�oβ��`��f�yx5P^ 9�EGj�N?r�F�@���l񔞓����븞)���`^c~����#?�c�m.������T��i}u�*&y��%4�+
-L��.���oc'j�ڱ]���A8]�{��a�u�\%��D�\��������E�`�����> ����e�@M�� ��Z�^_a����&��W��F��}ڌVZ#v�W�I��0�Ю{��:h�σ90��̠z�Y3>���8(W�#��k�Bս�MG�`�i���0�&���HK}�F|�<׾(E�+�/��	�7�����bhg��E[ý�-):r�|��1�O�A}�q�a^4b�u������#Hf�a�d�?4���`GY�@D�T}� c�^�ccf�m��c�TEVg�'Ia5�6�"`���A�a>�>S7��S�KJ(�F��u�Og1�}~G�u�Y�)�C�m-�bB$S��J�e]�o�OM��S����;�<Ɲ ��F�����D�'�w���t����ѿ�����J�/��+�1�Y��ת�Ǟ��/��l,t�^K ��>O��5J���.X/�֘�bن��f9��Z�����z�.>K���;Z{��>̡���G�2iV���X��e����sߵ9>��)�Qo��>���ж>��w��:����ML�u��7��Q]�]��>���^L��;�fԅ�ءa�t`�*A�� p��.����d�+�p���54h^�nT��ap��`P�$�?
M-��n�Ĳ�\�_��PR3�}Zv��3�sW`y���5 �l���y������,�چEKa}�#�x���@9�Ҟ44~<�g���+W2|"�F�zh'b�>LUc������ۥ��`�-@M�m9�Gz���m�u͇���9�3������M���zS@���P�q?cV����M�Z��m,Z��M��&�4([����yr-n���6o���"x�j�լؾR��g��h� ��{hX�����F����/ׂ�Zwk4ۄ7�AjQ�ϋ��uAy�^�7�S�����kTͯϮ`6�7���t��3��q4���/V�� �b��ՉMW;v^_�u����-X���e&_�q�ܱ��&LD�V����!�@BU?@��8 � 8C�8�2���E�9�*$4���V@�ȇ�`��dp~�\�U;�@Ü�����Q�U���T �,���M���k��ż�����-f��G5L[�a"Z�q���.�>c�[�)��O�\�C1�Z�2_9�9G�z�ia��/��tg�F�Y?ig�z)���B3��P�i�Y���GK� ����s=�*�^�M�-���o1�X~Ge�s��n�?�^��s��8p��k��a6��z�n�%4%������m$�P����q�97 1�H#Pɹ60����cɱf�{v e[����@h��$�W|�i�s&�s-���њ����m�w�&�W�`
�A�<y�W׋���y�C3�6����rw�P&f�2b�P������2e��u��Bu(�W�J�x���)�RH
خ�)o%�tl���&�[��<���M�RT�C{��i��+�Iw�
����!��ySФ!�P�6RKe=�#y�)SX�'w�)|�ys}�>|A\���Rka9�� j��Y3��������\���H�Ԓx=��9ǐcr���a��f��@�7�v��Uψm��s}%���k0��\3ع���F���fl9���M�3�X�%��3u�X>L�K�ت�m��]C�5�k��5�9���
ϾR�<)ܓ���d�33���2Xw�ޣI`V�� ��N��ej)p�(�mS�6��i'%|�K���	�/��uu-ʁ$�����$��&H�.MA�,5#I�)jx�߱&(IS�¤���LW�2d���Q���1B0g
2RK1@��~'�\0�"�-�@��	0��ضfЖ|�cMHΩ��:t��N� BЦfDs��K�Ϲ����w�}���6͊1�y��w�0�O	��g.�u�'��~��'�I��@hU[9�=��҈H�����T��9+[;F�9���U=�g��+\�� �]��+՜����T́���$�٧�(y
�U��ߒ��9�d�ԩ���I�D��7�ki�IƚY_�cK �`3L,i��kjq��tJ�EeW	m
\� �*A�t�c�݈�
	���Uڒ�K�F�	>r�ѯ����O�.\��dޟ>�^��>��r�%p�����9���u�oJ>7�G�/׆�z�y�twnf�J-������<�}t�� J`%М�v>K�[N����9���>Ϳ�lI�Uk=��A�2�ʄ׍�6
�5A���wNC���%O��%Z��g�����RNa"�K��֪]��p�� �S�Z�$�N�B������.�"���.}ɺfp"�qX��a�YK�@ɱ%�ٞ�H�Qj�� D��󚂝�阞����VMA�����@WG���
����rH��8ǐ��C??Sg�����a��*��I���m���T0�\��H�h�]�g��4o&@09�
s���6�ߗ����
�r��ܹSkbߒG�w���K������>��S��L���1����ܭ�]���K4��p�Uv���a�랾L
�A��$�[�x1���)�,q�ڵ�L�L&輣��#NБ;,�Ka�=��&- ��)�@�w�	Zl?�c��̼gƜ;F�ܦ�*�%(۱}��� !� P�@�Q�n;]��7�������4�Er�R �̴'H�>	����ۖ�����4�%�Sx&m�[���w�s[�v��oۧ>��뢶�̠�Ʊ�g~K��<�D��Jڙ�ڶ\��Y�}N�h	�����/5�^�%�6]�<G�C����>�>>w���u���y�9���0� `Jm�c>�j�E�\s	�,��Q�g]j��)l�r�y���D��[t����%�zث(����m�u��m_��;�n�@������2���/wc)�gM�q�����d�29�<�12�d��W0�0s���ʱw�%Z+���Q_��.��?C���V������XϬ-�qK5M��}�sng3hRx(������C:[��Qob5 CDR�W�^��Dn�~#_M�Q�݌��g�L���ŜǏ���%��8�]�F.!��HM�"�R���ƟHڡAe|��W���w�>K�M�V����]�U�2-Q��L
�F����S�!0�u#0��|�엀�g��i#��^�.Ɩf��j�rs�����������y��fN�B��
��d�w.�;��9r�2�?���������ZB��Xk����}ţ���Ư��ſ��m�� {�=u����>쮉��5Q����2OF�󕉛�r2'��NP��o���+�w���p}��s��fM_a�����Q��  5U�cl���#���f���6��8>�d�6� �~��*8Gu�0tw�d��Pw����M-�u�]-�G��`�Q�4mx�;��x�:g\��q2�+���O�>.�Cn�><_��t���P%j$�	�:gg]I�Ua�_���6�T���U����6Μ��xU�ʵ�v��r����Ǐuh�Jx�Rp���KՏ�umi�.��r�	��<6h��[j~���:Ac^��5M K���Q�2�/t�;g�qhm����<��Go��*�υ[��P0'��9�~+Й�MM@{��fIp���Ю��{��9��}�{��/v���ݵ�3��sC$�Sc�3%��'��]S� ���z�3�t��Vs�	l��@���ld��;ms,�7�3'����~vd���u�g���w����o�c(���1Su�;���W�h1��p���q(LX���N_���3_��e�2.���o�B��`�0,�a���w�y6�ZN 'i�Ra�5���EA��1���5�i*⳻M�;O�K�+�a+|��`]\c|��������
:t��8H�<�C}��p[hM[��a�#>S/�F}�j�Y6 �Q�� �&ޣ@LM�}�;�uh�4�����=���b��TۜT��rr9GRpfZe�\��׊��r��o���w��#D.��.���N��ku<����g7.U�+�9�G��B�x�B�X9����XO���Ρ�#>��Д{&}�
`��Yyn>?�O�T�8[�56	6՘P'�u �Y ͣ�k����_�"��u.��>i�f�g��Ú�	�5a��|�[��'@k,3v���<�vj0����	}�|V��2�3k��봯Ё�T�?��>C��{�����������o?�]�x;)�A���wX[��?������7��Ӟ]��ܦ��+Xe�0:��V��;�E�:2f!��p)���\�S�DhA���<2�4�O�&�ziGᡚ_a/���}�q=Mm�Y,>�Qx	 Z��Q���r�?ML|V���~�Rp8>��]��f�Ik�Y�+ �9��]Ӈ] ���b鱟3�꘎�'� ��ý��o�\�� ��>z�4>��8�h�|c���9a '�tB�@☔��˜`Ǐ��s�{��O�9����8�����I���E�H�UгB<G�a(=uH�]�Ƚ|G��G�8���/	:mSP#�A�Z2jF�+�+�yV���~�K��n��i�غ�S�������O�A$��>~4����,�.�t�h@SW��l@�x`����~`��3�P�L�o ���u�./7
>#|�=��S_��>X�=�����׿�c���L
��a/�`o����_�����?��Y1�_w��=���/ԩ������Kf�&�S�.�p���g�y��1k�W������_��ºˆ�i.�3��.��B�k���f��Q�*3H��
ZH�A��52��A���^���ԫ�75h	�4
v����u
4�f�ԧ�Rv�4}7���̶���Mf�҆��Z � �n4=e^��4�kFęi(xv�?Ʌ:���H�	���w�Yt�7Μ.�H�s�IK8�s�.W�g
L~�䩍�[��*���:�e���ߥv�:���\@�4S��4�Zv�}t��<���j�Z�@%�8�;/�g��U5��U@ ��~.��P���%Н�q��gấ�.>S�g ��9��j_s�86���|�a��l�ߩ�� :�,�4�\���0��s�]����<�z�{���[�߿UǺAoՙ��qS�����gݗ��/�OcD�x:�QR����h�hf�̾
p��g��
�L�vB�O&����	����@Fk۳߂䢯�I&+H�8���-+�=i ��Ԫ��R Q�>I���
e��H'ʫ�����8?�g9���ѯ���D�����S�9��cB8��4<�\�@@��rڨ��>Jd'��c��H��t*����8[>DM���|��N�z�>��P�2�*-N�h���x4F���Ur]9�[�K�	�����3���#�rn-'-��2��j�X��a}f$�ψ��V.5��G�`+��Ԝe;|��y#`�\	��h�S� Q`j�Z�g%�OMYn"r#!ݝ׸}s]���3�n<�����"�\��)�Aw��ݎ�>t���/|�ET�Ǯ;V��H���*��Y��Z���"�+rl2X~����5�%(QHd��ȸe���H���0���4%�l)T��&�,���~���+�faf��d�΁���H0���~�PKᑂ?�J�3p����-g�2��]��>ѭ��Y|�
�Ա��ꠏ7��遏cK=�k9�s�<���1�}ʽh�BUt�
�a�=u8m�h�s��7�.=^��K��jNuns-��J��P�L��8K���p���K��r��e���"&�S��N�[��k'���.)���
1F�3��)��	��td_����繑�X�z�=֙�;�|N�?>c1�:�4g^���N&</Ի��݅��Z�}�/�ɇz��/�8r��r�´`Hj8��Ӷ&(��Z���Z��PA�谛cH�A��0�	 jRdn\ל�`�w����.2h��BS��6`	`R�� -5M�˺�>ض�[�]�ý�n
K5LI缮��s�;kʧ��:$�����_8��-���8Qf�b ��P���P�2a�@��y$׻-g]��Kt�C�D��g��
#'D'��:��t�����z��/����.����U��*@ly�?ϩZ5{��U@����n�s>Sk��C�U�:���d�ڦ�2L�o�J����H	�5Y{�{F>o���g%��Ϛ�p����հ��Us������]�����ӿs��~�/�����ݻG��q�2��PP̚� 2y���T#�#���h�&�i��D�2�Y��)��Z"�ϝ7�ѧ,�BΝsB�q�j��� s�I�N�!]C�o��źS�	� �{��ץ���p��ԉ,�U���G<���ݣ����(`�V��$j-μ5D]\�F��wW4��cG6Η�IpE�;�떶^��HઆQp�z�=MSλ@H�j�vs�i���6ko��y��W�� D�E�5�S�W�S�8�R�qN\YN���r�~��Ҥ�f`6K�V-K9�y�+�� N�-�;u؏�3������?���G�JcP�����������ל��+|sQ`��\������k�������F��}�\;�/m��I�+��$��yˌ��i����P&���] �T�	z�g�Vd��Z�L1w��6�>��S&�j"gc?`~�t]$v;��G��I�h54��&41��[ڎP������oR8���N�HU̿}��$pt������B��d��P���2`���^��}��ƥӧ�i������ܾ�ky�mC1����#���`��^Vｯ@��Q@�� ��+�������������#5 /��#c��?tk ��	���8�r�~�qB�vBO`���#��HSʹ�3�,�h�R�@^͑ct��v�/˵��a��ip��ֲΘk耣;uv�}cSd_l�k
H/�J�S���:� �q�ƚ��_(�b���	ڶ\���rY}�H���~b����Z#�7�Dzm;��y����+k�s�{�vlO�d�%���#,�h0 ���=��wh��2������J���*ph�]d�ȹ'w��~0���/���k�ʝ��e[�=�7A��L��)?���Z��~w���1p1�ݤ`���]Ej4���;Z��)��m�Qب��B�k���Z�W ��g��E�Ӫ��E�u4�*A
�!9"��?^-\l� �0O�,��|��y~��5���&s6�ș�;t���`h'�����s�PϺ�l�Z�=7��Z�=M}�I���g>�?ۧ&^K�g�\����e9~�H푀n.;�9��f(���{�塇��w%3_�+(�A�EqKx���>L �����S�N��\��������I6�~
���`�z�����~��?'H2A���_���O_�OƞBT�!�w\)�65�O�f��D%�\Շyw<O`��f��L0���ǘ�|�2�Ja=חmTV��k�qj�ٖ��D%ڝ�ʥ�)�S��ꇽ���gW�ܒFV�X�W͕
�������NG��g�ȹ�C'Ȱܬ�4�1צB޵� "�/�%"�x��I�'�K�t�~纄G�V=�3(ʱJ_�4Po&6M^����r�!��}�����fc]_�;(�Aw�<����o��������``fa�a�ݧ9�l�\��Q�r�fB�� R+dX� ��-3�K���K�~�5B��(佴M�f@�ujB���̺�O���
9Sjx�m�C-T|kҹ�y�6;ʫ��!5F�����[q����cG7vT��t:���o��[[���e��P�#G�l��2��wog]v��A����U���o(/(�k	<�|�v"i��p��p^omOzۧ��t�������>|�f'�\[�_`�ƈ���6kO��#רc�O���x-}�����M���e�v�6Y׺��v����?�/o��u�;�7�9w��ֽM)��#������{�i�pȨMg��[
0&��Py���djf5|
�Ԧ$��$�L��a���&�ߍ�C�?��8�m����;�Y������
�G
�8&��<����2<�7}c�f�������<o-ɦ��0�\,�y_0E��O�:����2� ���j�a�q����aa�����z$��
X&�{9TҘH�[�s�ٶ�g�x}�1�;97^��sa�i7�ļ.?�Ƿ�5*������`���hI�������]G��9"��O>Y٩��4G��������3ꆃ~i&����W�����O����e�\
���ܹ��=��G?������o��#��p����vBxU�eL	Z�cț�n�sv6���w�	f ��T�'��/�1�%�'������;�x�jq��P�&����5�XLX	��tMa��uI�l�og׭���}U�������9\���h0��vW���:s�
 ��88���C#�����*O㝨�2Mo
�j��v�^|��$8|O �& ǨvC�`��>pٟ��y.s>�kl��;�4͠8�Q�-:r�`/AV.�9����u���Z��h97�e����䜽��`����S���~��������A/��u�;�kM�:qoT����ß/f��#GGdϒ$�]�&R�g�� ��2�����6axHs�B?�l)A�*&/N`#3Ĭ3�3�9pL	���m�fM�<�D�(����0ު&���(���	R`�I��^�ː�D
q�W�4����AB�J��`�3�.r�k�3���X~��Zޚ�zD��&r.s~�o�]�[^{9@~��i�h�V��쓟g�ϼv�{�U�o�*����ک�Ц�f"�=k��k|E����O �+���c�Ht糾��w5 ����?��u��Vx!���:��~� N�n��|���O|�[o��u���k���co�(>���5�k�dq�v����I��Qc3�QG	H(/�y�f���{�L�:L}�;��5i��Z�ZZ��{S}Ԧ��ERb�ޢ�Ӛ5�Vm���@�رG� �6�|����z��_�\����s�s����ҥ�;Lza^%�Ε�Of��i���J��Ma�_~��MV�"B	��\/�W���z�)�z���D���EOI���KZoZ�`���_��>a����u%���G�0�
��l)j.�T���z��s>��nڪ��0L*��(�:*��)����j/��TB�B?��7�7�s^(E�F�\��Q�ַ �G>y�&��Z�L�����n��\��vn��"���R���_��'z]
��n^�9����k�N����D��N�p-�g�ĻmD���ꆶ,!
����#��p�����r}1w��'��Fo5�2k�V}�6Bh]���}���Eƫ��z�U <�V�O�S0߀Q<^�")����2�x#}�6��|1���C��v}~�{���5'�$?���@ohw�ҟ�W+4J`$�1�;4��8S���"Ì�,���c?n��x6g����c�_�0�4p�������z�Q�I+���PkWa�b��s4)�����=��td��eUn]�V���z���!)�?m��S	($�K��U�9�[�6�aLP����C�?�h3==�h��]���ly7��Ju��t�S�5ۙ�[h2ۇ �b˼�1'�oԽ~�p��ּ���B��$��@]�+sΨ�ȸ�:�-���jݤ��&���}ʑM=�r^K�wW?�.XE��R�bo�'����7��
)oۇ��N:C��E�����0���sʟ*5��lx&�|��r�tsZ�PK�h�?�����M�e��i��-	�l�b�WՙW\@�Ҡ��IqDO!�n��r�;h�Y$�sF.��f[$��,?uѾ�����t���,O��S���g�8ɑj�g��,p��UY�*��L���dK�f������>)���3���|�^C&����:��+���q���%<"=�8��T[b����^gc�nnp�b�T��Xט7���y�����=�;ݖ�k�l�l@B�ǔ,��6O���R�QF��o����ړ�����6^��_��{L_�8Ű_�cyI�KW[�ٚx�*�f���"�$��T�*��N��/�Å�a91�T�S勒�6^�*�¬������X�r�j?|	2�U7 g�R�j�m]�93T�(�kY��={=a�S���E���h��0K�nb�2�ݓ�k�wϫ��,�51�$��j?����T���d�,���	���y��<���d�A�أ�K��E~�ER�6����Y���X�k|��Z栴�?߹]�1�R�`��_�����������M:M�&��B�\�*I�������a�d�3���Y_4l;� �zT{5|d����Yz��*`3�2iu��/Ua�훀�G��F�i�=Q���!]C�U����j..�v�P/����EA�N��k�P��7�a�Q��ǂe�y��{�>]>	\|9[�Q�K��d�ltU(�n�#pRP�
��Z�!�E������0�~I�����$�h8Jf��ƃ����������9�b�j�ϕ������T���1���3��LY����o7J6��ur�ߘF*09��-=!r�ڨ� 	C��C9ƑՕw5�F��!�:	Ɉakʹ ̧���M(N���Ķo�Tb��� '@�>1�V�v
NG���x����j𭒠Ȏ�p�PE5����˦��u�A�6�� (�$d��:���(���7�s`��,�\q����h=�G[/=���������V�/q��&�_�R�~��W)����I�r��&m�߯�^E��x�|Z��j�P�>���6����j%Ҁ�gp:�'���*���
#���Ԑ���*�	q��X��.�:%L�<0�K�:Y��)i,�l���f�p��DӣAдe�ȅ�Uq.B"I0��ʭ������� �c�B�Tl�7e[��d|�)_�\��F�G�V[s ~�͜U��T纣Weq!�����;�����R� ���.|�,�vX�;+�B?do�s�Go�-���#�=�����l�a9�HP�#�W��ي�1���	�tPM������3�l����Ʈ� #{j��hP����ϋ���{5��M�_��mmW��.�pDj��?��}ƞ���^���_~��.{��������#]�? � ��3���}�0��sM{N+�"I;�L�'�_r������s�O��_�m��$�����9�F�1V��\�=�RO��l\$�GA��� ���1�#oa2&P��а�3y�`�5�؜�o�I-p���!�����:��Z�nxX�'�i�����$V�(�{7���9r�X�1 ��-�������8d�&��zz�R�W[j�<ǧ�`����@@�aB�Z{��Q����H������)����*�Y�����D�Nf+D�7v8��sRe�d�?Gh ʣ���˚�ņ{]���}����ֲ��4!�
��Bډ�Dg�O>�2���@)�؟��[�cK��=�_��\P}���Ĭk��.q��N��p��_�+T,����+F�-!n���h�=��s��8t�Z9��B��$0C矛�<��)�7��y9;�"�3�n�ͨ�8מ������SEm�y��.Oٰ��z4��̺p���`ί����_�.�G�Gk���/��r1�ǰ��n�#����_Տ�x��ssnw��j�Om6�~��=9���$���9`C?P8��w�I������n�<����w^�����v��i҅�9�c2{	��K!�  ��78���	�rH���"�Z#9�(������yn��؜3�G��bR��è��#�)uI��V�\ă���~��܊"Mn@�e��JC������|�&㐞����DX�a�n,2��Z���@�%p�{�,��l|�z�	���S&��5+'y�g�?�~�rX�Ba~"7��]l���N-^�{���P:�qI�Qn��r.jX�%j�qe�.�pA��>�dEz�'�[�W��yĕ��s�Z�hk��熫3_���[�I(�S>�B�)��8�U�(m�~�C�10����a���!���LD��C�z�yu�����*�|�'���������T挠��������2wn�y���`��՗�x����t�_�Vc���T�碠��e�ԍ�M�g$Eꉦ�҃�G$}R����W>B�c�"�c�<�d�B�b�)���̍�7��J�]+L;����U��'��vR=8y��YC�}$q�3���
}&\s$}Z9��*8�g=�L',_�^?�q���&�-�q
�q�XC����}��C�"��pl�
�r�qD�o�̈�� 7��듛�x��� ��$�P`�����-�\O ���E�#�+����N���i-��$ҙ�h�8gÝ�'�N�}�;����H;|;�>%xjlrA��_�J^Ib9��f���<���.�PYO�h5ϡ���U͋ ��4YF�>�'Zzu��	i4��_je�{Le���}��N��y4��I6�*H>@U��r�6��X*�qn�m�5F�'O(�����Xs�K�7C�����V���3d��z�e���P(�A��_��ļҖ�2m�.Ӆ7ڷ9;�G�_K��C��Ĝ�-�zj�� ٰ��3�{��K/ ��r��Y�e�}N�G*;�|wT���,a.�05($�N�р��ԧv��K}��j�� 8�Q}dZW��a�<��%ŶR�qNg�"�D\�(�,E״3��ۑ�L�˟.5����ws@�ُ�z'P�n�h��e�g��s�N�Q9]C�+��VfC�0W�ƪ�ЌB�9�ʞ!�֞�A?���Sg9�T�\U'��9IP� �M�%��{��̫?ħFlݽ*���^��,���v�;��}eY��Y�K;�r��b�Ƒ�\aXE��և��R�>(��F�g�
��=}B��Z����
��5�ġ��	~Z�,�u�R� �C+��:��TM��i%=��=���W����t��H�}d��,e9�d��M��3�(�zE�A8��CC��N����|k)���p�>R<�vł���Ww�%rfњ/K��fB�%�=8[_"!�o]"�G�_���V�����.�a��ׁ�=Q�8 Vvs[� �;�(����[�	_>~f�>�l]�}d�Bb묜"w�lM�����B���2g2�=�#/�P�v������Y��c!Ru�o�$O�)�%�f��5I�9���{J�-V�$k��c ڤ<�����������e��迾)��)��W���hx�w������.'Vu��d[]F�_�z�ㅾ��gH1�*��rex�RX�lq�X�����s!��|�P�I����eBbqך�����BK����/�9���e�1�gB��a�}��Q�-�����!��~v'~+*�%$phű�Bj�.-��al�N�r�V~��
�L0��R�M���b�(����C�4H6�i��V�7 �k]��NO�C(�
�Ԁ�F4��@00��ƕ�qB��/c{��+��L�����B���TӒ"��]�$i�Y�����z!�<9QeW�',�;���'
�|�w	�{�}2HH�g<өm�$��ٮ�='�0Q�	��9��H�i]n��d{�EMeP;l��M;ULZ���)x��%��YyW+�[�'��-��f��8�t!�.�ge4ڤ|�y�Ȥ����{���4�Oph�|~���QiA��L���ˌy���RU�Bͨ2�lҏ,�?����bQ(?�u����lنkS�t�1*���5v�T� 󌗆�h
�ZtȱɆ^'�*٭�x��{���K�m0��*P(՞��kЛ
��'}ӂӐ̈́��w�+-���6��Œ'��ѣč
B�q�ʅg��p�}�P"d�؜��앇'Ȟ�ió`,�^ޜ�A8�ޖ�y�D�	w�_�0���nب6]ƺ��S�F���2#�d�O[��%�ј,l2!����q����"�NҢ���-ຸ_��B���kl;�/WU�\�}OUK�YMӜ��s8�/�Qh��
���	8�+��~k6�`/��"𞝁h���,u!m��r�d�=��iT��W	��/d���A�����#�V�d6RlB7M��"�2v����J��:��c��J��@]�$�j�3��%��;,rsm������-�{=-�Ů����+;��U��DJ3ݘ�p!㳝u�	Osfh�ف?�Dh�K��̥�k��BC�ؒz�1�kBԪ��G!�+�oJ�L�4Zw���&K���yWl����A�M���V�YS"�{dU��7"/=��"��	vE�ڹ�眰��x�ex�),(	�WV,���gB�=��Vo��F�������_v&f :84v:hi����Ǩ4�89�y�[Ƚ�������*Z�槧�Q��E��u�|���ve�K����R���~�NC6_���Ү���;$���Z�A�+������޶1�j;D
�a��=6�<�Хi�	�j��AlH�Zj1�F7�qs�;k���~�|�%�o��v~��A2�r��V]y$kW���r�b�k]�k�RƊ��{R��"���N^\�ܽ�Q��3B6�.!��@�;��
�f�_f���W��H��~�� ���!�/�[���}���:��z�2���&����ŀ�2$'A�7?����6R�$�le�R�$��Ox(x!g�-��tK�
���T�#Q�E�B�C�q�[j�V��	II-T��f�a�U=�r��x^�\r��N8R�zԚf�����v܆�*���h駲�T_c���q�,�e�
��ywT�v��/�&�5|�%��O�\H�����U�/T_���'%��*u���pMf��I��S��!!�re$uv�^�"��\��e�(��AS��5H�Gp8��M�	x����`��_v��r2�y��m��)����qo�훂8����,����~�[�x��<�kW]kXb�X�p�}0�΄pT��\s$�{�r���t�h��2|���wMkT���*��N��7�����j��O�2�w~�Ry4�y�=�
7�����OX�*6șo���zg�[�z?J��^�;�
����W���x����:}+���cL �1/���AB 6Z�]�o,�)F�L5G����Ĵ�eićY���RQ�a����C�&$�3b�7�Ko��勈��`�ź�P�Bin��f�
Q^������+p0�X�� }D��i�1���˧��?�,/�#1�@���>u�1*S�����|�
Q>KͶFƅ{/�;T��p�*3���u�
쿿5V���j5���x��ʘ�w�U��6�bg��`��_�%&]���w3��M�ŧ,���?��L-��6hT:q�%�:<l3��k�.(�I�<�:p���QZW�z"a�Sf8�䇐��_�0�=^7���p�f^�o#�/s�΢K�lm��f��1�E���P����o�.A��2�{L��@<��a�	�D�H	_�.Tθ�e�*��3������.o-�	<{}���o��-L���S.�6Mqi�0�,]9��y����%EaY���#J�]�*b�:��pzQ~�̓�E�Az~��G�aFJ��7N����k�+ �+��,������?uI�]p�!c��� �o��~��/7���I;��q��ף��M�&�#\'A|�G:>�dܞ��"L�wHy���p�yI�{�m\0��*���nM]���T.O���}���꺜���	:L�/�����x�K"a}�zy�����r�#%)�Q��k���ʫ�5ti=�ӗ��ݑKx��t|���AZyR��kO-�{�E8���Zy��u=�61W~׮>����Ag\ĸ!�1���[�Sō�K�:zl�o�5�~<W9��¹_���=��{ϛ�����V?x��Q�U����UKCqc?#�9�%�F��%~��֐(5~���=��ﶝ��jv~Z<�.~�j���R/�]^
a!!rE��E��*���1��|���5�G���놔�灆�!w#��оi���{�LbE(�X1�a�j�Imcr֟f�<�H+�C��jf�\>)�I��cVq�q��̐f�|��%����u�Rx�a�4�J�q���(}�;�ES.�L�Q���s �:	T �vA�D5w��X-(�aQ�U&FS����(k.��Y�a�N2X�a�
�O�![���R����-%�lI��娇Q�B�Yy�˝ޫ�μ�cw}��������_U�?N��ݵ�-�qsu���.ѹ_��ҕP���	}�76t&k�|�J�Fo�_0A�$[�u�Q���g��0_(y�_�$wkm/�z��Vx0Y� �/8�d,��/֛�X�V�vg��^���}���ֹ{!C�ԛG�X��;�v�eV݀�@\�<�����V���&;WQƉ�@�_K�j��̓�zU
1>�
�Dke�,��>t�B�oM`��Zw��F�`�<���C 7FC��
ahr���{=�� �eB0�+앲~�����'݃��,���
˿e̪�<=��������X�	_�xG"�1���Þ��6[T�)��������{c6��;*�b��م?$��J��(tVK"_�(���~��.�,J��˳�ӂ���ߊ�(�830�i��p����QL<��{�?�6~{�ν���@h>���H[����(b��g�	ri{`�}!D�ļ��j�M��z:����hʨ);�V~~̻�������ڡ5��,.6N�N��Uh�n�.�r�7���N=��gi����C{��&Ći�mBx�8K|������A�M
�`��`�i!�{�(�'��w�A�{��"qM| � x���Y��&�(��4
�ct�i3^�3p�����~�ۍh������k\xlG���=R���w.0K?����e��{��kxl��z6!����_�|f��[�تn�n$?[O�Z<?˾b-ͨ6��f�H����}��jƤf�kl�G~�� �r�7vqM�I�D�;EL!x�{]�$[�D$�yk�ʰvf0N�+���a�\\,B�i��jn�e�W$F߾M��'��W��b���F@�Ѳ��:o�f	�;�yTi�M�����ܠgi��}媦���Or�vi+��{���8�+)�J`A�L���G�uk���)���/���
!
`�����21�7�\c�7���_�$�}����[�]b�[l��~ �&���Х�k�SF8�����F��զ�B�藧2��i'!k���ST�p��j(1�G�ݤ��g¹�"W@s��3���/[+��S'��q�f4�a�/������&m,��y"{����S7<|$X�c)�J
��\	h�3�b��oz���g؉4=�4�n�U��C�町�?SS��^�IO�b�3BF!�i�F~���zw��1�]⛁��W��C�G�J�_�b�NA4�apH���ˮ9��T�n/x�??��,H�Sh�ot�� �.䓵Jb�Cw��䴣��R��a�5��Q��B此�ґ��0V�>�ؠ�*��J&��%�1G��*��;W��)df��K>:n���U���n^Y�=�i�5�z���p�\y���<�^��V�v~s[�
�u���Z�/�G"0W�i���哥���PR���;��|���!f~��r�@�@5	��TVQ5U����9p8�Ⱦ-5��Φ1�������kem������y�c2}�c�I�g�T~�m%P��k?�nZ��L���}�Ne�i���P�&�	��m�'�s�БXd��!S� ��pl�e�
୉﨟NnQ��шޙb�?iJ�j�g��]�>��8�����A��t~���g Ǳ��n��h�xrsy���]��&��w+���H$�4)M�_�E$�mV��&�l�^!e��DE�׉��ku�U�e�zƭ�y*E��:k���0�Ә-p�j��P�q�����0��tBp�����'�F\�^�
,l��qR'1��$���Y}}������4�qd�y^��jI�y|�{��ki<D�܁�x+D��>��KRN4�����E*AM76a�V�0��'�qK�lA]������uK���|r?���Ϊ�ߧ��n�{�qF�������8K�*���zY_�4Y�O3)9q��B, ٭eLI� �=!�>E�[o�᳧����6���X�W�,'��*�*�����`H.��ii�ҭ�av'~v�� ������%�����fti�엯S��7��X�2�>��'Po����,�NfUƞ��	gLn*[oK\�|\N��@�L�	�+OO�Q�r,��\W?�,I-��`H�߫���_Ffx�hV�&�z���$��(�����}��s�H��/�7�:��5[)����£��/J9[Jb�4G�\=���W:���
]�ǁ�µFt3��s��h��'S���uz�� |i��=)�UkƯ�_�E���+���Kv�y������z{�m�%	�6eaa��e�����->��=B�o/.c��Ot2 ^cKe��J���ГC�#��?B7�~�>�w����{��x.�^��,(Z�|�����8��EPd=����
���!�jG?$!v����.RH\�"f�n�B�-�rysN��������13<Hو] �h*S�bk����0G�ˎ{���%v(�`=C&n�oiE�tO�p��'s/u�ִ�K0rlq��+��"�&ٕ;G�#(�C��&g�z��׾�V��>ꖦ$�2{��|����;�TV��Z6Ft�SUs�U�5�N�~x��\լ-Y��x
�oi��</^G�ԞIE 4~S#,X�K4���9bX��l������� d����?h*�v ��;�n����Ƒ�az���R�����)�ՀG"/�
�r$����LY�@w���p.���!j%� ���,���.{��ŜL�Vd��Ӆ+�X��2k�J�"HѴ1s�2�:���In���mR꿭PS��F�R��;i��s��h�1`�*%[$"G�ɮ�c=Oco.!a�v0c�\ޭj��f�CB�=�����s�>�]����i�B��tw���~�na�}�I����4*;�k*Y�a"U��;�d M(����a`)�z���&'��(�Պ? ��O�����-xL@{�WG�-��5PFL�%�s
^?���+�$���7���K�K�X�������lZ���.�`Y��i�q6d<����,��@:���GW��_0����9ڂwK��Z'Wb_$`ܤ���R��ڥ��J�䥼G��2����������s���[�E�JGS}���V4Uf�=�������JC�@�C<(S�d|����;��n�D_�?O|8�Jv�!I�s#��f�ZY ]�k[��~64.d�'V9:��UeV���"E��|p}�\�ڸ���<eYO.T��<�[N�������$�I�l
+E}�xs���Ցw?r��靮z�)���N��²d�KF��+[=!�X�=s����Z����z�/���)�K�1�rC|_�E�S���D���tw�l�NMG#�|6���<��]9�{�D��c�|ce�<U��e,4�bL;��,�h����=:Os�5�U����S!�wBNU=�Jo;z���ԩ}��2�����-����)%��m2n*�E�2jGmx��QW���l6�u��S5�KVF�
8��1Sg�+��=L����	_�':���jS��̧"���Z����%�OT��$�1V���Q�mx��4�:�Vso>kD{��V�t/�q�uu���Ϥ����w��</��Y�|�ܦ����&��ֲ�p����x���p��o�E���?kf��������w�OW����-^�<�MD�.���^K�<�SM��lԊ���*����=y{��{!��y�VqW�$U
d
��L�Zq{�T���A"W��%�o�y�T6��T��n�p��V��q�%/��98���ѐ&��<�z*{�iZݱ�U����n�1o&L�;Bt���/L1TAo, �1�w���fwj���(�V	�[fϙ���ˆƟۖ �"���_���ui~n�5~"N����4��p�K�&7����g9m���og�2���d�b����˪�v�Y�KǇ�彚#��-��d5�]���|��-�X�hfH+�j���B��ݡb�������]��{O'����/��M���`.г̃���5���4���J�v~-��W�!������:��b�0y��" r��
�K��2:���8pW�4_�H����t�S��7&fd�p}�( �V}P\H�{!�a^LO$��������!|�;t-;���g;/�C�:�%��w��u-L	;��ܾzwL�[2ٍF�Zb��9��&�4��Gڑ�)�lِa��ֵC���ꅣ�U�p�e��9����#ְ:��ZK�g7e��m����6Du>|i�9c�?Eߜ柮��
��LL:D�T��HDP��h�I��F��Np_�� �� 9�o�������1�:��~�P`��u�bL�.�1Q���ΐм�xi`tQ��,xv��k����[v�Uװ��>���V!<I�<�X�͒����N�u�MCx���nG̊1��Y��������s-9vAeK��qS�$.�&by��h���d����+�~Q���m�p��Dv�.�2T^'�����c_;¤;J{��ʭ1�x�Z���ӵ�)��!$��V^��$W+J��h��l�陠"�O�Q�sG_�u���	{c�j�,9H���d��~��Ho����:q����3?�����{��(���7p�#%���c�|.Cg:�s��D��ewq�D��Ю�<r��E]5��i�9��.T�R̈́AJ���˴��:7@$#z��bA�g���m�u�a#Gd�sA�n§vϤ��<�)��>��������+�Gv���0�(*xQzX�~���J�e�p�����	�d.cF��<{W���ۍ@c�_T������6PK#�8�¤���k�=9��o�W�<��;A�Ї��6��_���?�W.�$h�>x�b$��7t6���ӳU$����̣�	I&d���9@��=S�:{jqB?�~�O4'̻�T{��g��Q�;DYOz��B������kHi�ڄ%ׂN6�Є#l��<֯2֕A�M)��[WJ���{�W�x�uO�{�C	���= �c��W?_�8[2����O�!ySoM�
r=T�b�Y!.��N�֭��S4�9J�C��
hp��J]��+�K#�u6�#�Й���
��*��d��]�߭�tj��~k9)�A��X�7�c��їn�.��,��g�19^b�{�r��!?������x��z��)={m�Ȼ����0��k勼K|���>%p�1�.n4����������r���|gA-�R"G�F��Vrv3J7<�L���Q�
(f��62�s2�1��o��~�{L��q+6p�x6aw��_�̎ n�cfϿ� jQK0�*~/���[w/O��8��b��A�	�Ȭ�3���=��ۓ�Zn�/ -=��Nc���g�i邚kN��|g#�<�/����&˂�>���Y�$�s+j2s�52nxK�~�yM�^�O=�aæ%!�ݹ�@�i�;�F� moM�ã� ���'4��5��i�BhX��ҝ-	Z�KR("�S+�':L[�\�N�s[ﰩhU(��3�u�F>o��� �)G~�
�ﵞb��m�XՎP[&���"qF� w��23��C�=�B�����ׇ Yr���M�:;�qs�^3��-|ɢ�p�[��|h0�۰˞�p C�#����u��@�g�7O�ɫ��d[C�3����f0%�R���#gG�.��O$�ī]��s'@� cq}����l�Ǯ��0vz��8Nv[���J<l���):�H�Rt�q��~N휫�&���,Km�*t���x+7�����T=����+a�g���V�K%3��t��+L�����o�(4z��lW�=��M�W�>����h�)�W�b��S
��Zm��QJB,v��Ԉ��ƈ��hT~�f�}�0@�0`u�!��I��A�E�C��U?+�F��v�GY-r���ߵn���Y���)s]<u/8�������Λ��N/� ��50�|r�5��ǡᎪ{{�v.�q��)U92]�x�� �1�D{�Ut�Z��]$
8A*8�b����.�E����K���8���ӹ�|Db,���1kn�ڭ>�����Vu��ܸ�<����7���D��4ҭl��[
q�~(��E;��ר϶��a�E��$3'2������L"U
�~��Fg�iE���og�ě�s4�+�an�!Hj(*���]�.�88F���UN��D|ǈ%EMYў�{���;����ӕ�|�{e$iW�q�+��9;�RI��U�!�;�V=�K"o~�3��K6+YN���S��jk�m>&�"���-��N5P���;R3���:Y�	P&"ѡ����^ÿt��-�w�4&�����ߏ?�j��RcA�3`�:J���$Z��'.�>�+g�.O���y�ڃjG��Eg����'^qUc�j6W�ʄc��f�L@�?6Tc�?jQ@H��!�V�q�Z;�}�R�@��uXSj�d+Y.4�	���ۈ�@�eΕWb*��
�-�H�5�.i�z+d�cm��#�6Y��f 7j$0��lGڭ��q�f�BW{ͮ�2%�V~C8S�Ʃ�υ������1u��5��|�q�������y����$ƐݸH�q�<�L{�Mʳj�N 3T���\��~�7L*�B�C�2NӲ�4r���;]�TX%W(�x}�Q�,(<��p��V��w,�?��!�GWœ;���o�@-" ��cV���lG��T�@���,�V%v0Ě}4�����[�ﵼ�hɺ%�J&u��?H�x�Mj_����VS��
~��_�|tK@��M�~��d3��p0��T��`��rh������n�����z�����fC�u=�
%����H�BI-k�juT"JK��D��7f�}���!b�P\���ׂ��i��1�bi�Gb0(=�2g$��l������M:���|)�&��C�/��
*��/�Yx�`�S�^��A±�|0e.;
�J����h�e	�*��ݢ���أT���I\���e7Gr�	~)�V��_ԅ�-�5����D�U�/C�:�_Ƣ�~���q�$֚�K���g�E�U��k���[y�!'4�-̛��L�@3�Qy/s������9�̃���z��4�O�X�������`si1�ir�Dށ�y]���U�o��؆�x4,B
��z8����6���Dm����&�E�,�M��2��r6��ٸ�!��R�.(���*x���p��%�hj�%�K��M<��X��gk���@��2�ҧ�-v6�R���ma�b�婲�m=y��9��k���m�Z^3����3���Bp:�z���A�A��s9��j��3]��H~T4&ZW�Q]|n�L��������|�'>(@���^�>�	M�f�\.x-{���>�S�3���j�e�d�{�M�f����`#�� <h����(�N��9i��@c�U�6G�,�A�^�L	�m5�[�@z�F�?!炭5d�HA�dXD5g�`�\6��41�>~�����Щ���~��..`���o�X�w�Bݾz��<AS��������'Ec���!Cݪ��Q%Q�,��\�C$����,�2xf�M��((5y�T��K��Y�^�O�$�C��ڕ���뫸0N��	Λ��垭[��T�|"�G�r�PS;j'���Ù�s}T��IGZ���K�_�R=$F��8y���2����x���$������ iS�3�5��,zᒪ�#2��Q��Z[u�t�L��-���y����n�x��٩�T���o����_��b`�Ǭ����V�8����Na��A�|�Z�9
=�iZ��a���J���q]c����5��X���p2Y9��9 |�a�P��=�����`"`�!��E6��������eq[�t�0r�ΘE�B��0���p�In�b?� X�j�H�Vi[@/H����3{�C,z�B'���i�*p1֚����|�ݒ)mA~>{��h��LW3sʗ�
�<
&�~�<w�;���;Rׅ�$�t}M!�^��yi�_V�R��z<E~�0��v;���b��	J�����̔�to24!{��Y��@�}'���E��^M��'�v)��j� �]@����sBI8Ym�J�P�'��̎/S�uF��c���ư���9Rs/�k�1�}�dqi��j�D(挊�gWB3%�ц�������A4���O!�R���T���������D��H���?�^�in�s����2����PW(���]��'?`�/M������Ke���T��P��]��Y��+�U���+�[���x��=Q�F�x�0䗝���>fR�МY�BI���¸�$���\4꺦^n\��ЂG"tH�(�.��O���G֫�R����="E9*�H6�S�H��XS���L� x+�c+_���V���(��q0��׳Q7.ov樅g��hJ�ԇ[ ����ʡ���r$fG����/��o"����6�^���$t�%�$�H��/���CWôDs�"|8EZ�=��Y��É�z�zᑩ��=��+^���S\���^��S��/�+��?0�Ϸn'�fܒؾ�b�$ı�P�w�-���������#J������Hz�R̓:ZQ.>$���c�}QX�4�8Ҡ:Y���a��A�`�=��#�n�zFC»��uhV��rQ�!2��M��Eڎ~&�6s�u��Z�p\8T��:%�C5-Q�Q+���#w�˙o��\
\��:w�t�_�e�~o��<�I��y�z�M9a代�5L�� ��������~��Z�M�D�jb�2cSy\=�5~Ͽ���YwdLC�IlUI�_&��Վ�=wQ����E9�3�Vq����)q�pFIеQ�*������?`��^�r1�h�E������r4FrD\�%+�.�1.���rv-W�?��i(�<����y���'����e}��!O#ϵ~�)]�f!C����8Aҁ��چ�WSHu�T<'��|�}�1�����p87�څ�-�y��=]h�L�7��|~Ҡ؎�k�T��i�"���Y�[�w~��|e�(�eOZ���%��O��Cqc�䂯_~�10�Z?����b��K�'��_^7��n(l��W�k��[</Q��:=s���O̜��\�P4�]	��7��XHh�2u�7�v����k��?�}�W�O�m�/�H)ŝ�P�J�[q�	�
T���
.mqw�"�i	���޻���g=k>̇Yk���{���̠��vg4<���.Rc�2���eP���T�_e�����Ԭ�ָ��]�Y �3?���	�5Q{�7�<W��c� l�w�|p^�`�O;�K�]hl�bX�T�ow�3䬽�f`�mb�n����"�ߋ469�+��T-�X�ݵ�I7�졢���k���]��K
|2�b��Δ��2eX>�·�<}F�ҨS�,�(`�ꠀ\� ��bi�����!y._O�]X8��Ca��HD�t�C�l���K�
ؑ�Ș�<c2�}l��yu��3m�8��� 
�!p��r�^Sz̄�L7��4X��(gz*�Oqt����18&��~�����5Ce�eXeu�}0�J���7\�lu�_��C����[�ŭlj�]���ږIl!B�ځ��Ed�N�a�,g�4R5E�������x�ڻg��!���m������E������e���kv"q4�`g2�O �zx|�z�3G,m�A�����NQXG���V?�,�(W�f_KA�BQ[�}��t��N���c���7!��L+P�|�hU�H0�?
�}Cx|-�4�?�5��k����ְ��aw���<I��~v�:�4=��X�wf���k'�G�$t��'ǹ�v/��rۛ~e�����5��B��Ei�`�H�Ϳ�]gKC�p����~��0�7��ۿ�k�㚺K�ݪ���Nꋯ�$��]w1����o�R#7��炶=�d�y#j�^sl�k��&ؼnv@Ke�k�p#3�7%���O�#��R�퉞���Em.(���{�jW���h�CﬂS؏�,�.���*1Y�.��AuPށ�ך6��7�(��1����WbW`ǉ\��3�y�)�5�s̬�0���y��m�J*� ��<��A���^�5�t�I����)�|i/;r�,j��W�璦�����t�ӭY���l�<�u�cd��ቲ�qj�K���� :�����n�p�g��Wq�tD	CaB�	��c�\�b�$�fI&��B�����Ox�gS�ݬ�٘y;��Ȳȹ�r\�A�=���OpN�5���|ժ����8��aVq�G����kVd��5��:"�1_�
�����6��Vz>�]W��il�u�ӅKhc�8�x� ��*���������sD8-Ue�	�܌;�s���-��9�V���q �a�����X?q�H�$\�BG2(()�^Ӟ������A�N�GO��YI��ԓB��%3iR~6�k�|{�#k���uZ.^�k.N	!��~�.��;��|��V���PN1�Su�8'N,���P�@we�_R�Y���҇�u��%��٪z���0��g�?\K����u8�W��_M%���a�^�%��1l����̚N�:�E"L�������Y�v�Ҟ�d˸���YX�0�s��7.- �.+=�"ہwƬXs�{?����5��!��D����P��"�a���A�v��F��"�gi��ɝV�ո��|�ה��������T��6�Xc��翋���2��1,֛,��䋚8*�uC�&\�9<<,d�]h뎫S� כc���*���G���E�h~�\����=���6�]��h+>}���'U�]u*2m;�Z�`i"�]��A�3
������,��Cv�Z,^��ț��oksn�g�џ?z��K�l]��5��R3C��9K{9i���(���;f�$���(!���
I���7bJj����dS����e��Q��^���\RMk�C��j�m@����f��,'l�[���쎗��7��q;L�Xʄ�W9��hq�e`~%�����ˬ;S+��ֱ^w��j.��w�4=(�C#�'I�rC'���X6��i��I�W�P���Ls��pRm�t�MVi�<��)ʣ�RH�Ȁ��
��%}N�Z
����v]��W�A+��:���߬Uwm��S)�����E��[�셨�P�¯�o �i�ᎄ�0���j^&;iH>c(�{�PEf�T�������/�q���� ��(s�Ԡ3���>��~�)YNbg�UvΚk���B�E'�J����?jsl�	�ur�5a�oPF!@��2k�p��S�H�JŦ�Ҁ�(ݺI�u]����ml��ʎ�I7�Zx������GCK�Lv��9?CR0LK2�I�E�� l<��lnm-j��~��f���-�Qbwf"�L�e��B�Ύ7�/H<x��ן�����xF�-�������(l�e�v�Ӱ�A
�n���٪� ��\f�K1�p��:3�d���JZʠ&����y�&'e��HPB�W}0:׈�c�~�y:���K��Pr��V�`Rv��Z ��Q�hﵓ���Ag6��Y�6#�m�sjC73�~��ش_� �8�)?������.g�Fr�9i}6d({Q�{׬�H�{�)ut�0?@�w�\�#z����ƺ����D�.<��%y���ΊM�W
/�����5%Aw�NQ��/4��XaA����U��RD^�zKǘ?F�k��OǃZ�O�tT�KvGE���`��K����]rC�ǥ���'@�->�1q��!����P��1jb U��������\���G��4�.��s:|�[/��I<��8F�#�wa��Uy���X�$-K.=�lw����a�v��r.���i��Wm:=�1��:�?KF��+o���i�9����&�5:/#.B�Dc+o�u
#5�C���5�����JF~��]�����{���)×q�\�dE�?h��� ���v��h�^�6�L�
Bܶī��^��9^���9:�f��Y5f
��X�c)��K��:���k��2��.��uOT�!d��g����կ���}�Rk��4���e%kv�o6]�	�x�;�\�?P�&��V��u:�!�oocofz�+�܈�e���^���6�YA�D��� t�]T[G�q��>�vi�`oT�
��b���lR�.ۂ|��Q�$�>i~{M��Ȁ,{8���ӯZ�a�H��h u���Xj�+�������s<s;�]K��/[>�ӠǍ�2��JW�!Y5�5����V-�r8��?_���޲$#�w���Ju�;1������ [���r� Q��K�z�ho���QӰ����*m�$9��t�9%���1t�#/V�;�wL�Qfy�,(|ςU5�*~�~o��m�9�4�"D7~x2�3��K-��~eɈi�@�2�?�λxDUN�h���^_�9��T��B���@W{RϿ9O%��3��o�6���Õ*�`\kF����.+�ո�\�O��ͮӌ�we�7��\�f��#JN�$�Y�mI���g�7�W�`��r�=�^�sWS�)��F� 2�ȇ��'w��JeC��t�"���Fq�n�Y�Я
p5?&��'���D�#U�|W�/���d�0so$P�����{b���5�v�;�[|�#Ι�ڄ9Fh�u���3!��Y��is��_:�bo5G�y�Ʈ�d�ã��$��j�	�!�ǆ ^m ��++1��@��R'�<��_�Ä�~�؋�e��v6t2pl���\4Vd��Rʆus�nј$�pN{���߅��5+,�F�I�1�b(bYϘ	�;�VG/�]�n�y�=�d\f�ߝW)]��)/��b�v\;���Z}ҍlƕ�.$.�ҷj�\����Y�l�:Kc�p��Ap��E��/̰LHyI'{�F:����Ʌ�"��$���GcX񷒄����ai7J�����1�U-�f��5+Yr�RX�.'�-��^��� ����a����#s�.��dc��!�CD�,dC��c�����k!���QNxJ�Nx���|���ieh��K����Ă�;SO�0O�'�BɎ�X9�Ө�E�����Kc�΂�e���]��|��1(�'Q�y?[&$��������E��٭Ͽ�#䴳�i��_w�<���p)��b}V�Rx#�������{�u��(���為�B�(�� ����hq�&��Y�+F��:{��)�[��yS�l۬��)�Rl~Q�1L���ѱ8x�.D
��W��W�Q�ڨ0k��Ag��ݐlp�4�pq��3O��1�Jpv��$d[�J��˩I�jx�L�[�M6��d<�y��<�K��F���pa��	a��OGl�v/4Ϧ����2���q0O��H��6�6���d�Zȟo��"�%�ѿ�=�o�Y[A	�BV?���X�B~�@�W�&�� ����p�)`��s������K��7��	���T��4���kw=?,�t
,�Ia9ב1niN:%A�ڟ�i���W���i���d �ߐt��A���nmcL>T֫�;\��A�'u�C�"�tR�߷KpG�$�2ٱ@�]�	�� �^3�x��^\16���w��F�4�@�o�fF�f�;?H{�x#��\�N�&~A�	�3ne�I4.n8�22������T~����B�n|�<�-Ć���V�h��k(H>���1��Aax*/�4� `d�޲�T7[��Y�uX��ـ��\ѓ� �H�UP���6��*Ǽ�>(��N�V^�������������+���qfv,�}�iRp���,��鿁k�f�/��b��SǬ;i7u����KI���ʝ��KD��2�(�H���U�s�y�S�bqC�����x���ʖ\-���[+���|�c����ߓBdiS��<����Әa�6����htN@^L�h��p��u�hU���P(�ޓ=�UDO,aVw���aւ�P�8T�����W���	�
Y fX8�`5T�iL%o�EOк(<�OaG@R�X׶�賐��S�'	�!��z��f��l�g4�Q��ء�l�,g�<%3o߼�3(�.kg�!��w�M�XbQ��9 
\��i�{��Z��x�ht_�g�͵�9��7��1ͮ�RW�!�{�њ���n���C��<�^h�jM�,��]-������^�mR�G���v�����N�۵����{]`��h�ݲ��E����I���>�bEݻ��|��s]�)��\O���6ӳ�,h���뛃"r�7)���vi�'�غ[爻_�]z��U@s�ĉ��T-~akx�����\r��Ty9�˲��
�*��m�Pnu�"�O\ޡ�c���7=�5���儈��b%�W)�@g<%Ob�Ƅ�fP��V��:���)��v�P�=eɢ˂��Q����ͬ�v��R�[&��v��Yǣa_7<�WT������+5������.f�ox%��V�>T���gKm��o�`˲�:��_��:؄t�� j+,J���$o��ɴ�RrY��ɚZ`�/@eS���x��%$Ds��]J���	�����&Q����������)b��i�h(>�:iV�}8[���_#�����v)�1,���'�����{J��lLS��9�d��O������$�s�g�y�cT����I	��|	l�1���&/6a>�m�SW:��?����
���*�k�-U�?'|Lٸ˾�pEO���5���L�M�A��r�C���s�E	H�<s�`� l�1��R������
O*ƈٞ�p�����N%�Ur6��7R���U���7�l��C�N�#� ���BL��:&�|r�-�.0_��|��U'm/2,6���C��Ǽ��EeHe+C��$lp	���6t
����Q��4}� /4r��'��DĄV��&�퉮!4۬����E.���Z�_E6���o���ݮ
W'' 9ha�)��,
N���>�� �3~֛���dŵl�L���Y0f"F3��xk���<q;#m����Ȫ ~�a+E�'b���F���oX8�X}��"�<_|V��9�Y2by��]w�V�L�ǾJ�	wL���ګ�yJx;�x�5�;.�`ģ��ֱ���� ���)W�MN����~���2�	���.<��E�7�@�}�h�F�n����;�"����A�� �6N���m�����v��$��w'm�O��Z}m7&�R�6����l�@�'۲
A4�^2��1�<�Fc	)�\&�{y�(��M
n.քG<Ǜ��d
�����T�?6�A_�/�8�j�����θ�Y�n;�M3l*���o�0ìy��E���'��8E�AyT}u����aَ	��U�/L�a����q�p@�����%�d8�K��6�pZjg������C��X1���lq^jqK0�ne��
��o���E١��Pȝ��;�����:��x���:T`!X��s��k���#���2�D]����D'��r�SAO�]��obU�{N��o���OO	�'H�!�u�L�m5m�IC�,R���O�I�g�i�w�Yr�B�qG���N�p�0������O�'?'�7?��ё���n~�'�S�+�rK��m1ӵ�m&�w���$]n�����[p��$��g�!]�Yf-d�qw<{7?ZA��#��F���O7�n�M2�I�����/����lc��~'� "1X�CM��ӷ��d���>H��ۑ�}M�}��U�P�q�m��, .�&Ɗ�s˞�a�r��G�js��(�hȦK�f@zل-�@�@�U��el>��?:�v(�&�G0Q u�Ҧe�[ 1�^�#�!`BK�d��p�~A��}a��Wd��c�����<j����R�]�o!�vWB��'N.ӧOP/���p���W&*�t1ގ,�PWއ�L�)&���.<���6O��SG'�'�ݘ���hBpx	�m�[��=��B�f���%� %Ӻ"�0F24�b��O��[f��	\�
�Z��I��*����j�*����XE�/�tc������|����cڜJ�..AFl� ,!RUf�'}�d�Jg�9���>�3� }��:�-3ܶ�+���3S��l���SX'�?��)dR�f��hS��:��}s�O�	����|=t��uu���3��OC�5W���������
���|��<y:=vf�4و�S�/U��kz�\��+*��s����r��޷e��g���ț;�X�
%�	�F�{O��A�z���FZ�R�Zʱi/���y�C��<V��V�s�j�ؖ��v�X�fy�L��4�Rz��1�� �=mt*4�����{��K���BAW���_�+�mޝ��s^�zU���b1e3E��.��� �5�ʈ�nYw]C��W=�yW�Υ�u_�Ŕ6+~�+|�}���ۀ`R�������\z!�@��#�Z�	O��ٝrB8�O��a��A5�=�b=�.x�u������u&=c�w	h\�I摮MC�{���d��w�Y��wz�>uX���r)�����P��il2���drn���:�ٓ<�a�[�ݘ���H��n¥,�q[z��N�Q*��d'��FB6���1��r7<�aک�u��\S����Pe���R�N}��NO��t���o�G�y�n�L2�'�\������0z>��xo,t��@hD�*EZo����p8��R=O��`�Q��he�������p;���$ѯTf*��bd��h�2,;��s�iv���m�@��� ��|��Pd�XeL@������%d[�P��$m��{��s��Y4t��P͔��f�)�3��A�9�R�t<;�����z�O���F��]��s����B�4���D�H1��pk����I߂ԫq��P��x�-���Ca����W>%��^���U���X(H�c]��I����g鯃�����J�`�U=����x�����׶ޛ��_ᓑ���f����5fR�A�R���%�k�Oߺx��@�yfNƨ��	�&dc��`7�hc����H�*L�?�B��d��y���L��f3�4�;ۻ���}v\k~ʽ�!o�����ϡiۼ��IEurLô�y"��Q��ev9� l�m��L�V.����W\� �k�ơ�5���h���Y��\��B�r��̡�2Yg+Ps��2����OԜ@v�Ŧ?�q>:d�n�;�#�,&6d\$h�����q![�ҙĤ2|^rcpC��.yf+�=uP>��6f)�O=˔P�ᢣ�e�Ұ���[y:y#�5��l�4��ȆE��@9G�9��>B	&��g��xW*0�_�6�9�!���&�\������"I��p:�kXLY�9�nX�׌�T����1&�V��f�0�����(g�~Yh\-� uR�Q��O�l����0���%�~o����ֻ�û���h�4a���½����ɡ?s���Jڜ�O��/�Y�MD��b!C+C���X����v�{H��{���/�>s�)����>Q��,`�	�i��kS�L��.���/s	S��bB^��Nc����T:R�2��|f����s����%.q�͝�AE�۽���O7ݳ)��o�����q�O�]����xlXÒ�b���ވ��!�J�0Ǌ�u[�rj`Ed��R���YX��3����������ye�x�KVr�o\��1/�a�e�C=S�()3�>�7���\�{��'aL�>��[��!����_F���̃���~��M�NY�ڲ(Uzo:�f��cv-��������3���$v��a@ɲvy�[
�Qa�EͲ���Vܴs䕁}�m��Q@�J�QF��ߢ����J>��F�sj����B��[�Kr�ʥEeɦ��mMo��ֹhwy|b?�@��V(�Ko�`�4���uF�M������	˴�w~~鴥����V�%3���/�>�{x��9,u��q��]�"6�G�I�'ڗ�R�L�}����fJ�Jژ�n��&��yh�{��� �N� z|�5���W-���ug	(��d�;
��qq�6���R@�AQ������\�:�	���ĘH��f�U+�y��(\n���KwW^��N~���l�-ѿIW�����;��Qfim�/�5pk�����֠�*��n�c��c�,\l��K����.j���U��T�B62�+��OR�_���'zҊ"�My��u��H= t���|:'֜_7�t[�U~��,T�yQ7G���)�>����8)a3]WW��fR(؏�kH�6�Κ��5
����P�8<�0�9�o��Ŋhd�iQ�2#	ӸVҜ��Gd���Y�/�$��xw������_�����[���R����y�0��"Ƭ�]�S�p3¯fu<%料HA��a$����G����u��]N�����U�a���]\��Z�Wg�UAD�Ca*���3�t�ᕶ4��=S7+ᒅXs�(��4Ƭ�}O@6O������"�J!�٘���*�ؠciz?.��\\�[%>Ux��\�{�Qjy��h���v��-2�.?|9uEO�
�����ܛ��Iqʭo0/D�
"16*�)
I/�M�E �9<fTg/��O��I� ��V�V�΢.X�c��G;����  ����X�׫gg�M�~���B�J=Gz�@%}���.z�* ���:��n,w\\0S�	�7��k��.�]���kd��>k���[l!{z�ز*���Rc]}�rK��33�L�f߿)�_,��
A��J5�v���aϹ���P���p��մ�in޶o��J[R�����1��Ǘ�ll�~��9��
9�6U���b���������y�������ݾ���B�d��e:7��Ƶ�0�|D뭳��P���i���_�r7��������y��V���� ��O��[t^�0�w�M��ݣ�_�wfN#xO��n�27�ě�Z�O���曚HQC�1k���[��T�B��[|����W��(�_<:TAP�P�M��χO�{pP�E�+�`�g^��5��Xi����F�����&[r��Ozd3�2uq0[l��E�NZ஛oVGr]RǾ��rw׻�yL������ܴ��ecqN�����*�U��\[%Dc�/x�a����U�K����΁��d���ߵL@�����
���Q]YX]�C7��-�$y*�b�P��E���.�k��P&����rl9Ѧ��}tb
	9��ڝ`���Z�-�9�p
�s�~<�a�/{��`��=����\�L˜�G�/.sXDY\
-��OK��ȌW*�wߛ��T�[zm}ei��k�����@�dB`���񔾁��8���Żu��XBg����q�f�:��96�'G�j����8��=�I��}迕�E�P*k��[E|�����1�uT5�h�l���|�y�$��K��ʵ�vX�J�o�l���r��7-%�gh�P��=J¡K�!`�<,�&2Ͷ�o��uȑ���J2E���X�,^	�7�߄�^u7�}}�W�c����!�w�����C,F�sL�eߧvr˷����0��?�.���$�1�l[��d��g	��'�F��*��3���7���>a<r�ۀ�gW˒�c�Z�n.�%�K�D�R��!72��ҁ���W9�aIg�r#.����y��ԡ� �}/���N���&��)ͺ܎O�o�e���pI�u��֢g7���,�J���	 ���	�O5�ɽz�/Z��_^����w�I��d���r�#�����Z�F��;�
�Z������tsj:nl-�ȇ^�<��L������w������ Jrxc�STߪ(�9���nx8͡fg�`8x_�Y
�>�fJ*�*5�?-��f�9�!I�J��0jw!�R���@0���ol�D��#E&ml�	�D+X:|���������zP<P�KԢe"7�i��)������Я��"��Pn���&v�Et._�$43���9ZXN�����;�h�|d��h,��Q�f�Ҙ����{3='"���zJT���UR��U�A���=<<�-�)��d���e/��i׎2����[�7S��7�aLx�(Cr�㈢k�u����L��n4K�б�(��n���'�"2����c3i#:;�6Q�����>`b�l�[1=Џ�����>ٙC���l��ѵ�NB]�J(X*���\�u� ��W�D�>?=�Vϗ��D��j@�i&��Ic�&ԭM�e�T��Lqz�L�etg�ƹڥg�Yhč�s���C|mӦp�/+���L�HspOQs��XaL$�W&)�Y�]6�n��!�m���5��T����]=,E�9��9~y�T{^<U-�>PN|������>���~4|���q"�M6���
�N��-x-ZcE?�*F���g�f?Rb���D?pN�@5���FV[�����oc����0W<z��!
{�2)b�s���yc��wq�*J���N��A?
#��]�E��9�]z����Հ�|�uD����>��8JbU��xo�����ou�B���M��ֈ�jdɎ�p���q_�λ�]��έYL����[_ݞ|9���pj5]dD	�:�,i"�t쐦����.l.���d��DOp���B�c�\��=GeE����'�[�C-�.������.C�DOڿ��O����Ǐ�Ӏi�t�z��?3��]��~M�:̅[L�V�&5��e�&�6������=�>T���a�}8�ٿO��w�u~5��`P�}�$PR��].d^����EP����u�W�bz��GO_����A��#7f���֝ԒՎ�8^|�*��'2|T\I[_� ���q"��[n�m�'@!_���Qݘ�b ,�a�Q���iz����@Y�Ýq���AJ�W �;�����	�������g�k8���G�Y�F9�J]n$<TXW[QY�GI�������`�G�?|mć�*�+�}@�)�exF����J3�P����*�����x�K���[��#���"�L�=�t>]C�*�U��^5Zz�%�l��k���#��Wq$��u�<�c������Ma��
�����v^��T����n�G����Q@ʶ�r
X9�INH�|bw7�]��7���Y����/�/���r�t�n�S�^�Ei~֜ISհ��5��H����4��ڒ���z8S�rS�dY��0��o����������ϑH��pD�{���rc[��+�̀�(Qo���Ju�1?TG>�h���'I�v��:}�}M�zxm��,�$7��x
��TDӊ[��̂�a>afgB_��4W�~�c��r�d��VT{�|e�WG�eI|�`l��d��Cׇ5��i�C���;,?I�]?�T����6_�K_=���7ɞ��4Q&���=�����������G��s��uJ��g%q�Ui�	���.�1�	#����8�U��{�XK��-z������G߆�ޝ�%G�#%���T�;I%�p+T�:%�u�C׻~D����A�����������J-oz����%��5j�}�quvh��3������4����*�%�����_�^hU�Є��cS��������NX�f�q��
0��qu�塡�������A&��X�Yd������<�������3����CW�ǂ�/�7�mA���6��x�
��e�"�Z�YjI��m�y[!Ԃ�r�qg M(r��#�t?�z��l֎��3���{a�j�O�c#%ӑ��(���z��i.�ߩ
=i/ BBB��<4�o ��԰�	�~�R_c�r�����z�n��*K� 4�l�S$>�I�"'�«ei�=h1WB�T���F�v�T(��)�����LI^��n�
�
�c:�Ҕ��:�R|��]��,fgrG�fi�;����煬������T3҈�r�����ӄ��k�­�u�F���C���r�6rT��/+$yA8�v(�{���]S��1���d�<�h]ML���;�{���uo�׮r}9F��H�o#����+�|>n������x%�i�����+_�h�t���o�E�T>�� c�#	�{�Pu�i�mYZH��<[�+��:n�a]�G}μ�֔��+*"����������$� ��K�f,�`��gF����*��0�%�u������,e�B;k_�T�FqMB7W��%�����G�� 9�Ռ8�=��g�dH!^�/[�JY�=�I��sO}:_q(�ڤK���<�Lv���
ܳ�9{v�#Q��������Ȁ	?�L-��K���3���Q�0m����ve��Ͳ v�##̳�!7�Z'��H��O#r��>������&���W�bLX�O1�X@-�R@Jj3$�4T붰 �Ϥ�{�Ϳ��m0|l��R�]e<+죦_ZC(�s�EF}S��xH����&�h5S��\�K	�{o��7�Bs���C%;>�
��z��Ϊ����%����mf��w�*�g�/��o����R}���uo���	
���y<�W����a2�N�j��T����J����Q� -�/��<�$^^��s��" ؗw椤�^0�Xi��7����3Q��b��߳��Y���u�}���9橑��F��b��:
���v`
�����r�$%�ꖾ�����;8�^p��Z0���Ej��j,�.���ؐ���Wv�~�4y9�򤉔)W����L�$Lnݣ?�����t������(���I�O��Ҏ&�|UM�����:Ӂ���(+���~�G^�'91=��E�y�>��n���լH��>��-@Z�������C�}ѹ��o�(��յ\��Z��	��Dz��c뽞�o��3 �f�n�J(��gY����D��t9�=�s7���U�Or�P��ψ�C��+a�ѝ�D
ף�t�w������P�\is��Xv.!��ʯ5^!^Z��PK   ���Xͧ��
 ܡ
 /   images/d1ea3d2e-b350-4687-bed1-c7e59b56e556.png @㿉PNG

   IHDR  y  �   _�]   sRGB ���   gAMA  ���a   	pHYs  �  ��+  ��IDATx^��`G׆��Kqw7��ݵ@-�N)�Kݽ_�[��R�%B�����=y�����P���w���ّ3�9#ۯ��W����K���Eh��i�/#��RSU�����@��;/���Vtuu�mss3J��x}�G�_����+�/d\JP]U���6tvt�:]�Z}E{�����"�w������GYI)��@I	��XSx��4���U�Ew�M��}ٿ����yb[G'Z���q�7A�[_ߨD��O��7m:�;�y�_7:���"���]��?���F~��҂�f�7��s�ҩWx�n�SZ� �N���Ikk;���xMq�{\N:X��������:���ʲ�Ԇ�V�A���'�E�[6E$��l�����+�����Ry��Рʻ:̭.^�?��"MM�L�������RѦK_�g~�^��Z��x�u��������\I[�[Z�x�������s�.'���K���� �#�_�꟯�wD{1����ԫ�t�Z��	}�R'mm,_�߲��^Z��F������(���ϓ}����l�����|�����F)*��Q]]���
+Um�F��mg.'�}YYYoy�$^��+ۢ�EG�$??_�)''G]O����)�{TWW�g�]��A��)Sm�-��tvj�L�D}C����~~���-�e�k[��s�G�k��?]���ꂴ��YW検��+�s]������"7-�����,���E足��S�ffTU�ONU��v0�"W�GR�D��y��J�n��+�W�s^ZF/���+Ϻ����:.�=����F�t߱�P[�wZ�v��c�����q�"�r/�5ӌE��O}fYD�$��C?�7�LR	�RHa��(�F[�"�J&���e�U�b�w���ה��E)+�@s���lm�FF�R B�c_������V���żES�ʡ)@nA���B��,��Ϛ�T�w�-,�r�>"eH���9�-�l~��v����嵕(*%��z�L����3]*
���rƭ�������󪽵H�����G���h�Nw�4`:ŢKWu~�7��ё�ijd�zB��l�nUXD���~g{3ڙ-��<��`D�:X�zD�.VRU�$�#��r���5��j%.�\nu�""�W���I'Q^�Ɖq�̕��s䔾"A�Q���������u�g_�0{/�Υ�@+���k��唗4&U/�
����+���o$�RʨN�Y�AG[���v*FT�i�� �H����U�$�s���}��en!����<��$\��/��?�A�M9�uK�Q�>�~O��J�s��MM�l��E��H����k�����OyF�.	r�rq�� ��5�� :�e_�3jJ���ummuo� ����D}Q�9nT9�
��z�� I^�u�>��Ҿ��������E���7�uϯ�YҲ�qI�����{��������꽯�yjjjT��Z����Wt�QD{�u�yKJ�=�ӥOAA^�h�.��y��i��E3����<d��VO�+�T��*�ڲ{�AΔ���A�/-��pI��܃A�j]M5��J�TY�����f /%)	�Fbf"�r��D4;�{ȓ85����6>�DSE���?i�YC�0h�`:s��6Z�Zay���}�4w7���I�V�a�MsҞϺ������NZ:[�����[��oo@Cg�%"w��5�W�V���
T4�������:4�����gqR4�T���FN�K-�JU��MUs9jy���jԶԣ���R���Z�4U����R����Wd��.��5���G[m9�x^Y3��^�'���?�~R u`U��JZ7����k��$[Z.���e�<��� ��;#;CU�\٦+)��(o���\K~+��ܨD�Yk��BJ�cċ4���R������$���+I�L齗Hz����*�Q���������Z(��(Mhh�E]#wmʫJ��?�y�8�f�!?�d�$ҲIAvj22�P^�!�U���-�5Jd��#���ڤ���������e+�������YW��z^��A5�͌����*��}��kFu�+QmL��J�v%:�딴��RԨcM,D��h�/S�r\��Z�~��Ԩ��_4ؗ�L:�k H������
���f"j�y$�Չ4R�d�S��c:�ϵ��N��	
2D9��[�v��ܳ��b��� Y�U��� ���� ��D�5�G�)��R��S�_��{�.��oXOE���:;{�([]����h㧓�
��^�����N/H�!�&�E�_>+Q��(���}�� �7�����$�dyF��2x��%���ʗ.>:�kh�n����A�#�Z�K?�h�M����=OD]�"�U&	�d�_�� i*�=�g��H��N�-'W )W틧.;/�Fw.�n1�s����"�G9_~�����_{���J^��y�6��Q1�Y��\S�Or/���MG+i�ĳ&p������8��A__ G���H>��Dt��b�cs�r- [Q]��]D�AI����HV��=T�����s�	��Ũ(.FIN.j�P�����4�@���'e@k$3~��WZ�%����K�?��j�cTS�����|�F�\^xr�c��mlh�cp**�!�hu���<ѱu5l����b���)�$CT���`|*����s�PV���R�:VW�<��DUQjK��ύ�Eh,/D=?�1m+��\��,P[����Sj�΋����+�4�=Y�k������AC>ǭ|.L��&)�	h-�Eca�rRQ�����ćC��¤p�&G�,6��ѨL�@yB����8�d��)-MٗJ[AZrS�~٦1=]ISF%M��%#	��<73Ȋ�c(��J�>��%>��	h&D^�̨�Z��Ҋr^����D, M�U��`���&ӡ)L@n^4�bN#2�B/Ĺ��
��O��Ƿ�ؑ�p���8�7ĆAR�iJ���� Zg������H�	BB�)$F�@t�a��ًs�C���8sxN�'nǩ��p��a�<}PIйc<{g��q��!�;���v��/��@�>��AGx�Q��?��O"<���sg���y�w��	$&�#%-
ɩ�J�3c�����I@vn2R��I��H�C|\(��r,=-�q��9����j���r2��O��[����aho�e]���D��K˨�4�KAB�$���mL�9D1ͣcϪ�؄�J�%o�B����55=Y�)�TK-]����(G-�5!#')���OANA*R�����D��BUS�#Tt�Y1L�8�$#_�J�8������b�t� g��r�R���f�S{%+'I��mN^��oIi����M��}>�+�@qy���LT��Z/������jP@�q��h�T��B��2*�ZZs�e=R�#e(��Jqe>%%�yJd��"%r�"��Y��@�[�lE.6bW҈��a��1��8�`H�^\�F�q,(�F~I�3�ȾNʫ5�Hie�ٯ�.V0�����$��|�Z���w����Q#�+W6
��X�e[V^�g)T�}E��"6�����ZȣHc��yXQ�祔��a�V��֕2�EJ�HU�V���]}�2�X���cz��!R~u��K�+���� T`���J�<��MzV*�AS�YYG�����h�ǆ :1��k�ԁ�����D�#�Ȥ�H���c߼�{���y�/y(y)q�2��BJuu�ڊ�,Ƴ|�}��6��1ላ�ALL"#�|�ll������@B�t%��Q�q��.1D�h��L�f�!"6�qQ�J�dZD!>)Il�bx?�~��NC�8==Y����f������8D� �<��P�I3��׶�V4��*�z��1�o�p.�(�B� 6�z4-FS	�(� �:,�y��KJ���O��LJN�#��q$�űS����]��ޓ�z;::�s�FD ?$��JD��"P���(:sU!����(ԅ��:0��W[p:���( ,ݡ��E�h	F۹P����ڂΣ���N�E7�8s�W�O�F�S�8~�N'�y<Tmۏ�Aˁ�h�]�N�a��3�A��9�����c�^t���+r ص[I��?����C�x�N��;e���}�Vv�n܍�ow��|�#��
������"?n�����/�O�>�	U��G�7? y�*}/�I��(-a��T��������+��7�G�.6�����n�����?G�"��w����S���}���}�*�R¾~�?}�ȯ�A�7�!滏��'H���~�"��a_|��o?�w��mė���������O�O�A�g#����gJ��!�}��~�>�|���6N|��ڊ~������$�O����S�|��}�9����N}�N~sQ���JI���#n�.���1{v JɯH<��G�!��A�;��ݿ"����.$����!��A�:��3'�}�8ҎB�a����8��=��B�D�����,CYnXsX�+����":���k��CH<�Q{w#����;������E@s�r��<�x���S�z�@����T�,�˔`��cH>��г�>���N ��b��{����"~�N��v�����O�s��ߐy�0ROB҉�H8~��Q_X��Վn-�\-�F��)*U���L$�>��E�8z�N��G�@ұ��'�FDƙ�Ȧ�f���>��T$��F�!3,T�l +ri��T�>Z��_�^��B^C]
��Ɲ?�P���s�z���H��SH=����ȉD^���d����Ejx(���Ԙ�6&�����U��D��6�� �\2����F���X��=/�<r��!+"HIN�Y%�Q�J�/ 729�F~L(�c#P�����J�hi��H�ȓ�����Qs6�)�g�r�4rx?%�dE^�J4�ui��zN�'+"l�E����<����O���xWJ�i�&*@��pޓ��KG!����$�*IQR���BBUN�S���:�������df䢥N� ^,�}���r�U�lhFmI9�3�P����!=��DC�\ b��qag��A�p��Q��N	<I�r��{�⣐��4既�V�I�aZ�y��ף��O5Jt���z�����$N�4��X�������H�4�q�屔�h��ON��C�{���q���a�X�D�]�Qx�1��h�`Su�q����׮ 9L���xD���|*�'O!���:$� ~�(ΰ��Gjl��6a�y�,�C䏻p�ӯq��/����q'J�YP��x�A�N�Q���ޖ6$��ǁ�>þw�Ǚ/�6��	l{2cY�	��L�̸h��S�qv�v��S�z�E��6N��	���>�9v|�*~ލfS�y,��)
�A�/��G�)��'�|��)%_����G��"�������y�=����|�Ͽ���_C��=��+���2�<��'�C��g���������|Y�_@�cO!�ѭH~�I$?�9�>��Gz��3�97C��S(z�y���8��?��	w?��u�!c�#���y�CH_��K�!}�=H[�IsW!q�r$�^��ً�8w)�pa�,�����^C�c[�<%�g,Fμ��={%2��@��%Ȝ���ː:u���FI��S� k
e�"%��"o�|�O���1Ӑ;~6�'/F��U�p�����y���;����O&��d���Z/B'�é��VBv6*�E�O;���h~��=����A̬�[��KV�Ĳ�8�p5N�X��"p�<����EȌE��9!��#j�B��[��9+<y�f�B��5HX�'��ĩ�pa�2/X�������9�;a:N��#���?0n&O��c����q�����'�W�o�%�8��c��.�a&�~�O�G�/��Yw�ļ58�r��?��+�����qh�?sN�\��s�F�ҵ8�`N2^��܋�u,��!�����[Hz�y�m،��� F
����jN/f�,�o�?���7#���pf�[�8�o}��/���A���:�[��˸���\$��_\��,B_�y?�E�;_`��Gp~�&$��{��y��?�����yD�ڊ��_@���X1^ey��_D�#o"�[Z*�0����Eo]��Jm�jGun!"����oE�k�"��So���O#�m���"�c�Q�؊��AȚG����	���mE�so#�i����>C]p��X���=qх��D�+C�VO��I`)>��O���ǟF�r��Kz߃�{�)�lڂ���GҖ����z�q�nzя����?A��ߡ��o��ާH~�#D��&��z5T��e]�V��O�]%KU|����e�X-�u8��/8���8�e+7o���G�SO!���In؈�=��g�B�ӏ�ܳO f�K��2�^x�������9J�G��aq�U2�Dk�i�h���M{���䯤��9�dY���.��%�(�}���B*�r�o"��7���[H�}d}�2?�I����?D*��O�F�?�|�^��r��ch��n��[Y�z�x7���޾y{� �k�![UR�����H��F�w�"�������������#�v���? �_���7����4�J~��~G2���G�/��y�1/��*�R�K��Ϛ�j�9���w��?���!�d��3R����=�#�(8B���y���;���cv q�vh���N�D��}��j���mœ�2#ip����.�-LWT7�:.��#����q��"�ߐ*F衣HڻaL��]�i����w"d�H>E#��i$�ڏ�v"��H�� �ӫ��(cB;f���'폀����*�CVQ�
U���B�S8��'��|2j�����9�9��'PG)�}E{���B*23�ø@�G_!�����=�}��}�s�1��#E��&up)��eid<_�b2q��_p��o���8��G8�̫8��;8��+��ҫ4��+�������y��8��sԻ[q|�&���Q���^���l_�R���m��@��~5� m����o�#�K���w���;H�%�<�z��?h����]{p�mx�W?��G_�ȳ�����k�C�q�Cرv3���>�{���Ǩ��?����F��5@^;�@SR�ۃ�/"a�Hؙ����xr@��H?	c� � �4v�g �w:��f �&�GOG���yL�D�IH�('_Ĺ�#�kRFOF��X$x�C��xu,�oer�f"��:�3�s��9EI*���{"�|'#�g<\|��3	�^����V+���4�1H�d�ND�8�%g�h&��g �sr}� o�E)�BB��2��B3~��OG�X;%�/3e��0m>*�MG!���OA9	L�rйk��0�� Ox�y2�Bf��DG#�!v�Fd�Zň,����o2�m~�p~�,d�|�����l��@�-ۃ	8i2xN��d��G�v���3qܦ"�>�3�cm�$�	H���H�18c�3V�8e�&�J�8��H{��R��	3O�1���␑'��xs�<��{�1�Z�1��	+�/�z⨅7NZ����`����3q���y��$Dx�D���fj�#�}".��B��Q�jb�܍P�G��LD{�D��l��O�9�1=�s�"�o	�z.B�x���i�@��pB�࿁<m+���O�ؤ�8��<X�0"7>���q�o!�:�@���Q��U�,ل�� m��H����Sf#6`�z/D��D�]��Y�̖wy�ʿy���V ��
���װ�sN�$�| �f݃S�V l�DO_�H����D%��"r�r\��~p�m�;N�Q�Y8滈ϸ����=�L�v�U���O'���,��jpX��w-��/w�+��Q*�p�)8����c�+�/��j{j��[��i������'�>��V� ��W�72�N��ohx��-:kJ������S~�,U�e�t�'�¸L���:v���h�1{���7��8�7�i ��"��䅟윰��{'OR��.�����?x�Ǟ�p�����u�c��HQQ��-�Z7{Y�~����h��$Z*��ǫ_�3����9���b����_��a������L���)�m�T����������vG�,�>iL[J�k!vNY����C[F��ڬ%I�]�k���8��=�:c~�>?͘���fb��Y�5o~�3�,�/K�祋���ؽv5��Y�KWa����%8��A���q��h-�����O��Q��/,��_�WSV��y���������S����s�#��i���h5~X������Yk����i�J6�+���{�w�z�#���ОC(niU�%��t���Q�1h�D��|q�&|��~|��n|O���e����������v�|6>�^�_.\��V�ǁ������(��6lű��w�ط�iY��G����3�����d��x��C� ��[X�VPH�MŞ���_���[q`��J�y�2y�{q`��f�ȱ�/�(%y�]�Z���]�a��y�����~3k">ߋ��|������ �D8�}�5|6a��[����$d|�6�yN�wk�#�F��4�vnڌ+�c;A�$�\���87e��X��Y+pb�j��0����뢮�� [5���
�Y8D���8�
��'�0�&h�y�#}�#|�{����z�]Doz���8a�}�!��my�5���)��D#���Pob�y-�!O��k��6���Z$|��	B�rd��@�,�m"R��#�y,2\�!��r�E���cy��w���N��v�Cu�lE�X�3?�y!����~(t�|�#A��{<����g���J
���='�m�S��W���<F]���W�x������qJJ	��"�����c��:�<��we�y-�ޥ�bo����z"�����(��cQ�7��Ǣ�"���TR��LFI�TTLG��dh���^��_�z�*(�e�y�y�(��E!�ӏ��l�0ٮcQ;y!�n�~��mC���P��+(zp32�&8�C��%�_�غ�BY�@��ǹ݈��+�� � ��X�*|�X,�,���+�<q	:��B��U�dcZ2u���A�8��/�A�O�$���c��LX��)�x�<��s	�ޓ�:f"2'ME�T���YHGJ�@�B��>���p�:T-\��i�P8n1�l@;�ۼ|#j�@;�_'�J����Yr�J�'�D�и�At���y�s�FٔEh^z��e��2Z�mF���=/�{���3�gc@�U��J|�A�;%����X�M�A�/���д�M�?�6*{
x�}�������~�� �׿�ևGZo-O����_��mo~��O@��L]��6�]�uI_�k�*@�co#u�C(]�J�=�#/��m�؂������B������ۺ�4ozII�=���Rq��Y�Z�~��m� A٪���@��]�}�<5�T�,,䝻����IDL_��MϢ��mhy�E�n~Il��,G���^g�r�Z�����)�|��k4���{�@������ٿ��%j�xYt�����Q�C�7�c�q�ŏ���+���2Jz���)Oxʢ��yh3
�>�PZxG�P���G�#[P��5�E��9 qK�A����=Wu)��*ڳ�y�䉷Lbw1�D.��Z4�Y�M�H���{���F�[�ą8?a"�߃��h��I�}i���]����������{���3W�">`���W��J5J���Ӆ�|D>�.L߀���qz�D��>���9�pr�b�f���A��PXy7aa	�Y��%w#h�B�'�>�,�g�}'�@��F[ȯ.y��Y{�9E8�������C��y���^��2?>}1Ӌ�� ���'��|����e
��c�	���W���͈~�GR��r�b�\=��x�ұ��yɢVq,�.{��/��}�t��F�W�s;���1S��X�bc��o"~������G�����"d�}HbZ�za�������$�/6�� ���L�	��
�]+�KT��ˋO��m� uF �̺�pt�F���>�[��Vb�􅄷ر��<�gW?��+�G��G�����ڰ�wߏ������ǐ��a�e!����.�w%�K�1l���|�s\�G�ރ��X�f.Ƒ������8�i+��z�-[��K�E̒��Y�rVmB��'P|��(^�$��{9�>��U[Q����{��ZD�`Ek+*SS����k{Cu5��Z����W�^}ao��_G��7PN�_��K���J�� Ͼ��m�"����ܫl�~܇fË��y�ɫkEܗ�1�W"�{Rh&�Y���6�DW_$��"���䣶"I4����V'�9��IN�Hv��R��;_���AƘ	Ț09��l�S�NR,�D�J�����G����{i�'�JPK!ܥ�2�G#��MI����|�$��F2�L$Û�Ih����x!�������#�ϓ��}%��gy��|O��y/��~
��D4~cQ2v"��OF��错���h!����k�ɉ��H��$�IQ���#�z��x��;�FOA��U�Zyrh���\�T����0i>���"�g�h�����c(T&;�Q?z2:'�f�E3��� ��9�.�ihw��f����vZ$u�SP�Ezu	@�����I�B�YNZ�/$�zMd"M!���]H���<?䑰|�)���l&f��$"�>`�r���j��2vjܦ�-`ڦ/G�Z��h�U�1i>Z'�C#�q�e
B���&/F�ԥ�tMZ�N6dU^�Q5z�Y̻u~s��3m�<��n4.y3�W+X�\%�� �RY����EˊG	ɏ�m�Ch_����
<�"
�؄�5�QJ�n���K�G��[�u�sh\J�^K ��Q��}P��H�y9�|�vZ� I3r%��[א􅼶�<T>�_T�z��ף� _���{�5����?ܷMK6��N����u�߻Y�ݏ�{���\� :�>��? 3i��N��.���.�>��+	���Ԯ	�+�n[_F�}���r��m%�oӃO �����E����~B���z�ۨ�Fx�m�����'�!75%��Fޫ�]7I�+��q��X����7�A�ַ R�HHp+�A�|�q܊����G9�a�}4����ϠlA_�r�J�L��6��Ͻ
de��-�� ���)���7@4%d��r�J ^!�/ms�A'���̫�4y�eh��?��{�D�m���LC���ε,o<ּ�>4Zj؂�~"�T��������0�3��֗h^��V?���עs�Ch��Q�D�y��ML��?��]̿�Mϣ�a���o���Pv�#(��1�oy�y��ATÇ����y�/�Q�ڳK���!T�z�L��u��}��`�:0�Y�;�ߊVBe�
Ӵv���\�J6<���O�D��<o�sh~�]4|{(!ܵ7��7�<�Z�/ymh>��- �nޛFT.�){��(ڸEm�EA����?�z~�
�- +Bኍh����^P�z�S�<�2v6���C�!jY)�����%3m�� �2��Kdզ�!�e�pݫ���:�)���oh~��'�G�O����pv�N���5O�i��o���mh}�e��J_�"��DM&�� Gy�d�W��������t��堂�,}�dl"-݄���|�Fe�?��V��-hzk��+�W?��U������u�y��h^���<��e[���>��b���:�}�͚��}�%����tz�dш�Z�)O���g_A�G_"���C#����Q��[�z�Y������'^G������8��B�~��{ȓ����ዟF�/�g���8K��X��bh"q�8gO�:y ��SV���hi%��QN��ttQE�	srC�;���G���H�2���q"b��"���0O�򺑎ވq�F��G��!�ޙ�wG����Qn� P��H��'bj	�J/_d� �g,R��ϩ|�8������z"=<���B��F�5��E����c��K���JɄɨ�:�Sf�z�d��� 0B<y����y�H��{�-�15娈9��ߣa�H�0�f�����MC��#	\����3g�<�o��(�ۣ������a�X�L�5�./t[x �^tZ� V��0vA��#ڸm1sE�i��F��htZx���F��5vE��3JM\Ql�B3g��#��cb�,S{d�9"��y&�(����(0��|Cwh��Pl�rk?��MV��j���Q̽�m��{��Ւ�֣G�tYy��r4�-}�n�6K_����c�m���b�6+�ع����V^�����������1+P�ڧj\�����;H%�h@��E�̵��%h���+�>e�汲o؀�P�<-�|�	h��:� t��?�`��c2��r��y��(GY�Ҍ\Itq�5$}!�;-������< `�m#�m@�+�&��i*`?Y+v��ҳ�m;p����o)*<	��%"��(��
P�a%=�'ݵ�iG��_#�m9'�A���Q�H�2 p����i3����x���4��tY�g|x����4�����[���v��&���u��4�2�,� �����$"�կP�j���Й�.o����v��Ng�ɓ�\��5M��P3�y�p#:�|����m���=��	Wi����?%f"W�<�aY���
-�n�A��0�:p�Aa��,�,�(��k��땔%���������?=��X��p��ÏP�ɏh�JGGK3��=�w%OPo��|���Ѩ]��i�c���螱 ����\LX��iܟ�(e����@���5k�ya>���о�=�|�(��ې�9(�>:����1^4X�P1��<Z�^���W�"��u|
����	4Ϡk)�4���	]��C���l^�ʽ��I5�W��m�*�bLԱ��d��#H[�,�f�E���(��^4g*���X�zEJ�w�4�+�1Mœ��i��h�ô�������Ѻh-*y8�x$yW�].���(�����]�)ȓ1z��9�|��Պgi ��>�O���i,W3��4��}��Bp�C�����j���SW�m���dg߇����Ρ��9E������׫w9Ϟ,�UB�l�� �?Pp�6�[�U=��Y̯UO*HoY����Cۄ5h�yu��q�b�,�SV�u�BtL���ļ� [+C&.�a�*jݹ�B��3�&p�d������AC�QIc>r�&���y�M?�(�h4W�ۀ����p��(#x�݄��#��z�l���5�Q���������1�0�EX�D8!+����D�)Z ʙ��p��D�~�tv�ݗ�� ��X$�)�����
 c=���N'�9� �J�t�1}L'�Ƒq���(��tO��/]��G�$��'Ou�^={���ӧ��%�I�;��*���JqF��3R��ࢶY�N������qP4a4��s;c'���]��Q1n2�WR�E����IA�B���E���r�G��Z�Q.c�o�sg���K0�&N��r}G��9�r���٢n���6X�@�0�P7��G�8�N����Y+F�<���v�8�\�e�������G����Q�o��3�0�Q0ʒb�ƵD�%��P2��C�a<�jO�y��Г�sF��=�qI1!�r�1����%B�U��8��%N�Y-_������fN袀��4 ���P��gʕ��!��ϼ�&?6�3��2�����s*�'-@{��|Z�� K|	�0b�$��~�4f��	t����o*���2�H!�򐖃��[PgM@"<�،A���J�z�D��ڈ��8��`�F�l�%���P3~�9u�������3���:�� �'ڈ�'���!��V4?�4N�Q����xٌG�p)���ta��n��x���3�o��g;`�_�&��qp�G�o/��P��������"[e]@�׊'�v�5��}��Y�"�eW��nSo�O��h�V��n�y�6)�NP�P�1ծQ�8��h���d�<��R�Y���v���C�6~�$�N�PiC8E�5c��P���9��QGX6�Ns4�z(�0�f��4�pʦ��x����'tD�3��fL��y��C�)���y!�\P���^�֌�2�������q�u��&ש����'���t���\��qK��`#R��(�����ʲ1��ƶ��Z�u�9�򛈚 ��i����F�ih�4��P�fo�󘅄���"��-Z�����h�X��q���w�x��6�1��W�;	Z(�X/e)���B%e������^sQ�6�w��d%�Q�:�i,�^�̤a?ec�Z��o:��D��Dty�C�(_�zy,T�K����X����Nƃ�j�y��]��H$<�
�z}�Ґ��z?�,�m�S�F�f�".�OAJ�	����>����w:h���Ӑ���K0I;[��Ϧ�zT�W�7��ھ�𴞼L�壖`���ȝ��.L��h���v�٨�t)?+Q�>�6���2��{��T4zNc�S?�,D��d4��j���(�SW���(�#$����'?����cQo�R�s���y+���yx��2��G����?}�	¹��!��-��������W?G����'����}�A3���E�r��`,��a�W�^	sqG��+B흕��9���=���#��Q�{�sR���P{�y����]p�ux�0w£��E�����.�
4e�2Z�x�"�b+��J�qS�&��uqvn��uUo�D2P<�!ѓ0��M�k�=�ʾ���x"�#��`c]yWg%	��w'8r���D@/k�?
�Ǣr�t�N���1c�M�l!Hz����4d/��
�M�?��B�j�;jQs
nC�ĉH1�C��r�Pj�a��p�!�x�TQ�	jM�6k780f#$ '`'b솮Q.�0`�I��0v 9���QmE��x��:��Lhki����-6hԳD-�^�ۑ��!�U�F٢f�=�	j�N�:P�����]O�ϰ'n"���ۦoKa�.0��O�u��;�w�S����3LwC>�%�Ll	��7�d��xS`""�F��%�y�K5�Iy�(HTP����+�8*�6y��$6x��Dؓ)؅���هPk��E��=��.�~��*�ق�$ j5�s����s\��� �v�s(6�G;Oy}g�a�,�ۏg����i�<Җ�i����	-����F�@��%Y������US�'��7�Gqt�6��z�Ԣ�hz�SyN㨜���g�HF:�y0��@44c�l�A�@c��7D�Pst��B a�n��M]X�g��ßymBA����]���JW���T�5w�8<1��&��f�Y���m�4��3��������IcJ�`�`}�QK4���:���^�|�4�A����44�~H�G�"`��,��R�=�w� 1Ůf�Vv#��PfF�@�y�5Z�jE���1��Z�DZ��m4Ԛ̼�lBX7�C�%���=R�/S3��.$��l��-�i�k�ҕ��j�)hƬE��D4�z�ƒ�&��Q�h4�F��*+oTٍF��
Xދ�=P%���J}&]H��"b�-�!���jԖ���?A��1��Es�Ѻ�TZ-A��8���/��B����7ٍe|	��>�ф�	�r�\��򟂰iQ>{-�<砊u��o%
6�$T�^Bu��=�d	��Z\Q���<�f��#���Y��P��{��#�f4�m�i��Y?�&��q<j	yE��P2a�FOF�;u��i4�@���k�}2#Yf`�h˿j[z�PD�擵�t^��"� �����\ԜAº�h�+A	V4`lǣ���0儽(�0�=g|g"ǟP<nZ	��Z>O��L���I������ߜ�A��8i��na�Z����O_���tR^�4#V�4Иn@�G;P<a:��ڗP� =�iv���̳tӮ�a2Mܙ�4 X��'+�#��{ӓ��:�Eݿ�<Y~�����} 7@ȿ�Y��n�Q�xX�#�y�<v!�GR�ݏ�E u�=H�y7R�.E��%Ȝ���W#c�}�X̲p�3��e�<��F��x�;��o85�q�e����eZ�"���ܞu��9g��up�9;g�����A6�J��:�ڞ�w��](N
�.� :�}9LH�@�
q�B(/�m4"w���Z�t�w�B��;�&�x���)tuC�#Ş��f�H��t�F(c����	4F�����̼_?K7�H_O^�AϏ�OP��xz"����4'7�zR_M���	ʻ�En%���h�p�%Tz���� ���e�VB^�I������=S��!��\h嬺I���Q�(`���Rװ�.b�ScJȳtA+�k1gcdl�n#6���f�H����6Cԏ0G�1Q3{��K0�W�������t����V�<W��6#;m�Hi�ӊCB��@l���L�yμ&�F@�G:��������5�T+uJ�����f�����V�77F���m��q����-	P6Z�3�Z��7و4��7�'PY��{en����܉0��
K/��� ����&as����ok�A[���	�VZ�V���T揼��_�$������lev)!���gPdHȳ�C����.��l��Q�3��NZ����� 8h� �䛤s�7m9���(/���c��~'�ʒ���h���\�b�m��j��4�5#�Qu�!j����D��sJ���z�ꯏ��F��v3���o�W V�@�y��yI�X�d胼��bJ]>��-` O��X>����K�Q���{ޥ��;F��.}4�X�zh�?�F���!(�}8���峂���������2U��C{
v�Oy� ��E��n$撏j�D��؇(4dc{�*n4D� 44핺Aƨ�s$*������41G�0��B���h�*L֍ �[���Pʪ��☼k�<Y�-�?�鼄��:��*ֹ�Q��`�&1e,G���{��rX3�3
h�fј��N�F t�L5��̽����h+&L]=���6~��/A��T���?D��\�mo�Z­�x_;T���l4넫V��+|�o�D�ݓc2e>�f!�e�'!���d+�az�@��Fd8@]]���L���y՟�G$A#�u
�X7�N2�̊�b�&��h���Z��(v�$Godx�E��D��Z�&�����8Z��� �.�B�,�����vE��:��L��z�J4�i%(��E��H[��X�e���mC v	@��T5�2��~�g2�g c�\�J=g��u*��'��������燁j��PC(:�|i�MD7��(��_��R�]��F�{;Q�K#�i!��k멆%P��� �˶�E��˗+J�cG�����! �N�aN����-o�����$T8���O��v*�� �eIV��3I�߬ɫ�7c�g�C��e���q���y��k��p��A�ݏ����iH���F�򤷾���؍cs�@��"�(�;������@��lEN�m�r��v��F�[{��|/0x��Q�� ��@�C9.^=g�7aOzQ�qGO���it��,,�'�����*U�c@�����G�8@�"�p�R"�#��{�Pw��	��xB��E��"��q�/[w��>K�����B�L��B�����c&(O��,�Q�yD!�'�y���l �]e���|�	���&��C(A%��y��<��
�tp��*6�V�+����B��к(=c�ȾֻewQ�P�n+%�G�RB��I�Ӊ������M����nCt�+�߃��2uQ^<�<�=�(�("p)��t=�oe�ΑZQ��k�uU���݌��C~��zl@Z�#�O��<����E�[�ʷ?gڪ���� ��؁��>A���Nʺ���-��@�PK���2��@�0SB�����K��@��n��3:,�{*�L?�9z6>��Iu�JP����d,��B�Fݩ��^���&�n�������.cؘء���4 �+��liCﭣɣơL��h5�G�x*�}g٘�Q	�\>���H�nPAS���ېd;���/4s#��q�C�0[��d�������]U�\n���+)�IOI��z(�7���c;	�o}TV�a`�������<Wƾ��!#*Q����N )"(��2�B�̓	W�Qy�0�ܢG������C���nA4E��'�z�q�p���U��ӂ�[Ң/���
A���V!!F<�.r����&g��a���s��0N�;n��[�����Sэ�㛆��.3G�uz(�m4���g�񙆨��Gw(!�iM[�6n�=�ez�+~�M����0b��o��`Y7F��&��e�ಘ Z2�EL���^�4W�9��<l�3���<�����؛_���V�1I��Io`<t��+w
�sJ���E�@�0{43C��%
�[�t �w �� K��۩��i�%�ԑ��P�����H�$��t��E���L^�ʵ��jA���9yy�/-B*!�"�������@6�C�S�2NìQm�A�C;!�Ɇ0g59Ʈ����F/����,����[C�)��#D��=^����4Х���,@.ݴ�t�!���,��<�U9t�Bִ��@��Uls�l�Q@#/��wu~0�P�(�ǸLRc�������aKH.�e�v��t��gG�'�cI[���x�	�Q�L�J��j�<�Z}��S��\P�����Mr�3��s"��o3w�ދ�|��y�4.�mPM}�nンL����/嵅��?K���gх��ș�$���(2�C<��<�=�g:b��C���H���SV v�R�L_��Yː0���R�l��F�Gqd�����7�^�k6#�UVШо�Z!O�mMu"��Bԓ������%�&@u����]p�GN�;ᄭN�:fa�严����� ��׉ ��� K�>B��h������F��h�j�]�g b|�!���3�.�*>J>ųH��z�q�`&��A���Y��<��!��2�C��@#<fE���7�͗��pw �v����m����'���ܐb�:�4IutF���=G�Y��|�\w��ŋ��(퐠˄�C�t/�Z�X[��P~�[��x!���i}3�X#�FyE��B����#�'ֲX�2�N ����*:Z�}E��*"�H��L%��P" �t���y��^��G�Ư{�Ō��`7����x�Z�c�
	��Tm�nJT<x_��J�� Ozڸ�@^O���9=��iBp���5u��A�F��9�nT��%6����<J�[��H O�	Ǝ�"��8�)+S�_��?�HuQ7���B.���lb��g�e��S����a������-�+e��5_�]�(QB^��PJ�Y�3�Xx"����B\�J���k&��B�� 
�5�٢���������$~��p7p<BZ/�����O��� pixz�:�yk�G��ĺ�G���j�l�4�B�u#P|�`�߮� ���Rq��zB�-��Wy������zTg�[�C�˟���6�7-�6�[^1���sҵ��ފ��,�D��?���3
�����恄�A������Y�7�R Uy�jo2B��Qq�(��'d�V:���k��=�d��ѦC��jc��8�6
���f������(��Dmˮ3F鍼��樸��>�ƃ�k��XҬ�vs��i� c$�A�;���a-lP�n:�S��Wi����V�=I������E��%lz�ٷ�BAs��9�p�r�S����d�S�����C��V}�K��ի|dl.+����A��KPe ������Q�Q9Ȟ�k����ρ��;mPv�-�۩��փDC+yq����'YoS< q�!���v㑾��������{]-�� ��Y�2�@<fUY(�d.�R,}�9�
)�L�J.��S5�o䦀�T��z�b����+GB��� h\�S�>[�F�D���XN��K�-Ӧ���T7��J�'FY˱���H�_Gx��ڑ.��Znᨼ��Էb��d�0+w��V��h��)o�����V(�&��MB��*��c �R���N O��x�J����9.D�H�Gϊ�b���\�G�J��]��#�˄q%��Xy�����cPkO &^ |U�h���W�/�3�D��LhL��0��L�pϩ����q�ՒG1��勢�.!�-A��e���K�#s�Zįx�<��>SC@�? O�>��/8D}��k>�9z+X;n�c��ӎ8��vQ\{a�X���ik�K䤍Vt�OY��9� +��7ι�(�u�&h�e[���}4�e��t�(�$��7Q�.��g\�������Q�Ry
	`�l]Lh���^�^�+Z$��MM.����*ݼҍ��ڹkŁ���{e,�tG�h��%غ ��OcZ�3y��`��Y���
@�,�׸N�R�
�:���	y�Vih¶lf�����АQ8gd�<y%�Ry3�� �'���œn6�Iשt�
�t���.V�^�U��~���(:��ɕ ���5�
#,(f<�pH�2H �%�I7�#!�m��Q�<5�]�Ǔqw�n;%�7�g��/N,y�����v�e�>�=0��b.h0�3��H��a2QA^�;_ ďyHz�-���jb��Q6���F�S��nnOx1B� }3.uL[<�R�ϙ���-l�Z=_��
~�*�W�ב^����!s�J��>�L-��6q6�J�U���I4U�-�wQ���#05E������vkԏ�E��{�ȥ��-clD_.h��Ee),��Rݵ�Zd��,b�'��3�&��9#��>j� l���~���L�������(��0,�w)X��n�;LX�e1�ih�5�*kz9�G�/�����ˌ�D�w���ث81�������(�q 4���[�)ob	��z�V<����S���ʼ&8Kw}9�Z�2C�F5�'O��@�2 �9�"���ƳP������v��J`!��\o�қ?c���Yy����8��H ���7��8�Z�c���Ǔ'�ǜRްk���9�t_ҝ�G��d��0�o'����#�ws�/al�<T���(3�7w�v*��3W��=[q��/ѕ��=y�@^^)4���4��(�ʍ��T�Z��i��;z��PJ�&�:#��S<�Q4BOڏ�q'_�۸ �:���Y���y�M��Nir��NR������مH��<=���s>K�@�Kd����<�i�_�K{�C��d�lBq��b����S�i��xs-}�����Է�2� �p�ڬ}_m�׈���]���
��JQ��!Dz.G�I ���G���Ѣ?r�d�N��bݐf?E�S���G����ޕZz�r_I�,���/��W�hU�^�vȓ9ߪm�+D�ڗQb7�zlt��#u�����QLBy����m�c[�o�D�rg{����4���'OC�;yZ����!��P�'YS�}�Ac̼`|.Xx!�c
.x����EԄy�0�S"z�b��\� /y�H[�1�6�uϢ鵯��ɓ�j
*���ϰc��w��<yG�lq�����q���WNػᤣ����u"���	�ٻT�{���'��Y:��ٳ�Ӂ2�N`� ~�փp殎�����%l��s�G7m����������nrO¢'	`g�V��|�� �@[�����Iױ,墺p	y�ywr΄B��<���|������2�#��)�'�<=���+ L6;kg]F�*)�� O��@��[��j��R	DȓO����#����i�yS�Q!Z������l�fc��(Z�Y��t�e��k���.Qgw͐G�@� u��k�f�ʀ}�.Ү �M#l�J%�Ak�YS.y"T�r�^��?���h=y"�#	x#��J i#d�$y��^�+4�vA�x<:|W��u������4�U4"����@�,��	�%����������Yx����PK��]��X��*�d�~#�fI�>hr$�=��-�א�0�~��򂆖x�����#t���}z��b�V�<�.F�L�N�a��!�(���&�d���LP;�[-���|�f4w7R�\>�t�'e[�&H(J�)�ƷY+�C��d���V�^#-y�0��jH���~Q{���n� O�
X�n��f�1i�M�I9.���
-��u��v��/�N��^��t�J����/�?�}��q��5�v������]�x�2By�4�3>z�P�4J�
n�������1�E�����Ͷ�+��񾽠w-�����&3	y�Ƚ� ��@XiA��Wz;!�&}�!�	�w�B�]��>��G��*�r��W���;��Awp*��E�����Ղ|/U��X<�|A��w��4����e��#�d1N�qK��%TI,��@9o�]l$~d�pt�=8��i�|�tfU�g��\Nz���A^n9��}���TTrF�]f(�O:�EwZ2��Q|�%ʆ١؀q��J��*�w�e��#��������}�ro�ȓXv���	5�5(�(Cjq>*3sQ��.��^�Dwd4S��:�F؝
�
h0��ﮀ8�k�����\�8�`�$��<�����[���U�B� ���	�e��	<�p�g���%��[Q���J�|}��K�g�O`�Z���.�4qayvD9�.���:Q��"���@�)A�̃�r�-��ׅ6�����2~��I���d�i�6&�!���P沘z��#�;�L�b	�Yz"� '�x
��	��*N��N�1�VKv����}��:��aￃ<�>�g�六5�1��Tz#�e)�~�s�s"B|�#"`6���A%b�|DO_��Y�=w��F�����A����^c�uqL޿����}�Kl{�:��aw���aB�QB�GV����1+;%G,���Jd�����^�9jj��&V�p�L��;C��;@&8��ﴽ;N��B���<xA�г��!ﴵ��<��=��Q��E,ݸy2D�O�t�L���.ҝ��5R�&!i�x$x��ר�ȸ=����K$�f0N�<��� ��m�����b��Ĥ�y�Y,ȝ�-�����B���8��}8`愣w��ށz8�G+��"�Wh&�h[䎢��7G����̡a�|~9&�	 ��k����(k�QdƝZ3τ0$K�����̭L��ғ.V�w���;B�qr�=�' )5�1*�6c+��&��Q�D�ʵ�
�t��w�"@�g�ӂ�֋'rEȳ�Pc�ۺ��٤'09͞KP��G@m+����,HM�kC�O#�
E&^�S�Z8��i��F^��
R���G�5�|����(n�:#'T�[�lPG����a�ht���/��yR�ټi�I�A������B�<3|$^10��ǎ{7`���u.p�p
C�Q>��@)�S��@�0������P=�I�.Ud�R��R�W/����dH���e$�C����\��H�Uy�	�q(2�s'���D����)�i�J��X<e��P�G�d�(�1���!M�z��;�'C�d6���U o�%���m3YMw�w�@d^7 �7��F=n�P	��8L�1�?Qx3A��'�0Ro���(_�P^�s/Y+P����(л
��liu"ۺ�-!f�dh��A����`\
n��� ��f}�1.97A��Cն�v}�Y���n���˾C	���-xg�/j��ݒG�� ����N�Z��D;݃�[��p���C�@C$�\�2����;(FH����m�/�0I�;IC�Cs|A�ی%�s�c8��Z�D�s9QA�T=¼��K�M5
��qç���#�o1$��"g���Wt�������j��Vj�`∝7N� �ޓ0e�V2ȶ!�L���"�Iz)���|'�؎��T6ԩ����ջ� �c>b���FFH�o��FHd��ţ��x�3��ÝM�k�t���MC>����:��nb���j� �c�(�-+��eJ�d�?�t%K�mYf��9���k�2�S�W�'�'!t�١�FO�m�
��x	+�"Æ�9����@�u5K�܌�e5鞫���>�Kmj�=ȓ����:���Ǩ��}QI�,�׎����u��%� )�N�h��fR��L�����5 %~3�=�^t~OȫnTy�r�[]�t"ǯ$*��[§;�9����2s_��⬩#α���N%��D��Y��Y3a��(ȋ���V!r�2D,X�s�����E�;_��b���r6t#��c�7�a�j9��<	o6�g�'�({���O`;`~Q���7l����(68lA`�����68aj�S��8e�S�Ϊ����4a�a)�y4}ԾVx���<�ut�I;G�$B[�x=�y�[�����q�Z>� �^�K�}�@�sՎ˓�!�?��<B��<�1jhi�e2�@��̍s�Q=J1��x®@^&�Igs�M���uig-�c��d6Qo`�]�ֆ��\$؍�=��V.82�����i�ΓW`�\CK1Q������l=Ҡ��|Ҵ��t���ʰE1!H��U(ji��RY�d�Μ�����xW�<bj�+AM�e:*nX��z���H������n 5�U��G0��'��x;�;�k�n/���+���U'�����Sݵ�c��e�>`����<�i��\�8ҍ	��Be��3j,���0�ɨ���Zs'y�>A�5�Q�F��@yu��@^���o4:��B^~)��_��_@�f�#��LEl�S���Y}c���vlބ��A0�w�>*�Y�LQ�}�����Pp�h�2��Ƒ�dc� 8�g��m��u1FZ���Q��!�ŏ~��zc���e�@*!����!H��.$���=�Wx�p%��"�"@��o��D{NA�w�h!5@-�L��j�9E ����ERd*�_���[�O�ߠ���!�P�s�~��P�ͽa0�o��̸jdx�R�9#c� 5O��߅<ՐH$�֝~�cDL"lZ!�s���$�Q
:u�'�}3�z�`��:���@�M#��<,�m7ф��	8���!o�`c%���!m>]�52�G!̆�̍^���"�Id�#�DI��@I���`ÜE=�&��&\a�����{��ؿp�zy���Cg�vv���r��_@^�c� q�\�A�fc��i��;����w��������kڝ�����AsW�a#��:��!k0���3��B^{O^�H=i�lCNU)��4�~�G�t�uE�Sݷ<���ewD����"��Y��j�,�"�%���Py5��f(��S/��;�W�����2k���1����;���'�����#��n{�OlB��h�|='2��ܔM +�2 ��+����JR��Sg�V��jAΗ�&�B�����4�KQ1����P4���P��0��D��LU3��G١�v��М�0vF>���~
��1q�����=�5�"�/��e&3��HfΚ�㬛BGOB��
����ą�3z o>��.F��E�Z�K���ݫ��O�����izq	���c,YHs�8�c��b�����+�6��nK{y}E<{:�9h��@�of�� �/�$܉������y�|���	_G=p̑�Fh��	t��iBV��h���E��hy�Y"}Oyg�[��	�M�p��s��2�P����3��;j��	ԉ�� kg������r-�R��|jf.��x��.�qHf���t�<��yk�-Y�Ȼ�/�>_y�J�ǓW\U���D��فS�>�}��!B�C/���A����u&��Z��WJh+�b*�pB!����Q27� ��Wnd�j;4�;��P$�>e҂��+c�x��ǃ�}�<�b�<#��7����J����f�c�8;-=��7R�j�jE���v���K������+@�HK��b��Z	�͆�)#+5�@���kq�����[�	T"�ˤœK0�1e����(��5;��W�g�f62�@�'��i!��֒����
������+��p�k%Xd.x��Jب'7���Q�nC��O�ccS�K�,A�f�����F��٪A28�EF���!h�a�G�"d�l���WY�I���A����_f��k�:�f�]��|7�,@-�$�O�]Ex��������#���
��\OX�a�<���4��B����FM�>ۚzJ�h5�Ճ���<��e���!��h	z#� %�ɹe8�n�_���)zj?����q�@�ޢ��;� ��a��o� /y�Z !Ku�
�����(	�yR��^���ӑz�t�"�v�&�X����S6����%��}�d�Ba��o�W��!�gPb�k!�̜�~�ʪ��r$eH�]P� ����D��
$_�q�'O@%�ΑZл]y�x^2-�<m|4�gM\���]�O����ػ�I����j�C����r��U!��O�@����pE��f��+�Ȼ�A/k���	�	���B������-�M�s�(�͜l���'��w��<�Iϲ�z4�!��p�n��<�9<�|!�,c�0패7���D�iH5�L�c���"�s.j��	M�� ;���	y��vBH499(����#d���!戦^�'|&�D�&8D�v�=8�d	N��"|�%�l�j`��*���1qC��$�-G�k�ҴzL���y�<�0�<����	o�Q8��!HlN�:飧!j��F5&/�� o]��\�-v�G���<�#6`!�_�ￃ<���a�|�D���0��`7i�ΙP\|q�g"�)�i�F�O�,��X� /t�<��_���qd�j|���h��gt���k�SckyN��@�_L��qX�*����{����#:���^�^��a���;`�f�^'=>��^���<-�9�a鈫{z��hr��	o�u�3�2,b�� �wB��U7�L�1v⡓q|AvZ9I&:b�䄽�X9㘭]<)�8jc�cvvv��Z(vn8�s�D�(˻,�Vf��^���8W�Zy�^j�m��/2�Ǫ�u^j���@\��A�*H,\��M���B6+^jb���B�G��xh�)��3�ȷ�@���(�6���̐od�|czZ��S^;ZzJ:xz|�ƞ,�"�`�������n]�Bb�����jh�;�AMf�I���n�>�7y+F��7Z��P�3������Y�|�1ҋ
�J�ԋ��Q3����I��I+�Tb�j2y͚Zf��t�����E�3 ԍ�Ś�d�<+�⽌�L hIȓ�ZR���ٵm�KQ�ʧ$�f��=9���oQ�z��h&�f
l�8�Q�5��E��H[w?� -��hn�6*����L%T�8�����h���y��+bcr�B��f�Ҽ<��L]���PM]eN��H޳/!��p�*u�!*n��!yƨj��a��`�'�|�C��w�L}1�̹0>{#ڻ�}�Di�'��G��T�O��-h<��G�!a�d�x�1F��	v�Q@p+�~ ����yx"��y�ċV�s b�>C�ݝ�6�!@��i!�*AN�Z��R��Y��8���H{�U�gي�MOy��3 �y=��~���#�]wg/���i���>����<�y����Q���<��4|W򆂎V����D;�F�VH�y$Rn"��$�E�(�c^
�eݪ����#���u�H�A�.혼D��� :O�ڵ��끥k�<Y���H4B�V#�&�3^�w#xk!/���J�0P�}��j��M]�N�q���7;Ol����sW◻����BG�߇<ѥ��
�
jQ��KD����Qz�4��!�e�n�|Zb ���e2B�`3��Kl�s�d��1�;yCiT��!r���<�|���=3Y{���|'�WyR/�%#��P��v����L��0GbD3��y���1#l�<qcf!��i4���M��8��LC��_�*9�%%�-m�V��C^A�:yZ�+;�s6 �ԓ�D�l���4�����av�}�	~fc���8���0���%S�e�8+ �u�����'�K��I��yR&U�v"nӇH��C�sB� ��ȋa��xM@��X5�7��LN)d��g(k1: ��Y�2W_�D��5�{���<u?nu�H�Ҟ�%Q�5w �ͯ��y��Mf�K��v�Q�����U7�yy39in/�E�^��Yspn�<�X�;�lC�7�/�䵚^�<-�������ˌ���$���a渫�X;^"��v	��t�����Cd��,o�m2AJD Pu�Z�����x����$�D��q��G��q��g��㰳�x��������������$����S3n{�N��S�v'l�	��:w���0�&�!�!v�>��{�0(����w2VP�O�Q����1z6N����4dY�^�؉ș4�~P�=��7����:��
��0Y黼�� �HI�GĮ�px�z�&yշ�q#k�2�:yT<��g/0b�&�)X�V�N��1�Rlb�@O�v2)@Y~��[�+c�Dt (�>9��\��9�F���BM���a�A�#,�{�� '�s�<��0�7���[�����'l���7�_?��<��2��9�!����D�o�B�����b��6�o��z�� �:Yj�ܣh����dܟ}o�x�d�@_��s��Pϴ�7o`�������OX������h �^�iF��4�sĭ��[Ҭi1�X���7"�˗J܀pg��;�Q�mv3�8SQɼ�����N�v���'_a�Y��]����F�"�	<T�s�6�1��Dٝl�tRQʟ|9�_�Q� d� ��R�2P���G��[鮭�!!���x��8%��LN�M���V��{� �R1�y��'+�Yt��~ 1�S��g����"��(%��Gv��<�-zJd�Y�u�!d�������~T���b
�D�BJ�����7�����'$>��H�k�x���2-�<�ɼn��'M�h�7# D%��%Ku������QG���yJ1�3�W
ʻС��`w�[O%��Q��y+��fޛ '��{+��	�JW�v?��H�u$�Sy��o�T6��f~8C��~�p��N}u򮥻V��6);�3k�<`<��"8�1v���;F*����'"޼����'��Q4����KZ��O������K6��ߢ]^Kv���S��4�L/I39(��-$�����*}2�=М��4d�Id���Q�?�܆�7�)�g���}Ԥ����Hc��������ZI�l�Wi���G]���O���j1�637ҝ����҇�#i X��h��޹��8�쏈�sU��T��e]drW��?�y�F�K��"-�2��PWp�]�x�3��XMa.�4�MQ.�2s���C�� �ГzÆ�g�BnuUB��E��t/�bCi�0;�А�`�bh�c���i�H�(~�uA��Kj��v}Rޮ����bU^��G_G��dTQG�s@W�4�8�\��&p �F��,SG���D���en�������Xޟ���F;d��H��է���j�2/��)�����D��͝�7~���~�D�%j�2��X��	0WM����ً��p9b�/Ǚ����{7�mzM#���􁼊
e
�?F� ��1;������|�غ)����#|�g%�[:a��v+���#"]��[9(��k�?����c����v�
�����9�xktt�Q���(]��m=��gZɲ.��|/~G	�',	���8b�&�����':Y R-�Ϫ+�01�u|�ݸ0f<v�Zb��3"�L��8�5g�F+ГY��2ۖqok����C��Y�If�f�����s�%Θ�����p��H�*��Hq
��yK���pڢ�Wz=yR����z�<M�4���#r�8�a�9��1��!}3�7�D�9[c��S>���g���|V0�Oy"}!O��
�r\y��2v�y��rM�Y9���4z�а���Ԗ�����QF�K�B��o�������|�Pl�s ���G��M^�%B�s����x|�>�:/���x��x��ԇl$��Y�S'�����q��&�0�<������9�Ly��ZG�����N�ת)�ɚt�#�Ee��� ���{6��B�K��āy�S꠴w�G��j�8j���dc$Y8�̜iHذ���꒬�Y����K� sB���å̛2}4qF��,�>��76r��R��б�_��<�O݀�;�Px�����[�l�ST��‣?!�@�o J���d鮕�E���7��P^Mk^�^�،CĆ�@q9� ������'iu[y7�x�dAٽ�V�y�Z"��3n�!!i0�X�d�t�\�����D��/c�rn�N���w;
�(F���-��h=-�%�W���W�'�S҃��[]}?NS�$KW]�
���)�kE�3�C���pw�E�K	]</�?���1�?��l�o�B����x3I����U�x�̘�������Ȣ� �d�C��,¯x%mDd\�@_�IW�tI�5D�P#ı��(96�~���Io\DT\)W+}=E�1DMق�!�KVHལ�O2S4�`'q��n�C��
��Z���|��=�#�������ݬu8��W�*nQyr��'���W٥ЬzI����w!�=d�9R�=�
͑�C	p���I7s�J���$��!v��� ����7���T!��5�K�U�)�9^�����_�y�eH��L`��1~�-�Ɗ�g� /�u�4!t��N�NF��%�[��cf(�������8� ��Ҍ���	yŚb������}E�_Q��O�˒1y��]�qt���O��d��Af��%^z /f���8i䉓&!@]��}��� �Z�afv�dn��v���M�$"��P]W��4�Zْ�ʖ@����Zd<�*4֓P3�	%�!h���If�ɕ�x���"��	9҆�K{�s	���]wmڴ����g5dGy
&��]+�I�S����>�3��g���6���}v�����Sp�"B�@�ܕ�����"t�D�\��ً6s>B�,��ek�����~��^������҉�_����a��\?r~'��F��͊[K7��qR���Q��~��汈�n_k��a?۾C䉃L������;�Jxs%�1��z㤍���݆v���Y�=��C�@3�<�/+�$��5.e��ÄK� "�'3t���G	{'�x.�6��C�8�叠��T��I�� �L���B�@�,�r�������DP�|� g�<�O����;c*�V-E�¥H�*�Hs�����\ȕ!O ,��	������\��4=!�;~���k����[`��Q�3A�@-��Q�(f���A�%ݴ�գhlP$Q	FZ\}E�/�ɬ$�sH���0y��#�.���F�6�{�$$|��V���.��@��8^$�8���zϰb=��o5��sB���$����׆��A�x�.=|9�o�>[o�O\3���6|;����J���f%�8��[1�e2�N���r,��
�ԫ�z����+z�l
��l	y�h�E��K�cC�o O*+y��m:%�T��Y�%F� ��ii��J�F�(������������1�i��Y�m�;����7��*���_O��m�'�5'�!j�:��� ��lL���d?�8"7n�>� 5i�D�J<@���y!���0	�E)鲛~�c���6P�;t�;-�\-�94����	J�~+q�������q�@$�LI�������z��d�H.�5�����w
�1��_Es���N%ݓ.r�+�Z����)b����0��3l�R� x�㽯�g�]"7�i!�Ɗ��O�u3n�։K���B^~�J)�<%��U���rA�'P,^F	Ż�l>	�w: �Q
X�	��L��E�ӂ� ޟ!�`���#� z�j�.|M[�]+��.>�|�Z�I2��6�����M@� D�0�7Q���[ 9@ƿ����:�G��&S����gh�~8�/���>3���{�﹏ѩ����j�O��Q���Y���]�
b���f�#
q�
�Ǥ9g���z�yyq#,i�;�4ua������J��!����{N�$� �e�Д�(=~%Г���e<%~�Œ?"�o��]�C��'�L����5h !���]���h�W���7�G���ZB"p��;�	y)�ȱ��GOt:�]a�W*e�m>4��|�eiP��N�_�(}O��L����/�N&�E2n�i�7r�1W��8O�u�z����Z�5�y�S7َC����<6�%j`MU��|ߠʿXk��oF����n.j{�h��iP��pVC�ZQ8y#�n4R���N�4f�=�mQ��4�>j�E��8��.F������C�Y�k�"��^d�MF��3Bh��r���g�g N�O@Ē5�Z�&-Aȸ87�`7{	"���<1N/Y�}�?�2����k��u4�#����~�F��4���a��v�9c��v�vY�]��Gt��=��vS����w����𐱳�}L�}�8ʺ}�����v�I<d=��x�m�~37�#���C��$c[}���r�)��ғy��A��	Gw幓پ��;lN���*��ݣ,���Sd&�V>f宼�r��?ғ%ƻ,�,�Cd��,�"޼8���_$�g"��OCҔ)ʛ�2}.R��ԇy�X���P��+@^s��ϰNU��Ry��ȓ���
���w5�p��>Z��C�(3��G��l5�B���(ˢ�Ѣ�cA��R�ă'[y홒���M�Ѝ�S��z<y2�@V5� �Q�1��x�4����x�?w��[㽡���VғƖ�d�睽��x|6w9~^�<��{�
��<���_AԶ7��3�99�v����xz�ple������6
��2�]��7!��_A@j�U-�Q��w���;�U����(�í�d�zSK�X��ʫ�s�{��_N��	���c?�
�Uu��Y!_���,p�� s�,$��(�˻���D!/�r5f5Y(Y<y�T��γ���K@v�5A� MoCǊ/:����A^��j�ܜ!F8�����&����C<y�E���A^&�]�p+�0��b����Q^��Ɗ���Ղ���3��H�����hI�"�y�z��#F�����4nӮ�D�AKe<�h���4f��6��㼍��-���D�U�ĥ���������w?i��k�oe����E��C���!��LI���u�>�o�$�@�����@��e��^Ȟ��ZY�K}!O�z!�2A��y�W�3����u�5��i�C��^O��i�s'ݶ�m,"�'ݵy2K8���<���S��X�8�z��RU=�W�&��u���g!��h����R�C��4	�~�&���XuG��(�� 0���[4���Ǯ9�a�S�1�B{���>�.��n
��i˶!r��wD^d�	�2�X!�qN�w��:;�
g�լ�(3y	���d��c�x�1��#�������AƧ�oz��WG)kLdt�rQ�� �З�"��V��A�x�d,\�@�2G���W���"��/��ސ��c�P��~�媃��Bh�6~� ��92ƳW�[��X���T6ע��������1#<�vGO�1AO7f0b�9���aB�a��pVϜu��ٞZ�'龽 �ҐH}�T�d�����\*�K{�N^-��/�'����H}�c�-A�`h9#�N+��ڪ�/8�F��/��y.Hc�&k���#�� o�("8�C��RT>CC�����x��y�m���<��&��}�jng���k�S /����x�Ä�8?a��/F��\�Qk�G��{qn�}ػfr7>��a#�5��s�{#��Ʒ��w����;m]�~�%���<�NK�Kd��������<=y,�{ܱ�黋e��ք4o�#��b���fI���e<~7{�-��kph��82uNZ���V�����P{=)N
��p�j�����At��������,����V�����c7̼��#��Ἓ�v=����d������VOl��?r'�FڄI�3��##`:r]�K�[wZ�c�	W�<�*��ţȢ�j�qK��C�/�bϚU�k��z�8�o�Б&�䃶1۩|:���E�E���Ck��BB��jH�e#	|�.z�d�]��v�O��+3�4��b3GhF9���%�dF�*he�7-B���>o����xf�	���b���^��o}
'���O�0*݅�j*?��hj�:5����I�J�G̾����[xs�<��G�ͱ��axy�^l��n2�kw�o�/��q�c��;�MM��N��%�Y��,~|Q��8��r���[�5�CA��EB^ÿ���/��#�:�F~(4#S�f��F*�L�G *�,S���6��x�d��r>�,8*�.︕���=P�<��m�������V���7�~��J�'�'ﰅ5� �[^�,Բ�@��'��
o��yy"�}+�c-觇r�)�~�3��V��G��[a]�+" ���r!c�"5��p��ɖ����qv�!AD��*�L�]?��,�7�f�	��r��P�'���wG�C���0�H%�R� O��Hy�2�ع�I��\�PG5Y ��P�\��D��� �� ��uK#Ȉ�HERd"���ԙ����׍ɻVȓ���=�o
�;�X��(��ԛ�#���L�H��e�&C����WQ�Nuk�<��E��C�?t��<�N!/�������n6���X�j񓜯��y��~��y!� y� �]E/�f�}��#y�(D�f�pp8�AΏ5s�A��4R�,���w�'^EsA��&WW��&�e� }���4B� ^&˳@���'c�Y/��0Uk��Ȥ��!�Էv�?�a�w�!���I=;�E;�8� I��/��qy/lSS���.�$>��-`Oэ�k��BܖAc M��������ī�┑�8�`���Z�6� %K]n� ���c���P�U��"�������V�G� ���b��FC���xu�H��I u�/A�N����c*���p��/�SW��#��
d}O^ ���I�p�����8yeQi�),S���k�<y�����w3�ٖ�Qr�7
�"�.sd�Fts�HCn�8�!/��.�)ile��'(﹕�t���>ګ My��B��U�D���>G��d�S�*X�;yߟ-�p��'d`�ҵ�Y�g���B��8�hBx,�Ǒ�j#bV>��>��UO�nАy�;��c��~�f|�<�pw�{�G;7|O����;��
���l�t���_-y�m!^=|�|�ʹ?n���^�A��fnx���Y�}Ͼ��ovB�ʸDT&��$.�q1�JH@md�b�	:�����|��^�(�p�����t>8��;�6��g�˼�8C:f����['�}����p��'M]h�����>�-�Y�g�=q��Y��̸��TԘ=�y�+��[��D{�!}�,d���,'?�L���?N�=��� O&^$EG#�����*Ү�N�g�)k���;�=�eF!���GL=�-�tbNd%O_��3jL�Qi�}=�t��1sriqe��4�T�WF��������L�������6
/ݩ�m�6x���y������W^G�p�%g�s��h
�C��(����%��C������.d~�;
w�B�YpFPZ	T����i��>�:O��7�����xz�9��?���6|�bF:��v"`10rUc��i5]�,	y��o��&
�`�z����w�z�ʿ����NT��A��%(5�t�@6�3�����)��"�R��ʻ�Dy��5O2a�|���z�7RH�4Vd�Eº'���y�e)��4�!5&��Y*���5�_x	��}��k�	�e��y�Ԁ}��6����~�Pd1yO0ݪ�=Zċ�׊Z����H� U�jd~��{mƲBMҾא@�FH�7HAU\�����e�z�4
���l�QH8��s����z O���� )����� �O��iǣ����83c1.PyĳQ�����6�zʍ���L�d������{=y)7P]����2c/����F�1T��Jc"�e:�M�l)omG�0�d����y�7)��� �,�������w��G)O^� ��E�ȫ�`9�mPM ��.��?I�z�$m7Y�b�/��LG�4Hy�d&mu����� ^(�J0�c���Ё����Y`7�RYV�y�����ESq�
�WW�<���T!��w�?Ƀlwz
��Z �R�3V" �����H'ַG��;B�'q�䥖P�@���4�ĩ7�yLDM�oG�qΞ�&!�p�=�g�&5�D�@8uE�`#����4W�N[w6^V8;Jf�Z"daj$!ˌ��3��MJ6�DA� ����Nt���a;:df���m�S2i#2����S���4K�U��~�y%K���v�9N5f�DУ��O�����C���<yŕu�Y�	�ro]~])hg$S�Q���̾�G�X.C�]~��L�e��/�g��x7��ćL��<%ة�y2�V��g��}�c�iț����B���ɣ��@��\]5HA#ׇ��"�V!i��k�o�ߘ/����%B���L��t�x�'.T�wn�
�\�Q�E��1�~�� rV<�ơC�_ OΉ?��=�/���'�q�n��	z��i!�>��D~�Ҋ�=��]=��y���?����]����O#���ڠ�b�U1�Jh	f�*Ogf>ڲsѝ����q��D��u���0��'���78u�3�;}%~��. ��wJK��;ȶ]�j�Z:���c�������c�#��,�|��y�쎓��
�½|���_��L�pG��G������c�0	9��"�w*4��U�m������� �t/�~�	G�[�V����gh�ǌ4A=������X`��x�D��dY�n����v_������dad�<���k�J,d>O��R"3ƶ�c���x�@��I���{q���"=�P\���}��E�!�}6�X���.ZV?2N�{�gS?�j=?Z��n�y�X���}���hZi�T0h �~�_�=u���Go�ǖa���x����7���!6(0�A�9���B�^��%Zh݊4S�y�]ȫs���g�d�!��KȫkiG}h"bV��l"r�ܑnh��(V"�:�8o�z=R���j�l�t���|8,��2M��>҂qtG��Ĭ���3�GY_�K��l��उ-�}o�ô�d�0���)�|���͓ٙj\�M�Ԥ���L�g1Q��
�
IP��]M���Y�*n܊�@,檰T�9i	>���	���01>���F �:=$�#(�G�.5�M$��He�2���[	��n@����AP~`��4�X�$n��Ճ���j���ma��p|s�f�� �hT��d����� ��)"�:����dl�t�j���r%O�D�q�]�H��H�R�k�{Tuo�].h�O��;�ȧ?ǅ��(���7j!/�V1A��r�H��v��@��|�07ك��7d$��B�`K\����O�-2S�O��SI�@�@�_ŏՖ���[��/�| �َ�u����[�J�!���᷎���#��w�V}��}$�0Q���M�O��ܷ�a�}�s�U3'�\���
�����Q��DMQ�2���1@��� /e�%"�cN�a`]���
#H�FO��[����P�W��bۧ�3XE���TIJ���|���x�ة&^�y����B^� �uD4��A�0��X_#��"h��:�76Z��cKUW��l5�Fuww����>���,����hj�qß�/���ZyG2���v��z�Z!�#�,���a�@sۋ �#h�f�)�Fśbl���EY� đ��wіY�*&�.��z^�~���zu�����#�f���1��M�=�j-?+�X�#�p�5�Iu�&٪�^(��W�\eیF��d$N\�tBM��W��4����X���~Hd^�c�(+�pQk��r����8>n6�v1B'-B��%��Gg�@�҇ԛ��'݃}S6�`�f4��y�	�p2
?.z
_:��/����?�=��F��.��i'��e��d;e�I�Ud7��I� l7��g>�q�����N�8#����C6��(:��k_E٪�Y�R��1�B������?�	��"���X����N��tD�؇}<��=�c'�r��끳�]���Nu��qS]�y����W�J�1����e#�+ ����Ui�{!�8�� {G�ثw�F�x ����H��G��xd���L�j�$�18����$��k�<���)�<�x�����#����1Bw��)M����&5w��J7�������<�&E��B��"x���6&���V��4�D��df��D*��G��v5���f6��ع��s���'Qt<������G�}�!~�J5��﷚b�u��������]�7��N���!x��@�P��n$@�i�W�ɂ58����]��Yz�-<c녵w�V}3<=���돷n�������T���0�3�����TI+O���y��x�#<P�0�^"\��k�k�����*h
���j]&y��y��6���G�o �i�f�n�l�A��#U�m���Z'�ߥ����Ůs}��yuL���<$L�ɷ��v��z���v�QM������.DHp-�Җ�J)����P����]����$4hH��7��J�~o��r��2���ݙ`R��#�@��ٸj�	�4���L���xe-�����}v�{��Ĥ+b�B32�yRXy��᜿yl1�A�"6�z~�Y��8<�s���Y�o�h�Ԏ*�_tRȓ�t��M[�S��ت��a��1�!����A�C�!�?����h��Lť�k����ې�pǐ�F��"�'UVR룒p�$g��ޣ�"�P,!�[���9�ތ��q�=p�����Ŏ��J-xx�v|�M��Cy옹H� y�ZH'a7!!4��rt��i]qy�kȻ�YSw⤪'�	���k"�&	q��uAp���˶��(��(^��7PJ qIѐ��.��Ņ����[Q[M���U�; ��fX��Ǩ]|�f����� �<>]��V
yr�T.����˦��3�W^��Du?	B	8J��˨.-qh߆���r�l+;��&@py��n.��sQH�bJ���Z�
��6(�t@���4��V�C�<�|�Y��!�m`+Vbip��ע�L��.�C�lz"c�:��*A��{x��&bT6J\N�d��^�ΞP��MCt����9�8�7����4,�^v|E�p�lƛ8!F�
��[��1��� ��4O����� �.�Ou���5���� �P2�$ʬ��r'Th��T�	����ȑD}2AK��-�I�m�(��=���6]qþ'��"þ;"=���S�߬#��(�&��G%��u�,�n�"�N0���|�4̵��Щ|;}��ރ��D���_��!� �)0
I�~�9�ϊ'�A뿃���<۬�m���a�@޻@=}F*�>��1Sgz�n�o��_��ړW����x���M'P4q�{�B�뷈2��N����
N�V��a�П�����U����|�"���(X��|c�O��ߺ�L��Gz|�}�g�% �O
�x�(g�a�?���|�dŇ/�[>����x���cG�!�v���e\{�[�
���p�d�D[gd�z
�Ɏ�K��M��Ȱ눰	�Es3x[�	y|����߹� ��Aud0���*��G�
&ŔƎ~�6]�=gȣ�/Ͳ0��D��Q(X�ӉPe$�I��n���5`�{�6�u��Q�8D�xvs%�T5�:[/l�|.o�J��.�� ԍ߂�.��W�
���ba,'��FE�u�3tͰ�f�K���HQif:G^��E�ԙ����F�Zʋ}~��~��U;�+�ؔ���s_�A3�����z�Ц�Q��%�:���yGph���zx��O�g( �^�
�4��H9�r�--}]��?t�yҌ���<Yz�Z���E��J;�J���H7����_����5|�Մo��&�c������rԬ��CJT��5<�c�I�g��k�����ey�
Q�{�n*X�o��㦠j�f�L�����z3�Vj¢�&�e��G}�R��ߎ�r�׽x�,���9�A��XI�7Ӌ�b�h���Y��gg��n�����|�0���6Qn�<ea5�iN`ׂ��n������ �`���s𲨬Q~�qy3<��{�E����2d|5
r���yȢ	J�g$�dK�˵���5��۲-��fR�HV�Ef��Ş<�8o�
y�x ����E��@�t��lE LДG΀ǏoC/��Q��ళ�ec$�}����5�>?�ɕD���?��0QW����(;~B}5�m�U�p%3�4�GlkuĴ�FA�{�N	k��p�w0�1�%������ ��y=\$0�݇�ԬUxv�AEz�w�H��{��M#�� ^����{������|�{��6��8�[It+]�!\�A��� "I�i�� �w�oPNz�����%B���^��|Ё94�/��G@e� �?.��ߍA�IgԴ�D��9JU�P�a.��o�>����x�l��H:;��"�$7L�R���}{��vb�,Y��K	h��~�VÏ$�Qnc����.E"��O�&�Nd�t�L��F���JTLEX�$�>���e�����H$�J%���Pk���_E���(�^Ho|
�qٱ3u����r��9��-��(%�̣1�@�\������,Wׁ ��Z&�2�D>�[��5��;jpJm;�F����7�\N�y����@@���4����}�?�I;N!�}82u�#Z��ʚ8�c,,�I�s�����~]�� ���!}�Gh��<p2�DN�oө?�|>�����*�	�q��y�`�W����w�c�) ﰽ;vH�q�� ��6}-��!Gl�3Ɖبc$j4��X���s�KW����3Q?kʾ��P��d�]4��"n�K�����~53��6����q�N��4�!=�1�n⎃4����ſ.��I��m��;�ˣ& ���𣱟����M�L9G��K��6����y#G\6unV8:�=��>?��X
���z�� �/��!1G��#�\�Dg8u@
_�}G:w�}�^�w��!?J-y�	V���Gv�\[{u4}��j"C3e��8��a*�Hӷ�3�^�u7���K�&�A����>#yN�H�#a�{�d�Ǐ샎ݓ4X��5F��m%�1K��	�6Q�(�@�e�i���ݭ��1�9�D#lj��e�zX�e��F�ch�����iD��`6�,�[M�@� 34t1]Si�i�c��V)�cn3%Lk���4�o�3
/����cp|�o�F�ſ1�>?]N��;!ږR�[���{�uP�g* ﹆��,���
w�M	��B�wm�D�$�������W}V%B��P�����ə"���������9b0�t�my3mqr4�I;Tܕ��P�R�n�4�D뾈7/s?�?x,������y�W�!���8�v�#�N�e�%��?Y��kW#�sgy������Aǅ���a�p�!�Cg�#�buK��\I��yN �J���s�
�M��	���bl=����o�b�P/l�W��Iʛ��e2�yR�SE&A� �&
ȓ3@��3(,���Q%H�'^�|*�
������� ت;�	49��"�`i��7�l��(R���~9�F��F�
��䱥�����NF��O�n�)bĦ6k'�� ��Y����6��y��ᩄ[%-�k��j��x����o ��O2�(}�����O�;��)�Z�#�&lŻJ`�V�X���t�Oe�FWdiE�V�5�h��M�yټ+Ny}�S����L�|�Gd���<0s��#A޵�4(P����wY��9�GX�V5A./���ķ�G����t�V<�g��~���Wq��@D��V��X�����Z���\��?�R��^� t��(6����8�h�ZD�⓿�m4	�	�h��'	�"F �m+ /\]",~y���P�t/P��ݾ�;��'y4�~YG��Q�b4*�$��n�K����b73y�6]�B�Y9V��2sG&_���$�(4�|��ͺ"فÚ�nsߗ�O�<�<}��Ƃ䥇Ph;7<�ۛU}��������OE����r%v�����sݺ��=P��+dv��E{�;uR�k#��&��|J_{oⷩ�e���Σ���	���8ib����z�۽�]?���{'�h�Gp��g��G��C������v$�G������Z.^�سA���D�v��V^b���]�4������z��
�	�6��Kw�L�����ҵ/,����N$������舳-uq���`7��S�4$���{M����
�����Ԕ^3�1sk�0��1b��J:8L���-�p�q 2o��\#�������1����iBq���Q��?��ӓ8ኅ;���	��e��k�,�g�rD~�16N"�[�")_��v"�Y��2�8�E��'
���Ky~y�y�����Y�"x��8�9q��#����y�~C��xi�ϭ:��� beg�y|Ђ��}*�5�g�	
M=Pg�qj�X��
�"�;�~c�����s���g�m�L^�0�8�� K	P�V�
u,���G4>]���f�
�����Y�C��@� 5��/�yD���hjc��6���b��X�SH���Ai{��(�~�(�!�%a�O����W�.'E����((!��	u��	������O�񅖭���Jq������۠�[V_ w�"�����7y�~'-����L����(A�ِ���xz�r~
��Ƣ����b�i�k4��� �!�ĆPjLW�D�����7�"�(�3���!�����������'��Qk�5��
�L�[��m�ݑ�%)�{�i���&��86�L8F� ��ڸ�BS�vJv�
8J��i������)M��R͏N��!ñ��'6~�y�v$�놫�;#H[W�!xȡ�b�Y��y�$N�7�Ѭ��]�6��ˇ��{�8����Ps5�;��@}v5k䲕��K�<��5Smu!�Մd�f�"������$y;d�-^0�	y<����}I���-�,�;����^Hk�����Ȭ��2=�{�o����Ӹ|zT���!NI~4����y�K�!�a���_y�<9j�M�F�J����i�i!�yW?c��GM\�)�!OK@�ESO���'�.Ó*������,�z�3��7u��5�pŴ'�5�ũZv�����4�!Y4�e�6���=��L�˥�*�S�a4�%��V1C��%��<��x���%(��|'䱰n�Q}u�=���{�kƣoN"���"O�hc�kJf���M���p��1l�4+��&�ɾ��/Y��-"tl����5F� ���4�����!&ꏗ9?��sR�TO�f�!�i�4�Z���9��2PDP) � 3��)x4�d��"�ƑlG����SH�E7$�}�{�P���˵��$������߃b�a��y9�fHѶ��x���w@!M�򲍭P@�>��+�1�_X�#ǥ'ݾ����F�\Y;�W���F���4����R�7v�8�@�N��c�=���c��H�/p��w83`�8Lp��P��G��_��H�j����S���O73>�w:����n�opк3�q!Ȳ�~3=�=��k���~*7��\GM�p����Nu�~��_~F��Tv43̪����ht�i'�6�� m�:A������������k���Q+{�7��>]S!�-p��Z��`�Ց`7��T��-�!~� 1�g�(?��]�	��b�#{"ც��5�_��܅�<v�̖<��X/�z���3�O��ٹ��z�消'�ek��2ܐ�D���7����E@��ԔO�<~dK޽{w��i=���CuX �'�G���tmC�c���ҡ��z�S��G��B^㒭���FRa��5$@4�|]7�k��Eʦ�D��3��	�j���U#c�
��vƞ�8�l����X%1�R���z&��c��Z����l]#y�k`��f)�a��kK0WM�Q�I41_U3��kK��W�b]�a��M1��g�,"�u/�r��!��X�e�?	&��l��
�H5�G��' qV��Z�x�a��4�|�f*�"���Z]k<Sw�-ۯP<� �7����w��c�+*��a��)�&Eb�rmc�����?���yd�+�J(!�ͧG�Tth�PG8}.�SO��{[7�鑣h� T�2�N�Ry��Iy��#��#�x�ma�:���͸�gN��#�f�w�頪�6*[렜`��fY8\�D��F7h@fȋ������ѵ>�dJ����-E�)����7�?v��YC��twA��~F��X�<�LJ�т���RȋWs��I�����磗O��^�_6�����Ҷ�<>X!�x$�����F�hN %D
y��K@�/����<.E����r��+2�{"��&��J�����']�}y���֔���4PgiY FQ�����kIW���Y5x�����y��e�x�{���W���#���� Ϸ�:�Py��B0M�[�#��."��!��n	�x�������pABE���={-���Od���F��f+�l��!O�MQ1D��!R�	���5�� �������p��>�x�*/�F*["M���]��$ <w��Dε
T\7䱰^��^��:�u*V._��J��ň�'
xn	���q]�JX��I:�z瘶q�UM��NY؊�ȡ:6#]ơ$�͐,q�A޵e{��������Q|�;N�d����q��!j;��k�Wy��8�ƛ;O$�:���YxlE+���� �%߬3b-��l��k��5�e�_@/9s�|q�"g�˵w�_/���xŐǱL���n�]�%/�t��<J��P`�&�,��Hr�
�����[>9�+��<�G�٫�1�]��kW졉�|#,utǶ�_�ܨ?�?yBg/B��MH\�ɫ�"q�f�O[��)�������mߎA&G�X�'����%bN�cg���t�!�.�؅�>آ���K&{�ͱ�走�=4���w�2	�펚`�����I_d��F�p��Nș┉� �}&8hi��F�J������a����#�v� �	�yyv���-v�[b'�=���rv��{�4Wl�������I����H�Z��1�{>�m�
o��&����qS�]MD͠v��������8�4q�@�[��_k����8��8"���v�<���_A^CRҧA��dm%�*����Ǐ�P{_�Vd�p��bd�0*�t�D�{O��A^G���7y�l���ZyN�Nٲ厅?ǧr���ƽp�3}�j��:�XF�� P~�LCɴ�8n�	kII.T7�b��uT�sU�D�TX�؉�mC��3&��'r'�W�$-LQ��Lm#�Փ��e��ں����y���ZF����I4�O�Ң<�b=���?�;1뷐�~�Ґ,��S%XD�:CE3Z*ሚ	�YwD;L�N]O�喙4��@�㧤���R����4�����C��zYW���>�:����v4��#�`���x~�$r����)���9��,dc�P��];�,.^�<`ӒT�6H�,w2����������<����v�|�M��e7W4܋�;���٤�+^���+����iLV��!�\�Z@���O��7�&����<H.is�p,����?Q'��G��*�Ho�Nă}}��`�i�^�7 �80�E+۠��x�[,Qp�~�Q��b��my��埁c#�#���qU�@XSd��<^��]Z�F��͖Z��L������#А�/�ݱ�faE�i�'M|�nd1<����Q\3��Ԓ�jo 	/�JE9�Ⱦ�R����@
�T��!��k!V]Y����_�؏��t�g���� ���z����pV�;���#�SDD[�9m�R9]n�?ސ6z$h~S�tm �鬲��:�Ǘ�0g^ܦVL�ϗ���J��P����r��w�Ix��ti9)�|#[^<*�*�䵣�n#��bh?�0};D�� M�f�Fݑ<t6�|�=C^u5J+�z�M�{SX�߻s��Kj-{����2�����ȫjg.8)�$�P@���}�E��H�4�ik������,���@�Ӻ�H6w��9cTQ��ͳa�:�'$�c�I��z�ڊB�/Q��r5{T8���Y�uD�r����#M6h�N'�E�Ub���0wP�c�x�~��p�Uw�z@챓B� ����g�3�LR�y�#qO�M��Q@ �K�x ��uF��&�4��[#�@!�ʋ!�����]P��E^���:�fmnԊ�n�B(���7N>�X�ݭ�#�TF% p�V�9kF��3}��^DZ�?R����ԄH�'�Va�S2P����q;��^�̙�P���@}q炱��?���K�'�\��^��cf-]:m�}&iVb���X��&p[���'����l2���ON����Q� ��̄�n�&�[�L���[���01�v#	vJ̅3�&��C��n��{��S���ǽ�~f�2�3���S�G��1�u9J̘�O���O� Mٟ��M-	�L�E|�s�a.��I��݇/�n�3MP��;
p��Ԫ��jK	v��آǖ��L�y��]Eċy2*,�7o���\B�_ޡ���o�3K<v�8w�Kw�<�wxoB����c#����0�� @=���� ��DB[,m���jV���W�n"L�d�h����Y'����X`b�YT��l�D�RX���b����K;EI��0Q^�����(j`��&&���0��A���=�aA�dm}L��=NS�u�1M���O`2�
8��yQ���`�m'L���r=LV��!�}Ǯ#`N�E��&;B��SR@�!�.��L�w��E��5�X	��G�{L�":�݇�k�w�N�-.�� ���@��E�����i@1�B�E\9�S�����'��'���v�9eH�KEvQ�>�;��f�R 2K޽��u��v��L�^W:��r�Jd,^�S�]D�"��1a�$fE+M�6U��	&
�����:
�����q�<�����Li�`FĢ��'a��5ǿ��I�����׌�IS%-�	�ڋC2�!�(�2ȓ-��5W�wcUlq}�"��+��	��#y�S�1�<B�����,�ۅ������*"�>[��^�Mm.��!��*��F���6:k.A\�Q����Tl���sϥ�oO�#��eH�<q-���\�MZ��Xd�7�I3�HoC�َ�A�,��$�'y�?G�����j�H�J2*�
�n�@҄]8����A���v�Jy�o�!�uaP��u�x$!����+�<��s��89u	�TK��ZY���Q,���C����B����<��Si�b�vu�H�OR0��,g��V�bO�?M.}�M�g�hX2T�o��C�@T���M��U\�.�8�{��.=޸}G�c/ꞡ> �]�u��S��ܦ9,^��Iy�llq��^��<�Y!X��:&��{�솬��q7���5�,>��xR������K�,ڃ�oP���R5;�0rA�����r��i�����0�u8���4��3�L���G�g�צ�*k����B��7Aj�)����a�c���$V��ǱK��`�@��ȹ�_!��)}��+����k?�vH�� �Y��5��<)|!�Ϋ�(�( 8@ǿ��{�-�q��j��ܢ9�C�\�E^^�������x�$�?�
|C.�l�y!!1!���FaY	�JJP�����$D�\	,�K��>��5p"��}���� o��=��1��&�����v�D��7�B�H_����S<;��/Fᤚ5��`��vZ�b��1�b�M�f�@������N�JvDn34%��[j�4A�Kc7[�v�Z�zβ��G�m��Xیp��
'̱K��������;��]�����-�j��_��7��e;��0�1���mq�X��{��s'�٢��*|�q�M>|�F��j�,+W��y���=K&�������J\/)Ey�/b�MF�������[�sg��@3��fu��.d�'���<�+;!���"R�_i��LJ�{��c6)��ݱ��1�]G��u�ä�����
k^VYb���/�6�e-L�S�y��^��)�W!�(�a$���WP�xUuLV��tMma���i��Z���G �����z�fd��S�$�\��<�N!�z�9K0Q�@���@�9��u
��|	�����'��6�=���o�=o%�	�x��HO�^"7���5'��u��h�����:ûW�vt�Iw�%��� ��N��S>�����9�+G�����ػnΝ=��n�>�?���#����^px�;�Y��N�a�J8b�q����D��8L����'�r�0��Z�Ne-TQN s�-_;-z|�"�|��@�)!b5ޏ��&�:ɔ&+)>fWs0�� u���շ+Ͳ�E��b��&-��L�6�MK��PC�#`�/Cޛ��gy�b �$K+I���Ǥ��^��lD�ٍ��qQ^SX�d��J�bI!ؔA�K
剅㶲d�U��#Z�!��H��6"�.��]����^*�LZ|��%�l���t���H�:Io����'HY8�
�2Ko���p%xŴWG0I��.�hF���Ap?����c�v,o�|_��x�Ո�Q��إ�T�Hp�VT�D�V_H@���Uʣ?[�:�(iJ!O�G=��Ĕ���[*.�����*�Lԗ_G樥V�(�3�d똢Ȝ�i��ss�+w2	��Ҟ ���p�r���Y�Glɋ&@LU�G�qg������h�{���v���@�m�~�JxO�HF�w�H!�:h݅P�.�!�A^	[�ހ<)�h�!M�'p�h�B��gȋ�4D$��E��Ȟ��S�q��ܯ�#�<~��0Mw��Se>*VE�=hkG`\����g��n�/��M�a�if�ȡ��*ʏl!�3�E����n��퍪�y�j(?ܚ��r�L�o<�j��pK�KD��Q�rR1�Ǟ�\:����#�����<C^����"�(�4 �6P0j1�
+�aΙL�
y��'�x�72!'N_±�gp��I�^���Gp|�>\9q�$A��#��/���"��
���".<
��aH��CFb<����$�����?�<�LZP��0���VKw�$��ne�Mx�M��ʌe7������Ǩ�/U6��!���k@B)�������&�[������,ͱ_b����A�m4	�J�.?�){hB"ޣ��K��/pA�v#lё�ۥk�=Tw�h<�%���mG��pR��������^��D��8d�~���{�b� �8\0����cn�0'�:�#��-��.��C�}G1a��'��y��¢cm�xK[$Z�#٦r��[�^����?ŋ��������� y~:e5^a��S�N�x�L�G����*��ֱ�;��*�X���*�-yB�H؂�Ҡ������;�w���1V���\��������ըc��<��̱��|C	f�������c/"�K�˭S�1��"~m��_��1LY�+��kEU|��K�����i�'zE�7NW��7����-=x�t����B,�e�/L���Xum�����?����<�K���#0I���Lc���Ѐ�G��>Ecg<!E(�<i�[>xq�f�4�P�4 ������<��ED&a�Թ�6o	�L�k֬­�l�;�S�é�#p���^��iHHIŸ��1i�l�Z�K����a�)X=y!6�]������O�<��a�?�/�+��! /����� IE�tA�♸0i2�v#�3@~#�6B^E+u�	�k�QE ]�NU-4�Gm!�s�I�GO׊Ԩ49o�H�>���qs�e0�0�NHp� WW�IDȭ��M�-�i[��A����q8/��5�9����{�l��?�7B^� VrL�51��}W%O_"�dN}3I]�F��s�S�v,�M�&[B!�㶲d��@���T���8���9J(ja��D�cG�|�T��a9u���������=�o���,y�y$�rZb��!/�����N�N�s�
};Oi`yʖY�c)�1X�p��/�֤�|���a�ԻȻܢ=�Z���m�+���Q��#�͓��6Z��F>r�y�8G
���Nt��sW������x��,� ��˧��<e�*{"S�R�_���ce���Pb	���KR{=�7�>�.��㔚>��%"T-��L:ظ��b�ib@����p��>�cߧ�o����n�SGD|�	���}꺣B��K���%��@�T�D@��;oO�Dg�f��7�ky�^��Ι��߂��Bjj�QS{[X��,��%�º̐GZ��4���!�������ho�7v�A-C���4S��Z��5�P�mb/ /޾�g��/8/�����G���5�ѨR h�<e��S�L��i� '�]����g�L=K!���H#��!��ӑ	���s�l��qc�z<`����"o���%䱃����8�m��b+M�ϟ8����a���8�}��A�E�_B�y�}� ����ƅSgp��%��8~�N\ē�H�Y�ϐ���:'32~���_a��;v m!x�(!�2s �s�v����&.�A<��ʌ�l��z�ōK!4�<ǝŇ�c? �j����X��ae�ff�O�w��E��K߆đ��[�Ml�I�Z#;l�p�*�;��4!XI����s��#6[b��	�iKp��'����O�Q����q-	Ι;�(}o��n�#k�	�ܸ�]=���E'Ěu�Uk����3+��8ⲕ�X�e7*�v9�Y��;�<{�%[xv�c���T�lga�X��D�K���:�dʥ����i�<V|��ƍ�����jd��!��Ϝ� ����8"�H6�������p!��{�@�!M	�H�s*���kN�r��=^��kV]Dȗe�Z��c����q3>c�>d
Nh;c��.a/�1���h&����-LS�K�3Tt1Y� ���Я���L��0��v¢_�����ϱ�1�'qsCOM-�$1Ǐ�Z�MCS��1IU�icU�,m3�ԑ�\=3����J�dl��u;i�{��#�0��	u�D�����H�F�̲�PK0[�eH����7��q]�Eν�=1�j4x�ng�2�X�����������8zr�m߀SGN!.0Q���s�0�>�� _���ާ���A�ٳ�����qS�h�8l�9'7���c��H���:�_8��E���yfK���JFBǟ���
7� IQ�:�!d�|\�>\{!�wE%q��� �Zm�L��8���a�n5���B��_��(�돗�Li6�7��nn���V�����^=�ۻN��"�`>�ID5��-�_E�H�L	�M���k����\���&��D�X�b�\<+(���8e�GޗdJ]�O盡�P�?�,�!L�QD@`tl�K ��oA�DA
w�ּx~�!ؚ����Oq���*J-�����|K��cp'M�.�^��s��v-$n���E8�Ml�9�u�~u�	�
-k�jY���M��1ҩ_fQ�Ƞ~�BJ�O����L�i���O���Bq�Rȣ�
Pb�����9��݊]�إ�����G(�{,�ǟ�"����6������RA 	?�k���r8G�9�8�h�!8�`5jʫS�һEV����.S��[WQ���+pQ�#rT섏��v�Zє/.C�F�
:�ѷ�
��y}\�v@�D�S�I'�X��_��PH3xj3�d8q��۷o�;��2��w���2��"p���֜B��0Ty��7��i�Z�
��vª�m���l�(��r('?	�*�#� /M�	�pɲ��DeJ6�����������.Ko�7Qv��X�|N7� �t�i�|�j9w䷷D.�PQ2!���L��9�L�f�t3�A᪄}�eS�9"϶�m{�z�zj �����D%'�K��DRagm9�\�Q���tjce��H:�]C���TW���6Y/�4fDZ;#����(v�$����_)�%�p���	��W�ߏ��Դ,�8v;��ǁ�{�k�V,_��V�Ǒ�;pz���<Ac�!ݵg$ُ�{v�♓���+�'q��)l:}i��㹝�yBo�U�Ą�Xi7���b'�!T&��fn����n��L]����$��cfI�1cqҢ�41i�������ε��Zj���%�]�l66�==����6=�{i,^G�7�&�3���Xb����c0M��D���#�Xt�sl"8߬f����;tLŖ��T��u�p�&:��k�u��s/<
���}��-;pޥ?M������=.�w�����w�~ߏ �Ü�2m0�{�u!a��h�H3'!�N"RU2��<[TY�#��A�GH]��/�+�<>~�3��!/�1��>���.Q�$�I:e��E
y�R�Q�� ���"a��';]��^c��y�M܅�yr����#�'g#k�^\��=m�1�
{&u��,�<,#c`�qj��NY��g��4�E3�\�}�B���$��3qP����Rq���/�D���AK?*��t�1��M%X�Nל�j"d�q���m�K[%,��n%�yL:v;�t�0��*�(�cVSDS��ںG�h~W�Oh�{���D��5�{#s�"�^-����xs��;�?w��ގ���&�" 0������`l���@08%�9	�
�����0�?�|���4{VM[���Lp��?���.��}Ry׃���Қ���q
j�����k��b=�;tC��9����ZK�;��mE+�W�.8|VQS�ij�R%'{FC ;�}F
DZvLoA�L�ĝ�Wp��s\t�D�o��8a<�9� QIM� ��-�I�W�%�X�P�`���9�	��a��"�,�=/*&e�LX�8���j�ˋ&C�����N�b���1pn58^��9�w@^�g���Z�;��Kk=��qo�i�����W�1������g����R���L$����֮Hn����
���MՑFy��2G��%
I9��0	kl�a�K'h`�$���P�A�Y����bq��W�\c�|�s�=�C�Ƴء�pU#�6k/N����R��QE����x���MZ�#����(��<}�Cw0툃�����u�}�eDv�w���3:��s~���<�q�S��zd)ڈ�$im���^1Tw)y�'5��6b	�8rB*�U��>.�J�g-b�Fj� S�⍻�j��x�O3x�m��'=�/�<���&��R,��W��!��ky�NߣX�%��S3D��D,+�h�K!O�`3@��9:�5G�ĕ��A4�F�#I�Qڎ�`�9�:-�׫P|��5ը��e�$ʎn�!�@U<=�n;��oQ��E
�yfT�"�-C�'܈�ÀG�y�|�!�&,��z��'b�z��/��2�\ܶD}q��x����0}7{�)���
��T^y�(���3���ؤ�T�4Y��&�H��I��#ˡ�p�_��%�����,Ë��W�b�JoBޛz�C)6&[ir�e�nlX�k�.Ƣ��v�r"�[�x�O�����	#�c΄?�d�T,�;;6�Ù���}� v�߉%�"�����^y�m��-;�U���Ӳv;b��6�%� o3��F3gl��Y�o��4��En��>�u���@^9���C��7���`��)�[:K�6	}��p5�=�����U7�Ds�zb��#qz�\�ލ�}�v�"�����d�o�\�_)�`���S]�ӳ�zM	V�ญ�H7\��]4�o"��~���h�"a�R�f5�D'�П�`�>N����'��p��~tW	�8�m��=�M�q�`�!/�`NH#�E�䀅c!�p��Z�4�ɵq�ud:vBа�@� ��F�B`�c�c�A�5�"B=��ƌ�)'wR6��W�Hd�<��zvl��Z�d�ty��%u8^�}J�[��=�>3/�0t�ɖ������f����oxO-6�#�bm;c��A~!�Lm���󍬰����$�m@p����Vpi�
���1�W�'$��7*����|��O=��@���]d`�ؑh���z��@e�A%)�9ʍB$?O���'��b��ٸ(���뱐f�Z*bh�R�>u;w�S�E�U6C��	��1��r���r�Ȟ�\X�g�*�]���v��=L�s:�L���g� :*L(���\$��#>%���)-B՝��JFd�E�߰
����z~/k�@��*�haз?!#'��y�uv�2��� �&0��C�����z�QUåNnx�g�>�+�!W�՟Iݤ\#P�A�Na�c?y�ʹp�)8����>Ϡ�<%&z*���+%)=�!M/��n�~8f�I�G�*��.['$Р_�L���-A^K$,� /��^se�Qe�S��Ѵ��$���_$�^�"��F���xgbeY�������2p���`_V$p��f�-y	�5.��q|V9����FI���$5i'��&� �7|�ؓ$�^�ȓ)�#a���	Y-	@�j"��2�[*!����`��%֨|R�yZ�b�=���4�@p�V,���F���2錐�3�<�\\�9��@���M?w�`�q�QuE������OK5x���*�����0D0�ޥv*zR+�_[5���.���Nh[a��'���C����۔��ĻE־ބ<��c~����ه��ݑ��JD&a�{m��K�|�"� �%���8rZ�'h �D�'�Ç�ډ�6~=�T�N�VV���'
�LL�߰�	�c�	y���u�������u��'J�KP�B��j����)�K'3�g8��n����;�	УT��D�P����-����q=� E7�P^�q�W�<x ���$ʊ^[����J��/�~�փP��Y,ײ��T0�R���Bl&�*�Ҹ�b`/,{N�ᎣO�D�-��4������]�����t��,>G�\x��;��r�N"��)_N�4%K�9!����v��p@"�O�����Nݐj�tW�8x���/l?G�o��4�O	n_i�#��ޛz�C)!2����.���E��� ��e~<?}= �|�~�-����}{�����C�����#Ι�m�c��E�|97o�3[���d���Ie�9���_c�yg�  �db�-x;�	Ќ����a�Elж�^�l�.Y�e��cIw����8���i�‶-A�=�l�z�`hEPf�M��b=۟�Z�������������_������wk~��h��N��;`w��1O�B���M�sX�Nl����4Mp��u��K���E]L"p�⦭�q�<{#�����t��Lh�fb+��A���AH�5M��X"�\ނ<�%�MȻE�(��P����\L��.ޖ&�>|�*RoC^)���LD�>��c�;g�����0�,y���<��7!��Ώ�1k��Ii��	/-;	`;H�MQT�\�.ذ�ȴ�ێ�[?,�A��	S�O�����9/�N���B����M����%m�B��Tz��n�V�z�zl���=.�?����8�m5����UUL&B��e�E�,�Av��Ժ7_�Kh�0����_&�!!7���ե�6U�]Sqzw��"h�I��Rm͆Qcy�m*�_<RpF���O�WyO��7+�m�X�=y�EU������X�b�ۍ��l*�'�w�������1N�߃��h�7�/t�w����5k�6͚�i@����#�@ai�G� :�ܤ�1^,�Ra3�ew��6V�$pN���U;�.\�+� ��;
�-PMWE��59a�ca����٪���z�Q�CҀ�I��E�7nX�pz�$߄<悓�f�Ox�������ݖ�HV�Eq9��6H`Pj�)yIMŁ��ߜ��g,��$D�ۢr��(*�#����,�g���O��s+r�<��l�9g/D+���M��1�� ��.�  �C>h2D���>�(��*��Mj�+��w��qb�."�WW�D��7�.�%`I�S'gڐ�ppt�,t��(/��o\+uUa�ˤz�l����&�6���2�L\���o ��[s�Ty���8�� ��Z�|h��~�R���z�w��D��Ώ�ӿ��ۨ�4勽��>����{����_t��X�2�ӵ�_�`�!xku~�ر5C/�Ktuwl��ӵ��b�l��EC7��~3��� Q�Z@ޕ#��/� ��'��������ݻ�<���bT���Vtb~����(���;�vP�H��J@ڞ@��V��HD�`��l9K7tC����$�T2D��a:��'J�BMN��<�X]Q���k �㍰X��D�Q1�)j��4*Tn�B^IkGN;d��#C�H�Y�A�8�k`+��	*:���e�L���D���L;�l�J��VT����M}Z�� �\���縺y�TN�(R�GUv��p�02�eS���Y'���,���4hgY�#��y.ݑb�ţ�Ir>��#����<.N�lY�-̝��}	w[X��[�9�;�9����bٌIؼp6̟�+����w��i$��!4�kNE�������^0�=lx���3o7[���S�𡋭��y�Xo`���y��F��I��3�C���`C����j�UT����8c;�����u,�^��%��֘�b�i�qq�&ܯ�D��'���G��x��/���E��
�
�~Lm���ar耾Jz��g6�-i��u4�!]�K��y����*rV�+U��d*�Qy�
v{~�K�]ӥ�?��]p��\�����0>��GO���q���8��g�]�!ﶽ2l<4�' +���G"�����r	 ���=C^A^��<^�=��s�f8�e,.�У7�;uA�9�Ka�{}��U�/��5>iː�� ��r9X�mWkX`���/��%���r��[(.����{����M%J�bd�_���E�=<5��{�$�j����X�����N�G�ٵ7:�H,�F���c��C�ݾ�Z��'-a)dG�˩����4��Ƒ5�~��b�g/dQ�G�M\�a&Q#��JX�^�h�{A�Z�xBP�@ ���e'���E���uD(SoV����J���1�V^���l̝63gLŅ����'/"�J�/c�ڝ�?~��!={C�iK���	��4�-G��
5�#Ǡ����*�O��M6���^gȻ��ܞc���B \u�����`d|;
4�.��Zs-s�����8�!ID��6��l��tER��Or�Ӆ���P���+%�5�hn�5�'{��E�n���G;����RF�\�g�+�8���+�nAZ�}&'�*6(�}�r���A�܋��ĵ��~�>m e�)���={i�N�X��4��#��<����:x���O��N��Jt[�]K������B	Ҿ�S�����Bo�g^ႎ_uZ_��#� *�� �ISUтÖ��BUsЄ�-	Y�| ��J,���m-$�1���a3P#ݓ��ߒp޸5�?��3��UKOฆ.�iص��/7��-�(o��ڗ�|��C0���^�r:8Mpu� � �ҷ��a[�oqx�J�.��Py��w	�R�an��o�h2��͡ɲf�*�"���	���1/��cL-Y�!/����Y̖�F40�
R5@<As��'.�N�ǳW�s�c)̓,1H�b0܉%[z�,'ORP\$��#l�Jě�Ba;ki�jC�*\x�%.�#���%Yc;D�8� C�)j��R��6t�EI7��ڄ���W�w��T@[y�[�N\f� �^�/^zX�P)k�b5y\nů,y��1�I��R4-��m%�mI2%�(��@�C7��^�6u�������@�����'Ѭ��+�}#P��$�)�*Y���,���TF8tB�����ecg$X��!�4y(��@��#��i�����EF)���Z<�+�����]+��#�Oc��e���/�������X0����6-��3'c֟�p`�
D��B\�7��BP������ţ�Z:|��Q�{�?�<�Hqj1���
뜿����C�h��-�Kx���m���
k�4+�ac�Q4��.ҧO�3����g�MT�����z���z�Bv�9c��)f�ص̣+Bv�&�����u�"�+������dί���������k�ҵ���ج�/���6��m#����1�fyM��i��<�������$��7��U7/��s�{ں"΅��A
w�4��p���m�[7���I�ad#x+� /��I�.ȶ%�#�J�vGȐ4�(�0�q⛺S{OX��**��Q��<��7Z@����"x�=�^�w�, OjœB��fA��,��k����U�;���Il��Zz�<)��4\b�	����B�JC\�a�G�RE],4��S[�o��c�U��$��Ѷ�Z6Á�k��oN��־�,�N��d�Q���}��x���T��'��9g����h]]L#Yh`��*��E�6K���,0UC�,pn�zj�w�:#���`���)�cA��{dK^-)�'�.x`��T&7tܑi��s��8lһ+I&K�H�ܸ�i̂1pw���[+|��wX�b�L��YS�b��#�f�;	�;8�R[�ct�䎮�]��f3H�q�=����Wyb�"�<�R$8���p�W+o�*R�e*z�R���ߌA��L�#d�<v�Q�VG@?r�O~�R�����d�د� 2�E�2�}��^)�F�y�� ����6�fN��g�3��ϱ�U%�2,[��?k/�)�`NH3y$&�QBr+����g�HU{T������ɧ$��ӧO�in�Q��8���q���N.AG�K�o@[��[�	�c��bl�J�I��<�7U����Yi���^Y��GBm�3��b��	�P�Zj�\VK���%\]�*Jdq9I�iV��r&���!SQ�/:��P�>y�Ğ�ڧȝ�'U=qNN>�!�3�5eG��Җ����Ň`�rS�S�ql�3T�Gup@�
۬:bg�!8�h\��xiY�)�O��?�ǻ4�xy�!����v_d(;�Xr;=DSێj���6z� /� �%��ݺ�I�c�f��m� e}�*� R�A�0)�|��8���G���5B�[����lC�C�q/���.A
i+V0��2䌑G��-o�U�9#�<S�j;!U���y��(�H}g�1�䩫_A*�J_����������J�v��r���'@pD@ɖ�7!����jyѼ}F��4Ч�X!M��&��!��hܓ'�<����y,��"P����A+q0�H���%����<�����
$N(�t@��;�I�rԋ�^��� /�@@'Ѣ(k�y�8�Deq5�8����a��?0k�(,�;+�N��i�0s�(���X�ݻn)b��!�,��Gw���JЗ�|��͌GE�l$�	�NKOŎ�`����n��h<�`a�զ��`J�fl�y�`'�;tm��&�������}p��7vk�a��5k�L�ِ��c�u�kl1�`k�c�����Ghhh���"஁�="�<��)�M���X���`�M����Z-c,�S��7����cF�wDG�#_��{I@�-LZ���N��I,�^tqC@O��t�(G/D9wB�sg���y�EJ��H���C^	�$�C}7ˣR�h�������4����G*؏X�d�g�zת*PRZ$^��#��A����q��:�8Dps�*�Gw�9v.T@- ϐ �8♡�8Y*�<g4�H�$+/�ZvD�Q�#�@��]z���ux�}����ǭM�����x�o��3�[`��O^�͚��^]q��\t��Tq,�;1�K�|\��'U!�4����[i��S�oyF~�щ�5&�a����q��	fZc
=N���d#S�9	�3�p�D �8u�$Um�<U��o��Ɏ�r�4dZvF����{!˲�\��"�2���y���w����i�>�G���
GKSX�ؠO�~�0n�,���~G�>ݠ$��m����1�O�����Np�ߠ�8}�$6�ۈSG���j��J� Yބ<6�񾼇y�H���f=P�f-6r_� e<�ď��Ӥ�2T���N�X#H�I>�슣B�U�L��l�����Ը�I�^���JI�B�|>�Pm��jpe�5�CPsE�4@��-Zj�SP�.}�"@���=��%�V�Z�d�ڤ�8Y��ʱK�RXqd�Ə%����Fy�/sǄ&���y�����݄R(#���+IK��d�/� �O�ɣ�F7SF��5Ҿ�YfG"�J����e����0�)�&#��+"�C�U�'�� x���#���8���Fi�m�N�'����pP{�gh��O��<��Υ�U#�<я?��Ut�����qV�>4��м��=JSMR��?�_+�����E*������|[M#�9L�i��;�|9Vl��j���u�)b_�%��7�?�y�.����aYA�1���T%P���"v.���"�lX�	�)��J�8�f�+Z�Q7@"����=������<v9�LS�t��5����&����[\��%[�o�Qy|��@� O��t�!�-x�rF��a4�� ]�F���b#���qt�D#wy�WJO��T���B
yo�ç|��1��nȩE�됭�����l��$Td˵2�6��P-���m[�N��?Yf�`��%��ӫv�/!����(�|-/{ᷳ��䍃���C^.��>^6��za�,[SEzϪ�F����l���I���J?�������{�L��;���7ƌ�=[6`��!�a`O��e(���#�p��Vڱ�O�E��E��{#-�
�s�\���Ayf�	�q���dc��EXn3�-:@[gj��6w�j	�=_kh�=4�Z�m��l�<|��C���X��-����l"��l�MF�\.X�k�yj&ǱfgMǽ�k��<�k;*G�<꫼O�D���K'�h��K��#O�ۇ.

�kO JP�\]����������i;���n]c�t���'���Y�� �+�Z��׽3���Dd�u�D q�؇g� [w�v�����%��@��3"�i�bn�8+[��{ �kw$�y!��7ݺ!�ڏ��?�er�'@��#>�q��:)ʩ#2�E�8 ^� o��..��ڭ+;v�ƭ5#1"�ktx�L�^�؇ǖ=���
�ݬXR�s�f���ֶ���X�/�"~�q�w膍�)`�����K�Ki ^g�" o���j��Z�=u��A�5�S��'Oځ�7s�2�Ʉ�SX�4.�����������Τ��nE_C-�������l�ɪz��V<*��J�ώ�����l��b�G?i����-������m��y[�y��Mǀ�>�]�����l���(U��'d^ԣ�~�,/IWq��N�ƔG;3[�v V���aC����^��0��8qz3J����������IE��EH��ĭ*�+��\� �������R�+����G��=�t쑩��S֎(]��7ⰳ'�ԥ�<�q���VҨ	y,y�4��)� ��Ż� <��A�A����%� Y��F��O(�B;�]��~21'�SA��)Z��V�Ft;a��E�<y�^7m��k	Ћm� �k�X�Ghw@���ץ�W1p}(q��zA�Ƿ�� �b$�w�E��%�����qsS!/�-�Ki�������8u˧���-X�	C' բ��ʃ��$���O���a</���A �.��_i���UG5$�U5F$[��rZ)!���[��2�|5��o��d=�P�kY��so�<w#rx�����O���(	��v˯�<L�8פ9.�F`�#,z��5q��
��U�	��:>��#N��!�<B��O�P�ZZa��_���xRŖvٕ�#����X^&e�)�����r�L9�]8��	�m-��L�M�VHP1'�3ּH�P��iaw*���l{=��E �]sa�
����&9����I�>{�q�q�d˶,��*�w�L�R�[z��v���K�����ҔuP*[�mg$����8U��-� /����v�A2G�(�I}�U\1�A�u�J��J�K^][z,|��U�#]�,���3k���r��F���8t��b( 4��7_���=;9�%�mKG7�@4Y�&�TVY�z村h�9�'o�~yW
&o�!H\�܇��F�<���\��(�sqk�ڛP��#��AXi������dM�e1A˔��i����;"� /o�,܉N[58�-ÝL���N�/��U���H;|����&ề�돃1���1���8�o+B���ŞM�p�� Rb�p�<|����g?B�. ��O������x!�Vz�S|f�/6Zt�fSG�1�;�6���F�[C�8���C�HO��w��б�6]l��w�w�r�J������Q/���1�x�����'�Q�d��0����'=�A��G�&j�\�妆���.]���2ָ�b��=v�;–ں་'�]�E�\��f��B���8b�>&�v�K�k�AD������ ��s�J��9�z!��!���؊' ��9]�:���	7\� ù3��Ez�Y��3�1�0�U�Ԉ�Z��wr�p�t��Y=K"V=�͔p�\���0w�R�{��,�9�S�������"�:M��YwF��%V�P�l�˼�D$��äDo؇5� f7W�m�o��5��b���X��}��Ŭ��nC���������7�fy�d�]F�LK����@�	��g陈��z�M��Tt0�fK���4��M����\E,RU�o��������T�i�������/ڍ������p����r�.�x�Y&u�@$D\�$���ȡ_CK����c����۳�zY��C((�C\b 2�"q�:��2q�*�*����u�#�fs��n��8'���3^�%��6�Jd�{���wG��!�q��e�v#m�j���c�T΅s[�HÉ�#�{+j��"�����xt�O�����5�+�Ȋ��Q��������S<����._〈��\�Х+|h@M���Q��(ǫ|Ȃ%��ru	TuĞ<>U�˹�����9�z)�|�]I�`�\���y��Ol!��A��� |�6d�A�G{mxp�!��.�9�ʊS?Ӡ�h!��r�������Q��R��Ɍ�j"-��"\��$ȇ�������CV�O�7�,$��9M�a��<V)��Mn��/;�Nn���&�	@5�)o",}�|�V� ���Eu3\�2'~���	y<����GY���>�wI})�Jvw��Z��U5���!��.B�}�4�#��S�t��1/[��E:�g7u���J��nGl�������k ή݃g���"H���������  ��IDAT�����uy�2
1~v�9!��+�`�RsMpy��!� /L^_��Q�D��&b�`z�`����MB�bE��A��OC}b�Ex�9��pz�� ,]��r	��*�K�n'���#`����E�v(W�{��$p*Aq��>�g�83w��%k����
Y��K: ��sdO\���|�ި�k %@ڿ����D����(���>orVP{��i�KC.����r/���!K� R���u��j�\�*Z��AF��H k�	/*#>*�`��	�;"Š#rm~����h�S�(��"
����lOo�`恟SmDr���d����v�6�-�3[�Zx��É�4�#�^K0�# �D��Se��y"���._�j�zq"�!OL2���D��O��k��Ȟ�8�8Ϛ��]�0tP_x�܇��`?�[W�Ǚ�[�]�އ}��c���pb;��|p)�&yexfc��@��ڊ�0g7��|��&�]�Z�ޭ2 ��q~���[b��.�u�5�y!i��g6�����؏����T��ve���S�ƅ5T�O�Op8�F=�U'l>��D�?�9��^��L߈6B_<�y+l?k��i�ܼ��������zξ��m'�I�Fz��1�]é���WB@g�	A��ҭ}�O����u슰��۹B]`i�K��8!�����xz-͖]8!�Nz2��Sg��D��?��y�J�<nO����cK^^V�X�e�;f��t,pT]O8vdȻn�;Ա�hf	��5B�,F-C?�%��g鉗yI�XA�����?�w�'�@������\yu�����Ydb%|������4#_7q
���L�U���w�����0 PE2����`�|�$��o�����N"�����0�f���D��p��[84d"f�W���r�`d�	�:8c���OD����\��>�q��O�X���*�L�9��|J�{p���r��,GB�Y����_����Ə���LòE�p��f\�=�������<��V��V9������0de�Rg����u^_C� =��_�b�1\R��0�n+�#�~���Dʲe8��"� ��<�����6��WG!AU!�EjV�s�8*�<z��+�:훐��.%<s�M�a��8ln���Cqm�8�:u@]#�3]����G�h��j���-yIm�Zx�%5i�T9\1rƍ�;����@BJd��"S�B�<z�2�d�z"�{}	?=#Ĵ���⛩
y�Xx9�!����&Sy��f�\�op})���m��T�ғ)�W���uʐ�n^x�*n>A�������f"��U,UV�<��حNu�n$\�d�d��6zH!��&���)��f�U��_�oqy�J��){KEި�Xd��)�����RO�ԕ�G�]ج��ڶ�Q�60%�3���z�p��^؉�a�Qu� "�/Ñ�����/��Ww,���^n����;v��E[��6�8_�=�����ܹy׫�PQV.,g|��!�*� �cW`��B�]6W���:��� W�q���Ӂ�����k �����N��uT�����S3A�	��qu��%W0chla�M�����UZQ������(!�[�C��og�0%jk�y�1G�٪&HW�F��6��,�o�_�l��hb�t#�ң�
��#���|�.�L/BQ�AE����wo���1r�x/+�����H#]�m�	t���H!���l,�j&iX7��a��XwD9!V� B�%�:�Զ3���R̿ǃ�'���"��J�}�뵱����Dv������H<Q�����\ev�LЩ� ���tm��k/ ���'���"׵�X�M�:,$P�0�?������'b�VL��8���G������b���8�}/�܇�[�����r��O
�;���ۃs'6c��ؾ~�-[��6���s8t�*^�g ��1��V=��1�n V4B�:ޓ�K��=��v�ۜvS�������iR!�������u����!o���t�r+aśڵ7��4��Y�u�m}"����e�D�/N��@kgL�u�j��db!_lT7�]�X8M�*g��#�x�Y��A�����g`�K���6�����! /������ɛ�-A�����Z8����.H�tB�����YE`˧�c+���O�<���1��֢0'���Ĩ�p�.pZ����db�R��� %z��	w�
���5��{-| �\�J-~��u'<��MK,m�����W���g#�,>gGM�JR4H�`U�"c;,1��|S+�1��O������7R+z���X���!��ߔF��� L�Ԅ�_<��ͭ0�*s�����K-y�t0EQ�:M��<ŉ?�c
�x��i�)�Ƙ��?[�w�5�N�`�	����cW��ȥ��3
��#�}Gn_ɧ$����n��$�Nm®������;u
�,Y���@޷�6�EX�i%���u��=<�W�[�9��MCzl8}6�4�����9y�W)��eV|��l�	���(N_��W�i7��ވ�E�qܵCc����h��)�pl�\9u�ǫ��:��n�W���31�}�D��z&��ʚU?"�
g��U�.�3��ig$��"��.��
�Z`5BKr+z����p?�<�7Q'�$qk�~��:"���ug���ۻ�q����r.�����ki����wq�|��њ'�2ܩ�G=�����i�
QM�#�5��M_��k=���z�C�x��>	�V٧�4G���g(^t�ڽ�"g"u-��ﶪ�Ҳ�*)"T��4	b��y*f�8aK0'��d95�4�i� �����0U��)l�|[�~����Gb��@�q�]�®!_c��=0}`l�1��mB\�6����b���iȷ�ק�z�����4!2�Ճ%鞩�����H�}EC��y��M���C�'X++�rmAu�s�1s=��{"P�
amu�Nۨ��ǩVj����'��_js ���u�����L�L; ֱ/��2u�墭|�v�)�i���Wx�R䭤��� ��b���l��[!����1a�b���^�,E�&?��� B\ƙ�#Yb-b��}��.CQ���V�Fy�\�߿QZ��kU�<����͆����A�m�.���B�aOk;�HUB,�&ܶ"�h@����Q�	�6���$���F6"��u�Ef=h��� �Py�o��e"@����Bc��~�5dN݄`��(P�q��-������8���Q����U��s�u#���Yv���늻��i���{�I7+�_���8��
�Jp��9����	�C��p�K�9sv�%�[�3�����?��N����q�oX�#��`���@b�[��'�GC ��x�+Kc��7X&�V8�m4#`���B�Oɚ����Tu�y�@V%����v���@�|��[�pT#�0��r=+�v�o�iu�0����wY�ޖ&���ZL4C�����ͰU�DX�v�Q�6�y+W ����-�ŧT!}�
���󺶸D�t�&l�MiRe9z�U{�;#����E�DA,�2��t(R���b��F��v�ȟ~2s�%��3^���'���9h�vZ��TuB��!�\�2#Ԑ��H!�E(�W"ݓ����%凌�p���m��m�1��
��BɅ(���ޯ��p";U���Ȟ޷�B=�#țen�T�1�%�f��
c���!����|�����a�E��%�L��O}y��/>��-�4�_��hV��,^�����Ř���	m�a��&)� T��=����3xp"e�� >	��CT�_#a�B�����Yy�|,q� y�F��ģ03v,�,/��4����+X�t�_�����&�l:�"7%�O��ճ�����d<�'pl`��pNd��H�����iӞ�W��H��ͬ��p>b�M�~�0�7i��f
Bކ<����Vw��@���C��Hu�O��+���`��5��%�>G��M8���ߌDĨ��������oF0�D��5	�����Zٲ-�kqk}�Rg��[��V{"����%&!����y������WZ��)�/�����H<�Z�y��j�� ū�wzxl��B��XB���������F���@��5xz��P��R������>������uJ��s�ϧB�R֤͑��K�{�e��WB������	�������ZS�h�h��Զ*(գAP�����/^��5�[x	���@��G��U��~?��:a�_`�������!?�ǄY#1c�D�^3SM��1#��^��j�9J������[BMM�'/F����^弱%��gš���@
y�Օ�*,A���l��,��X��=�F>�O/���[N�@O��r��N��ᐆ����C�o�	,�#|�F�,�'ڎ��$~�q!;0T��9����@��0D)�@�^�*:�'�
�1A��)b	�	�x��U+/>���H I�tB���Hr����B;)'�}���w�������v�Q�h�l]敧�����7�A�d 
��Q$/A&�p��b�������|$�ƙ8u	���h"�K�ǎ���9BHD�DӤ������D��GYz�H�t;����Qs$ Q�ǠĨjT<�/!V�F�&�svA�H��D,�q��`m��X��ڮ�Y�%��9K����l��߯��#�p[�QU����رy;V.Z�u�W��38�o��q��ٶ���V���Wc�X�x>�mX�5��bۮ���H��y����z\]y����䭗�`�r=~��ʊ�����/<O)F��c�A�g���GlԶ�V	�Ao�Z�k�ߕt��tj@҉5o��� �������1�2[,�5�z-}���p�"�z��	G\�5���P�]��_ga�����p��x����p�l�"b�^2��1M��5�-��mfA.����yNyH�~�˵��;!ӱ���4~�r��^��ç�n߸�ԋ�px���ጚ	�S�g�+��@)u�r;�D ����$-�������%OX�\�̲#�	�B���S�D+,���|��$6Ǉ��n���ژF�a��%[��YD�l��~42Gб�t�ҙ��sȺ�{����������;����CR�?FX�
K�_FL3�Уf�/T7�5CL�실#>@�u\5S�kb��2~�����
�5G5�[�34#�����x����q�ˏH��� �4b��y��V\����'Q��ذ�ؽe%u�5�����X�hV����x_�&�]���Gx�8�B/!�紀<�SG$ ��{p�|�Sp�����S@^�K\����^C��^"�4�D������/�kk�X���<vUO��/��
[����&�]sT�� �~�p��%�@�sK� ���
�CV�n��"i��!�ROA�_3�O"AK]�]��7Q!�Sx�>���x2k2���,�x~�'��w��E�" �+���]",���(*�P ;.��mD��Y���D9c�2�O�&�Q��e�.T��9҅���I ��By�Z(mk�le[\�vǣ�|��Q,e���Z�?��_4Z[x�+��c��#Q�y��֤%"Z�G�Ah;�M�qךd*G>�¯E�I�rt�Jh:#應x��OuɅ!-پA��%�;��	M�*o<��iˡ�� w�����}��bȷ1u�7ؽs�v!%����c���� |����,н��-%h۲\]p��Q<z� ��{��ƭ���x�V2�����R�)���~�pN�Q��C|JE]X�ε��<o�:>�r�����k�c��NqptSG�1댓]@̮�PG�-����}U��F�����5
[�*�b���l\U�3]�g.Z� �to��!�hR�cl�TcG��wF�Go�:w@*�O����	r��"�s(�x�q�}j��Ԩ�����6�1�T_��B����.:2Uw-��%���#���4�j^(WpD���TM�J�7�ƢH}{�И�@�Xm>yl�8Ck�y ���ڎ���%2��F+=Y���������e�J��V�+�Y�Q�?N/F5�t�l�(;!]� ��.N'�0�D��	L̩��e����Ŗ�l���q�4�l����^�<y����]��m7cݲ�زf#��Y�˗bצU8{l|N����۱o�J�ڦ�+�u�Z�ܱW�/"��6u���	�%���c(VZt�-xO�F���V$6X)��QV��`��)N�Z�zv�5}�Xv'���(�`3M8�t.�XaD��e�?�O��������8�o�]��D���	�.[�����@k��6��d/�r��;ሳ������P<�IACr����7\4p�������>Y|�k�1��)�^����X"	��\�N��{�Rli���LT�tDv��������qK�����N�d^>�S#~�1*�48�P5@�v�����4r�}�dy����!�O�r����o�^#�=��H=+,PR��T����S����ɳ���+��0�@��m�?�\cQȣ��1��~�5ށ�s���wI#�J�!�=��?�Q�i'���A2�f�y�I��S���F���NǉoFar{5LRVŏ�����`]	���%kO�v@�VlCŦݨ���n_ ����C�ylQ(��'���I��q��v�ܶk�,ö��r�\�8�)��9�ާv��}��FVBң�wA��"'9��b��Rv��v�ܿ��+���w����%�U�C���S����s�G`��5*Hm�)���i���
�n�$b�	��V:$(ln�,IOd�)e�Q�e�o��f㝉��z���XQ1����{%��k,�z�C�w#q΂ed�TEB�4Q}'���<=�ۚ��r4�K�VL��L\GX�d��>k[�)��9���x��}$������q�@�!/��<�=b�|�K������RZh+hr�V�iKyj�����HRuCX�@h��a��m����%�K.+>1��$_å����y͍�D��R��ۋ}��6���!�Cv����l�r%���3D��-.��h�.��Q���z}8��'M�b�3��=3/�������o�����j�^ف��p��IGV�Y�Z<���vA��V��f�n�.pwt��)SE�.�%�s����*�Ï2�����]���V?�ki��*��V��%%m\V�K�zg�pZQgI��$�;�a* o�����{��(�m<���4��4�Vܾ%ڳ�av���&K�W��ބ<.g>��0���!~�zx���o;K$��"A����j� \��T�kv����H3KęX"��|�YD�~���W�� \ �i�� ��߼.��߆<~�{�&���=o�\�>�O_����$�]��oP��	�JN�P�D*�aJz��wB��;�1��k�(�Έ�pF�~Gx;��ϓ� 6SJÔ�� <���ˈ�K�E�����"aA��ώ�/;��/'#R�+2�z�`���]�k�l#;����"[���^ȵ�̞#�7c5��C�C�M�������'�ᨢ��@��Wn��%�pp�~�Y�W."} 1�����D����m�f���/�V"���mԛ�7���y�����%�k�Zw�:����������5<2�[���%&89g	�e�!}�&l�xH��_�Ab�v��D�[+a��1�/^F� ��2�	�c��ǭOJ|�y�.�03�v�����0���G=;ဣ+vjZ�l�oq7<uq���v�i��xؗLl�k� �j�H��E�@G��!��
�f֯,yQvq� فږ��~�N�*��(�싄?&E�
y\�ڤ��z�>����/���4�`�2ȫt�;����M�ɓ^=[��u y�X�;��A�Sp��x,m�"b�Yܠ��Y�
+m�0GA�$��m�:f�-;F^e��e�S�7R��K!������]�=�D�٩�=����k�%&�H0[�@����R����zJ��q�b0v���0AM?��b,l���t�U+��fo�w��.��V�o����  ��ޑ�W��DJ��P��n�"�/��p~/Z�5�b���8rt+Ο�Y��]4{��uKf ��$��pN,�ںaW.��ݛx��O�Ko��Iv��O$j��ۼ���v�r����87�O���������9*����G�;Ino��6�kn#P~�*����y=����-�B9� 'A�^��Zۀ�E�q��x\p�+z��U�@Je�}Ɛ���&J���L���E���v���녊}G	>��*eJFj�#�{K�<eʀ�}��}�z
O��7©j^����	�@EC�RI��Q4T2[( ��"�Pc[��u*�#r��z�0X4�r{a�c��һ�	�4	������?i�z�+t"�CV;���՚�JN1D� O�c�Ҁ,������im����H���G�I��#��IVOoB�G�?�#����z$E�������s|�o ~�n F��-f���;�!���c����N,��~��7��^�����_}�%�O�� � �=~$t��ʇ�����P�:�Ez�d[^U���j�����a:�x���A-�p��.���>4a8���3�j�iR7��Gݙ��D�>���,\�,CIEy5Tn\�)���9����w�ID���%-O��:C!�QV��c~�6���D���"Ԩ��K�i�x}$kKaFI��	��̐��L�o���<:)/�=�P�P�p>x|���� =.ߥ���*[jS������B_|��1�>#b�� �χ ��_�W�Im�E��E(8>$a�1�ݐd�I����H3�����0��Gֹ ��{$`D�^�G��D���y�K�����ԇj+��|�Dw��������q��Eu�k����N(��\���/�[��3�����§�j������yy�7	�(�����g�o��}V����������݂��v��9o��������&���u�����y�+�{�^,p�
�-;c��V�x.\�ح2�r��I���7�މ3Q�V����鳮8��sd���N^XAz�����*LQ1©94�R?�q��'۟^��L��'�;7L���-���swl�q�6b�m���K�r��U�[خb��ݾAmB���"d�8��S��8O�t���f��d��.S�d��!�b�; ���vNH�s��d7�'�ڹ+��"�����5"n��L� O֐e��M���[(&e8vN�J!O� �
5��Mg�0��H#Z0�	!�cyf����e�/,��̱�8��ϱ�v���pe�n�L�G���Xjj������D��!��Ђ �k�0�
�[U-�9O��q��F.k���@˕���뢗Hˀ��f����u0^�D
wzx{�$;V�ӿ�k1��쏱����*Fj�Ph�(�3w���r�i���D���h�Y���W�"�.�?B�T	QE�mf�d���8q� N�ލ�G6a͚yX�~N�܎���a��y�6q���+l_���sǐ�s��#!"�~�髓��r��A�-,�b�����5��N��HY�1�`��B�t��a�Z* �`!��%��r�( �@���%
u:���<\�����p���G�>���7!�9~�:�{���7:a�z�,�2�r-[��Z�|��(����!�����Ώ�%�# 4�@���@�uR֌DRpkT��2��c��������e5��Ża�	im%Hj���ڈi�.��Ǵ�F���L���QH��>�8̔���:����&`�a����~�(�\��OO�;�;���!��	�B�v���/�!A��[Ӡߎ�����*"��&*h"K�PD��X�ѭ�'g�%{$�� ���(�tDJ�R���_Co�`�`�[�+��0j�̚:���3�a�ز~1�mY�K���~# 쇾=<ѵ���:b�#p��%ܬ�+�R4<}Dx���� �����|�~�?�yy|��V���ů�#д���h�3�>mI��==x���I�հ�&=��3�;.�vv9�f5��QVV��x���կ ��A���V��C��5��I�EJl��߻SyiG.!��i�b�!�}��_u�I��H>1����L; ٸ��2,"�럨Ys��>�5Y�u����p9q�瘵o�^��� ��#��k�{& ��96�j��� ���T��(��)bDk�"Ħ"\h�l�5�-�D��@D;|��nc���R*﫢�rv4x��ې'@�ꏅ����&˿�i.O�8���׋�4��í�P��b�t�n��o.I>���Y@����?	g��3�X���/L�!�����ն>�8�,�li���O�q|�z�9�>g�w��ٶ[ׯ�{����+�p
ϞAfZ�<~
vÇ��S�ܮ!�3�O ����i@���X���/�!��&�Xef��b���m�9��X���i��X?�7<L�E�	lp��|� �����X�H�	�&Ѥ��ĩxVS#���~z��3�wk����_�(skl��k$��ld�m��½�~�Խ�)�4-p�����+E��ᔆN�⬹-������@��A�Ma���؊ǐm�nTl�B�����Ξ(w�b��G�y<M�?��t�h\��Hx�{x�&
}�7�\t��o��چ��A�a��x��u���:��pWGd��kȫ7s�S���."���<w��s�;��Z#̰v�Dk��E�p'-�����s'�n���jژ�k$��M���s,�u�b"��&����ר���Kj��:A3Bq��Yx�El|���
����!��a�3��J���]�`��&Sc�hb���F"~�R��9Z��弄'�fd	�Da�gO���/Jr�����:��q���QB)"{�X��\�5N_�|6��M*w)k��w8V༔��!�SR��n�عǏ�š���*�߹�����0m� ,��fL��E�`B�}���B��b�g��n!_�������卷<sx|6�z���"�tʘ�pH��T�ܤR�4'�k���r('�+k���fz(W�$R���7��4���.?�dJ\���K�?=���i,)�	��'ऺ#��-�H2���9eı�7��G�)oi��6��om����4�������T�V��
������=����#'�φ�Ԟ�?A��0��6��o놤�f�nB@�TO,)g6�D5CNīZ#Ƶ2�LC�ѳ�8���u�fM�^�x�~��Q|�����s9ޟ��0�^�lj��V�(mc��:��z��I�pby)�"C�����|��G��{������,g�����(��Ӈ�0�E����z|�/�Ĉ�c�1~�0��K���� tq�[/���V�؂�Uw�/�o��W�]0�	�3\�<�������
�e���.F��@\�v����R'(y�Y�Rs��;"V�A����.�e�G����×P�S ��UVU���5����5T�Ox)�֝����K�����g�������2�@M���n_㜤;��!A��j��t��q�ZD���H�������f?)��q��	��,�������ݻ��wo7^�M��7_�6K��x�`5(i��#�����-���`����~�<p1FoD�C�:
�)_O Y�n�����J�{]��R�d`+�?�<���T�<�����|��\�`�W��K�?g�\Ir�>�+rF��h�yTVoʿM2P�)�N9��{����!))	aaa	
Db|4
rp�f����}P���xC^��� y�yj�#p�1,t����kLl�BbE�g���n����X���*��M��vh
�Gfb�����&[�lD������#{��f�V��	���|�����˘���2~����O�w�Ԛ���ΘKp�˽'�X����w��-�c��1V���嫉j�P|��^�pI���s��餩5��]�uye��5�C���+^�P(}�}����8���ppA��'��:�{w�����,��V���D�^ߠ���;\ �-?��<o\�s��� ���&�4����� ��h� `����{*q��)�m戇�.���ǖ��f��)����b�����9t,*"q�JB�qe�\�����M���
뽺`��ƹy���-xA3����˭�ҙ!n��/!to�����cL���pB`��r|i"���	�?>a;���"���J*�hl�ݓ��A\J���r;SQ��*��Uk�.���x�>�=���Cqc�:{Q9uF�<SY!B�0 �/�;8wlV�+..�����˱m�Jl]�X�߽u16���E�Gb��:�{̘�'�:���$ܾsSXy�2Ȁ'*�WM�]���ﲭ��Sz��⛌��"x�"����h[!^]��8�i��1��5�L:���Hԭ$(�-��Ɋ�u[�������K��Ϳ��8��j�#c�b�x��hOo7�������"O�9ZY��D`~�?P���t@��fDj��
��M��f~��� ���8�jQ<��\F"��+D�v�n�C�2U���#����;��w�� �Q-�Y�g��^����ƞ��aL6*g�BZǑH��,uW�j; ��Y]�j�]'���P��<<>�OT���p�#~�o[&o��[c���6�"��P?�ć���1s�*|�(�,\�+������X��ؾcX�t+6�9��{/ �j*�B�\�R�A�A�C�'K��%����C[�J�U�f^
υ"v�v�|7����\��?�^����-�j������A��5FqMJ��2m�8�  ��L<~�8��-||���vٺ��x�ݪ��땸YZ���8dn9��_g#n�x$��خ#�y8|�����c�=t9�-8���UP�S15����ˏ'�bY��}�Sd������t��߸���)��x%3�"�~�]�A.�{�&=~��ǡY��<H�D
t,���~��$���M���r�h��eB�&]~��PJ�i5@�]���{�i�@��]FwB��=���$�^���-|��"d��E\�[w}ފ�!M__Z_�Am�俁<.���\��c)f���zk/�7����a��,�5�L%%��6��K$l:�{��8?k֚{�ë����zG�5��fsvt��Bv��c\���=R9���c�
��-=^�?h�p�}.��\��N�BD�8K��q��|zvF�Y�X?�C���8d��mq���n^"�Y�{g\����.Y:ક#�o�%Iآ�n���E���+�K��E�����J�n�p��>�(4Z���۷�	�:_70j�$����!�eBx��B��x���v��]�l�~<�<�=�5H�=5�Z�^�4v���	w�?�q;����DU,��чϠ>� �S�
�-G�X��&t��n��k�J���� �"K׵�sϽgfz�qw7����!	!Hp��ww�hh����݂�;4<���fC�@��?+���U��>K���t7�O�J�!c�^?ס����69�dt�L���g���Ekctu��6�:6�Z���>��u%�ږV6��wp���g���X9~	ww\dk����A�\y�omI�or
�{s.���U�`HEN����h.ظ�0��lr�fW)�4RG�&sD52���?`��mL7�S�0~�p��N����ݭ]�6�Cz}��o.�7Ajw;�u��&�� <�3A����~�I}��ځ��aĚK{�K7L)_�ɾY�Z�����*�F��-nE8�ȉ���*�����0��=�bS�K.��������h�1 ��n�T��l)Қ����Q��A��\Fjgq��ޜC���XkQRSFg`�#�eP�s&���лg}�dv������^���\�n����^G�%6ck�Fl�W��V�6�����"(�Q[cu|��SVk�y�Wu�Yb�;灄�1CY�9}�#C汦B+��j��ҍ�^�)�ʥ��l
����ͮf]y�j;�r)�n��E�[�<���?i��dt�ez;-/]���u�9p��N����Ü�pZ��Ժv`���~dꆖgkx�Q{�:���тU�I�'�Sкv��KWL���g.�q��T��K:�cL���~(��R�_�%���ď�9��$�pI�L'q(�]�r����U�~V��,u�Y�s����ܸu��}:~P�]�p�����,Xƅe�9��㛜;&Lg�����j�TN�H�To�0�t�9��.S�a�3ǽ����*���w�٭�F[���pj1��)h��䣚^t���F=���S����6�V�>-~B��.ֱ��4��5�Sw�)����k�L�x��V}.��y�{�=�9L!"n��L d:���<ʰk�vzWjE�{q�(�_����F7���^t�U��a,v�/����]�Q�o�_���9����`?�%M����Y�iZ_�Ҽ�\�.Wv2����s�����?�����5�az!yOյsgi[�6���
/� 'K�d���dlN�Z�02��ʔ����?���f*?Xx1�k{f�B�A�ϛ������R�`�g+d��h��U�S�Sm6���6�y��CXg�oG�"����(%���~�L�1k�Q�A3��]�_4��)����E�lވ�B�K���8��,�o

��־{?���y*m�S�S)���<�}�͋Ȳ�
�[.K��t$U��֑{�sz�"zG�cN;X9]�z�'t�w���/�E�64�d�)=����5�P��h�V�ǡd�<�1B�V�J��du�]<O߆��*��7�Ty�.^t�s���%�{m%��8�0�n*����⊽̈I�����z.�XY�=�+������o��mCF�`.Z�q�ʝg�\s)���赿+�t��J?��Y������~d1�<���1|`͛a�����LBS�ln�3ZI>����sF��G/���pq�Z%p�p�N�u�ᔁ�I�����H�ǹvC��u/�,�5�J&7����O�wԄ�]C
�䂬��UZ��qg��F���,��x8z#ۏ������. �3�8%C!��n2�l��a4�g*�s>g2�%�Ԋ{�_�R[B��)�ٵ�pBܰ��;��qe��T�iK�TZ4��EO�I�c.h�2��f��\�V�4}>���ژsM���?�;&~t�K!�C`s�EX*߆�pR�5��B� ���V ���9��1�f�S��V8�xC��]y��i��8n|�_g~�1�¸G���웆}����wWǿ�hk��7]�z� ��D�.]���+�Ν��K�G�s7x{�2��\���\�{�sw�]3ܬ�wIA��E�\��*���w��)�4g�����s��-�]
��3.q�B��W�����%|�L��gp��e, cZ&衶��_i�h�e]�j�����ǿk����3#�賌p�x���3�?%�hHkj~�K$�:���j�{�5����S��,#����l��L��wc�t�H�Yd���!�s�}���g6f���!O���ӌk:���	�q�g,�ߥ�&�~������lJ�y*ed��.��ن��sk�v������2t��d����>.>�bȝ�\Z��Q%X6�CFK�ʭ<[���q�k�}�s�7C��-�OZ��6���/3u��ehT1~�,�P������S�S�1EX`q/�Uoa��:��mf^X�s�1�ƍ�vnL�7mgٻ���+����bo�+)�u�6�ݶ�x�<�������Љa�8.�_ר)Ϥ��Y��&{�"��ȥPM�G�%cڴ��=�p<�*�v��1�{U����#�m|��St�<�2��kg<����P�]S�3?σ����&'����Ɲ���sb�F��;����hg�A��6t�q���+]�]����nt��GD!Z�+Le���4�׷�H�2-��0���FD�5}�ۦ��z^�MI��$C��Fm��4�Pڸ��Mj����NGgc�E� RB�j�x^���S��D�?[�lkC]g[z��m�8Ayc���|����Uk7C���qѽǪ��6)�� ��9e.�͡��P�>z�-��_͸¥�������Bs�6�����ޢ�����t��.5m����Z�ӱ2B�-f�e�P�Hy*@�Lt����ft�ŻBX��Ȱ�u��w�IXkx� @@���[���.��2\�F�m��r���ch�/�V��:�X���a ���wh���̈XZ���Ì�s�����F^�3>TFˁk���t_'��j�F[�ԯ�JN����L�}0��$2��x%�J�M���F�a<_�_�j?��K�������D�g�Ǐ$�ɿO��)���"H[�5��*�:�Դ��Se��7F��BZ���O���n���[L�G/��`L�0&J����\X:'v��EN\<õ�W%�	�~��G��?�ѫ�Ʒgu��])xo�p�v��^5K���n�� �)�� ���A�=ꦫ�L�Y�ĝg�]�.�|I�P���5�<߽|���U��.>���~����.mj8i5\�^MkF��.P��%�3+s�5��5���3F]�OR80�4��,���"M+�޹�>���m�s�iX~$nҺ���7͟�s�7���:[�'\̂Sh�]��.��v��U@��W =}����i���,�ݑ�t�ڊ�N>��=o�dF�f�u𦯭7�=C��艎���@o�@��at�
�-_�=3�/e4x���R��҈?���$ �����%o%��'���#�#��+� �	g���(�#
36(��n>��`�g^�3#�8��KE�.w[�b�G	~���4g�9�������[��"�%�>��c�W ������o�<cwh{
F��`���P!��������k
��B�i@�%����]ǎ�Z�$��H&�h�M�w���a%{�v�L��lp�an.+v���8��Ā���^�!Od���_�0}��c��:����?�3��̰u6>��B/54���Gp��%�N�π�����\B�r�D ���.��<]���o=����|��L�ӟ��J!#�+i����H�[=~�)fj �;r��m�R�7���t�����O���]���NKK�ɳ�Vm̍��y��(j��/�4�*uh���(+kc̧B��r9�:���u溕7�|��3�n�8\��=(����n>�(�%3K.I�5`��sAx-���O�j4��O��gd4���{���>mL�Q_����ӗF���R�6��|�j/$W=x���j1�P{e<����f�
z��7��w~f��w������* <5�Y.�O�V�@�a\�5(�*�}yZF�������0��_I��H�-�
���#L��f�"���~��vj�eH2#���$R�5�7K����]*c<���i=�w�%2���x�T�>u����'~ޘG�{1�h]y�Lq��G"}��S�}B!'�=�B�Rwn���d�ךAO!J馀�V��]4������z����p��Yn?��h�P:���´��;�-�:1L'0ܺs��7�t"�TPU��g��<�} <�;�G'�\�P�����	��2�H�_������/ݺ�nݖ:�	��Obǯ�S?�XY�z�&�0��e�LqP�x��J��3��f�6��緆�����Hw��9���ݱY�޹�L���������٦a�n7�*?����!ϔ޹���ܽ]����g|ɪ��]<|�5p;ٸ�E{ϲ�1�Ɠ��mh�Â��!��W88���]G����C�u�f�K(=�}�f����R�+X�a��m�l���xi�_s��2#�|Wj9��?=g�����O��w ��d���e�����C�1�-����o����p�o��H�f�̑�)�������i���q�6��)�--��x�!��[��k��r�2>m��#o��@�hNǗcO�Bl)ŉ⥸$��Mec��p�4N����M��l��ktAJ� �xhf�;�v�[�dEP$Krڱ�Ҟ���Ey�m̖E�l�tBE(?�����Y� �X��=q�S�q�~��~p4[���^�=E;���1���<-W��gY�.tPl�Ӗ���wp����#Z:��R[��3*.�&�5"�$��W�H�Z��/��n*�I��R��GO9u�$�.�N�R�s���b��t�3�e��;��Ó4W7ںy
��+�k���A��Lf�{(������us[��Ɔ��~\��瑇��xd���o��ǝV����i�vב@:.��c9����,�~2w��զ}�7]�@?Y���,�32��䙤�j���v��Ec�  ���[�J[/�`6����Ҽȫ�!iF*��j��k����)�����L����	�����w���n��w�(�����`��ib�HA�P&P�V��=5�}'y�9�5M<�qK
�|рf� �����k}�n&�S���}�ɛ���'��T龾���v�=Q�i��t�{f��:s���1�*���ج�5�o����x`j�Ww���}�*R�zǨ�e���«��=~`H[�tF����j���s�����.�K
a&�S�N��8֘1��C�y�^j�	��~��M�i����o?}���õgF�ssW�_�ݧ����+�2��m�S�˸��w� <]<Y�ז��b���)�=����B��O��K����Ũש$��5�ȵwƨ�+5�4��|��4�U�ܘ��C�������1?߬�3��9!���Y�33+s<4$�|,��|̬��|�6�m�d�����Z�8t������5�hy��h@�6�tu񠳀P�<δ�iO7;��;P�/_�*2���qo�FT�a|�Gnz�z˭���c�c}�|�!�8�@)z(N��Y;�He�<��S���H�_�ʫ�.�|�TRJ�!M�nl�r������=���İ(6��̶�Lt�kh(w�/��8�w�݋����l�n�;����4'/f	��R*��B��y�<���r����+�
z|X�����cT$[󅱣X�&'s7�"���vC�_��ϵ�i���@ǌh���u������{79�b>��7�wYm��jGw����&�xG�����:
�9���=㛵��?������g=~���O�����dP�s9�4���&�'�}����.L]��b�4�ocgO{G{�9;���J�xNk� �y��3� �K�ӳHy�F�n���o�ƶ+8�cN��̩Ӝ=v�sG�sP"���Х^�:yR^H;58?�h�"vz�N����Hw�����1�a�n?����XZ�*����_Y��ҙ��,aa�Y��Gn��s�֎G��\��ĥ��n��6�����@�_[�q��	�<���:�Q��I�P7K���Fc�YE�O���{��`&`g��L��2`J�1`�p�ܫ�$5u��ȐDf���������O��yZ8��w�5�{7�@�_��"dk�	f�3ܜYfx��b�m����F2߷Z��J8�Wu�qNP�y
R;���j��Lc�ѫ�*3�ia��;Z]��!O J�XlR�S�Sw��La'7k�^�zWP��Ϛ,�'�2�IdD]1�U�<K@3����<��H@�ׯ�|��ݢ*1�+uB�yf�υ�9��<�/S����]���e�]��-ɏo\�s�ِ�ȽZH�V%����0��T�Rwi����4�a�y����)�]1@��e������{��˺t�ū\�t�h�������Ffe1��ƫ��CyE�o抔y�紅��A�Ԫl��ߐ>I��F��Y?g�w������i��l�G�P������TWf��f>o�?��~�ݲz;]�Z��'��~E��LW� cHT7w?cbeOg:
�氧����himE-+v����ut'��BO{_�@'z9�k����bg&��Ȉ���Z6��:ug͜�\;y����H�?Vo�0�����e�o�F&��M����G1^���{0m]����> B�қ�>�Lץ`�m���cj�b'��U���+/�E0�?��Aa���~@�BY��b��e:�A�j�����^ۃ#���N�l��a�����e{t4�+W�jѲ��	e�v���>y�L�v�jk�9Rj����mcLޚfX)]k��{y�4��yƘ;�WV���(��趵�敵���-���3'c9�����#{E� ���b�ӝ���%d�2�,�箃����g$��H��EGkZ�X���E�˓V��mu��o���P�<*ա{�4�nM��	���L���hS�*���,Ijy祶{�Cc�]����l���B�W �����B//�䥉G�%T?���\����I��?�(��!�p��<�<���|ܲt��D�G�G�-<��͞Kq���=�p-ľ�-��ɴ4����f�ILҘ�>�yW�f͌�6�5*f=�盿z����r��\f�c͇�dz�G������g�d	g�G�@S>�qA�Y
*���s޹+�sMn����gL����BՀ;���L�{w��Nǵ}�>%3�ik�/���+��qK@�S��' h>�V9͏�|lw���zl2
��.�>0�Ϝ׫Ҍ��9s럹PerǇ.]���27h��J�W�Tc���Q/�(+�O��?ټs�{���{w�|�k& 6U�uL�[����f 7-�@��������w}=Ì1y|���~t��1�����K�mCz;ZY:3�\2g�m�s��3h2�B�+��{��ɑn��twp�󠽍+��=��hkZvdp�*t�ObL�4֍���▓kvpj�N��������i�pG�Fdh�X�5p����}�2:��J$1#����c�bN�:p�&��b����*�xw��v�����~` 3�#�΂�h��e����]��8[��J��n!l�c�W0�<M06{���ߟ>~��)g"�s%����Asa���}�c�4�j�׌��H5C�ں.�|a�2V7��j���qb�����ȋ6 ��+� p�3Z������ڋ�6> p�L`졀�{/��xݶ���O��<�-ȥ��nJ��NT�r��C S���<�q�%-Z���[�N�˝f���;;:���ч��.^Y���JҿH!z(J��42�矗Ze�%�5�8]�
�;�0�����I��@��'m����Iι�/k3r�����y�r����F0F�-��M�\��o��tb� ���<���ƃ{v�ܰq����<\�.���=����g1(���ؒ��g���$s�c�ˬ/��1��3 N���,�h>aja4]�{5f�f6z�y=���b�_�B��̽ ?g����?e_f����?6�ә};���F�K�uc���O�|^�v?�L�n�v�~�����.�_�/�w`4��`2ŝ4�i��%���P�.�Q��oκ�I���c�(��v�����'��@�UN;R���66��I���C׸�� #+Ԣ��~)Ò�����p������r/G/�Y8��V�u����uW!���bHR-:M�m�D��J��t�_�N��� Q�����	ں82o���o־����p���3�|�R �g�OgUTE��2C�lA��\���`�$?���2N`mb` s����"g/V��k=�Z�i�K��_6�s 6�=����NDr&� W�sv�jKޛ�����<MК�hf��Ԝ@�kF!�҆�5 //�,\Xk�%�γ��U��N����7�i_���9�W�yy��S{?^��q
4�+Ⱦ�+�<y�G�"�Px惘J�,�H	\�����i,ϙ۱/o���,�ۜ~~����4��'/�孕�7����a%��t���g(�F30�8C��1�p<���}@�|����!��{�99�D�1�Ϗ�~�{��V"�N��b�B��Zӈ��qg�F��g���A�?�/�Y{R�և�	�D��nT1�K�ܱ�垃�mݸ���U+���ܷ�����E�b�m �wF O�:�2��� x*#a���S�
_��c�����11A����u��U����̭K
=
%��)��a%����I�PӸ�_z�R�.3���d�=>��_����+��;�]�����������j�/���;2TFp���?��h�زt�{���!�x�]��, ���W�!tq	����ml�I�t =�-����榛oqN�_*e�v�0��i��"0gO/g�:���ځ~R��r����#���t�dP�BLЛZ���WfT�J�+R��%k2!*�Q���� q�@�P��eH`>���3�3�1V�L�����2�t���P^p�N'���&K�:x0�Օi..�f��330�I�~L�dQH���X��f��	������$l��Ƀ��"'7v���×�~���"�3�>Q�i،��NK |�4���5QiFhH~Ԗ<�wq�2�4�gL�]�ە5��p��+�E��x-��� ���1��W8o�"y*T�D7������(�S�z��x��4�<��S��2,�����R�!�&M����2�Iuk1<�,ck$3�r}ʔ�G�B�)̐¥�U��ޡ4qv���m�B�R��^tr�K�ӄ
[G�yz��ˇ&�4�������gG;/W:yz�V�L��Q�$���Z�Ǔ�;�X,�_�������h"���-�	�x_�k��\�c�mK�ڻsC"�G.[{p6�	�}��Y�B쨗f|��_yj��f��{�S�q&}1���O��yFc֖���w�f�SQ(Q8�5f�ɼ�[�-z��~�5�,u�ګ]�����]L&�ɘ���}����c=�y��v=+T�/�rϧ��a�Ь�1�c�Ae�)��6��
���y��}y]\���k�ĵ��~y��kk�a|����m�bEל�|�ΰ���7�_���)�T&��ә���+�.�8���MO7/��{��������#�>����%�V����W�1~1��k�k|w�k(#�k���][�d�w?�08���Ф_��^=6�t��,��fV6o�81Y�l��S윘%n�(n��Ջ�=���,7�9{�A�\+n^)n]���r{�k[����\L��~����o�|#���N�(�5k��<m��L�� $�5 4s�$��%�� �`�4��zOh��G���>� {d�ī<����ڄ��%��_�bJ��L�4ffz+z�hN����J�a��4�ґN���k�X��jĢ�m��c_:��C����0�)�f�ad�J��wݓ�V�����>��C�\���!Сtu�����K ����1�C'sts�����NNT���C�2l�~
�x����_���8� ���W�]ƍ-�Q �{:�@y�|mŵ��ܴ�嶕+7��o�xq�ҝ�܎dds��_܍ٵ��5��c�r�3uϚZr͙����j�W�2_���/���hf
F���4_��F����wf��3f�*�h�U�V���X:|��������*3�)0���<W��<>�s��n���[��1FӶ�?�}3��ev����3���H"���������KF�ݻy'�*��2�4����D{'c�;j��1�vR&����8��I{7�Z���+KR�����n�� ��]�.?e���W���Lk��q�5���u�dh@0�c
3 0�X�E�ESH�띗�^a��Kga�.�����}}�k�c|Ic�G0�=����9��_3�WOtQ����ms|�3�v����x[gF9:2�C�N q��7c����3�˟Yށ���c����t�*?��3�с��r�0&�n�����.�@vnw����O8��"��ʆ����̵;C�
t��r���w�C�JyȚ\N��vg�Pn��Z��x#��->s�1w��p�k��{���S�`^���qp����M�Ͷ͘ۺ5zv�w�4�ډZ=��Щ-��4�X�T|�T'�>�jp��P�L�GPq��r��46�L�~�t뗟�[�p��@��h��>���{:CjT�w����}`�$`S�%ٺ�y�*�A@O?Y��ڞ����kь��f��sܚ���ej2&�m%�W�&;U�\i���`�����R�8.�_\���'�۸q�ҋ�9=�m�i�ɻ�ۙ�ٝ��g7�9Ű=�9�;�/�gJܙ��`�RR��W�����������������,-s�!�z�����9�3�I�9����OAUf�����y�z��=��f��5�ݦ�r�ծOI[���~m~�����ܭ��Чn��;������Af�)����O����G���C^g�@ڻ���u���7`�����Ӏ����5�nC�?[�Y��k�с��qo�1q'�����u�I�������4.o��?��C�'e�.��G ��^z������X�������Eo/?x�_ܤ3f���:[w���]Nk�sY1�h	�Μi|���\�<���+3�F�tb��#��jg�h''&8y
��2C�ruXA��@go�ͱwe���y��x�9,��!a�s�c�s ��%��)��.�����A�P.���C�cyݺ���$>yﶆ�|���wy�B^]V�	�9�9��-��Z�y��kg��y�L��ʋW޼��g�q�BJ�4�4�ĳ�B2���gl�z�oOj��4�ؑ��MiFx�f�k�{��$�ĭj�իcW��%�ӴO0G��e��r8��:�ܸ�h�N�2b�'��gl;؅�%ӤM�tiȤ۰h^g��Iz�bt�-M���Y��ڂ6�Hd���A�ݿW���'��o��`Hv{*�����rv�����}�R>�kbɰ�㢅+7�\�c��#�݇~���Ń��<���~n7��t��ݹ�X��Z�a	������2�QzT/����ע���&$S7�������{c���ʾ�+��Eh�_P鄌����h4^�Xc�O�Sf�!-3�)Иǫe��s���~Mk���O=#��n��_k��˨�ӻV�Խ����翘3��g����GC�Ɛ��1�A'Z���G�#:�
ܹ
�	L���#�N O +]XB�·vTy��<����-;�E��.4����Zr�q��{N1�� ڄ���?=�9�2R�b+�f�G��P��}.�O�����0gCwƺ3�҃�_���/���dL�*�]�D�H��˜oݏ��ř�ۓ�Όw�`��#��a��-�981B n��#s<���3_�3-��<�ma�\K��z1�щE��l
g�v�
�n��c�e r���-��>�.�q�0��	�y��fm�M��+ O�&X#�J���k��56��9��ڑ�n��z7��)T /�;��yh�f,���N��%�{.܎(���d4���V]�ֵ'}���j��l��&M��]��u�U�*�&T!gŚ�T�񕰌��&>	��:���l#'��h����J��Tonɦ�]�w�#�����١��6���2yi:��է��$&�h���1`|{�4N�G��o^�v��"̟�~��Mb^��Y��{'Nr{�nv���w���É�?�I���st�fn{��aJ`8���� ���䖵�츑ә�6<�
���a�w�'~�0�����{IN�� �����T��<}����q��S�e�&���ocn�U�f�3�ޓ��L�}'3�3�ߣ�w�1�
H�.Xs�cV�2KaK!M[�U�ם�|_fe�C���
G�3�ӌ��e��U�~��u
Y�,����{|I���F��BS��3 ���3�l�U �$i�s0 ������f�K��7����K�w5�<�4�ͭ�h�#'�-,�.�&��}�A�OI���$��
.=e}��J�����Hv����c0��C�!��C�zx��[��GwI��1�Ƀ>���wp��q���=�[�2GFN�xO^q�f6Wi�<�|�ۍ��ìl���h[[c���67V�>L p�o(3���<s��S�Ù���H��E1?� ˊ�`]��,�)�<�HVaST<;WfGLEH�Lt9N���v`4�}BXY���hfg�uV�qK��]'A���H?���e�-[�چ�X��Z�X8r�ћ�B�ϝ���6���xm�+_^����3�{a�9����Mժ�Z��R��l�FX�ƸV��}���%�¹J=�+��)��ձM��uŪ��!A����Wm�C|�bC=�./[�p{~��f�Z�w�F�^��=y ]�v�kz�~����l�U��g[2vV2V&�zʷL�~��4i^��&u�з?歁=Wa�I���ͺ����B�?��~E�lyH�nE�?砝S �
�q��x���1��jN{��r6t]_�io���,}���[�\����7\�)��F=�$��m-�ټ��O�#��Woiw����y�d\�Y_̿�1��]��U�}��3+s+���2C��+S8S03CWV)P���g�fU���h+�ڙ���vf=�S�Pͯ"��{�0�)����_���|1f���ڔߛ���B����xL�~u���kLn=���r4q�Kc[wcb����/]�:����V�^�֖<;W�R�]��O��w$�Α�.���u�av[��k�,"�T�����{��]G�<�Gfv�F��d:(G�(���#�vΦ���s[��҆V�jgcy^]��`IƧ����<�{L�hy����fV�����Ðn�ue��+��z�1Nܦ�7�Ύ	��̰�e�g>z{��}�*��?��'�a�L���y9<k>��������>���Ʊ����_έU��f;��_Ʋ�u�^�+᥹�_��~Ѭ��.�&^dc��
��[�i���}x�
g�,`M��,��2�W�g��+oC��[�XE��JE��W���JRM5nɪ�=�Ԯ-eS[�R��k�&{�jXT�����E�*���ĽrC\d�r�P� =��IX�KĲT����Hil�&�X�(ѕ����<�_��dkCzO�B����ƿ�?᱁�/gO��o(&�~[��iM����@A�.[�*�	�[��)��ֺ�O`��ul���u:3�+�������������ܔ�:U���O�XݶܬP�~8�r���r�r=������e�e�_��.J��l��=�(��$q�A7�����@�FS�ו�M2��C��`�Q���w|1��ƜYN/_��H���y
?�aL�)+���B����e�'�73������Pg�'����:�D����e�����kf��/�����e6��ޜ��Q����O<������R[���=�U��E��	�t���ݵ�!����D�Mqp���+ivN���#-��������M;���J�͹[y{�o�H:_��K�7sd�<�tĜ�m�.���)�/��"%�Q�Z���C���̙%�y��?��̽�{9�{
��[1ʩC�3�*�1����:���0;gFȾ�{o�yy3�?�I9#ﲬE+�>½�'�������������cn��ı���5e)������cؽlO�]���Ԣ�W�j����pP�bȗL-yY�X�����yzt�*g�ge��,�`��7Ks9��ƍ�M_��
v�<��TBM��Le\�n4h�FL�5n�k���U��eBU��U5Z����>��r�$`'���o9�&��t�+�¥r�j�&�~m��W!�V"k��X��݋r�ZO�ҏkZ�io,?̍��_Ztt�}wwf�/ĝ�u�t#����x�+H��5�c_���x֬Fh��ծA���7I�V�bT���ʟ�������������b6�F��j�м7���f���z{.K�����\�&��4I�u���6����m���&��Ag8�ݵ��_dL����d��2v����㨤�b���fԙ���$��Yf�3��`��t����>L��^��k�v����z����'f���}��o13�e���WM2����
�_@��5�s��9��GB�گ_{t�>s:#5�-�
��=/���i��E'?RU{�4{Ә<�4WR��h�l���h-l�\������G��75��@�l����f�88tw���w��gq��ȝ���r;��o�@�����s?�7��Ɇ�<_��S�q��X���w��+������5?s|3�.���������.^���}����柏�������1�۴�7��2'�?�*��d�vn����U����ƭ`N���>	vfP�1i1+����+r/Y/ܱ4_���FޒPޤ�w�y����'p��5�u��pb��S�B���-�����޼3�z�G�^$�脋 �WU��SR����c�ڸ	�9%��*���pg[.�ob
b]�,�q�P�JM)�ҝĮh1z�fL������;�q C�/"}`[z����-uy�������~�zڏ�w����$��8t�5M:��M�r8�m*T"W�8r�V �<7W��-ED|"+%� �<�
��_���蟿$��m���\�ʜq�ǡ?ې!�w�ډ˹����Fm���a���S�6�{.f��RP<䝻!�A�3����̉��$A���b�����'�.�2ݧ��6'��U���婰�9��k�>5�!s<7+��V?�6U����f���}�����?g�1@ՎOA�Y��/˘|1��h�,�ɚ��*ȓ�~+�=z�����sj�R��CM� j8����:�4u�3@����z-<Ey�n�
��ק������AKW/[;��ʑf��4�M�x�Rn��3��u���4s��{t"*7g^��l�f�dߒ-�]��][��u�~6��ʖU�X=s�NeQ�qLmЉ)�Z08�<c&0:&���0��l#�2�7���E�=C��o,�2X?��L����p����;���٫L�5��nE�P�ѵ�_>���g���]��˥y{��ؖ�5���^W��h���}w��>a}��,-���2\
)�ހ���D�A��s߮Ɣ�I���=���7�1y
yk��g�{(�r{�5�'���ʷ4/�+s�b5v��΀�ݩ�ޅ���U��s|mj␘�mB%*Uǣf#�k��l9K��X� ��U*S�Fu*���a��6�!3V3n�Z�.[���X�l{�a��cl:{�U�����qtؑ�k&���b6���K�9�p%�//a��ATo��w�Xˇkbq\���u�BX���KR��c�Иl%���DCrNĻ|�V�M��x*$��k�$.����:�x^�����f���\�q�Ln[2r��t5I�es:e���r1�g��9�͊K�|��_��;���ȓ�`�}k��S�ib�V=�9=��ڲ��@����߯�0��yfi�rfe��U�l�l�U[ִU�s`g�?3����o1�[�>S����u���g/_p��+pw��e2.z����>_A��b~�hj�,���w������3b߼��廼���u1("�jy<�\h��m@�������^��r�5֯M�5l��H��4�	 �������i���
;�y��J�0��-�I�|����t(U�>��ЧEzw�E��Ch?`-�!��`C����v��TKiC���4JoE�V餵�L�N]Hi�N�F�hӨ6m��Ӿdaz��_H8���O�>�i͸�����7����Mz�j�D��l��eZ�`����ip�)�ݗ��bu��� \�15�;���S���]�����j�(��|��\���S�B�WBޛ7��g�<�����f�yF�%���N���Y���H�����8d yk�µ�@\����9���s�d�����t��+��\%�%�3�>�Zu�ӤILX���Ӧ0s�Rf,[���Y��8��`��m�ڳ�g�q��~��YŲ]�Xw�Kw��E�8w6?.���]�c�����ɝiԽ���V�IT�ԑ��Q�mS"k�¶X슋;��&�Z|+U�)��b����(\��
oP��Z��uSv��zn��>�v�@��\���Y9!g&�r2Z�T
w:^/#��Xr>�����gI��n%�x�_
y�����Θx!R�3�l店��_�y��4Й��sz��>�/��k4�i�mZ����{�<�і/mQ{��%pen��,3�)�����gg}��yf��-F�B���ӧܺs� ��A��z
�_���9��*���yj�.����%�����Z�9�r�c⨑ˆF.�4�k��O7_���_��Ϗ�{�g<�5WB/R=�i�@�@�y��ݟ��^�8y��݇F�^�.C�I�oހ�-S�֎v-�ҨY*�Z��(W*%��MR(�(�����W_Ԥ%�[��&�Z57��J�N���ٍ���Ҵo7�z��k����֑qMS_�6c��2<*�i�j�E�?���Y^����A���l>,�(˂
u���DNm��ɥ���s��s�EW���-�Z2<����;��֗�ơ�������cLݵ��%OVk�f�{!����c�Ŋ�5Xc�g|�bv`0�kUgn����ۛ
i�qM��]|"�q	X�U���{��ؖ�L����K2`/�fc"�t�L�Ԓ��5s>O��½��ڿ�����n������;Y�yk6m�ȩs<x��'�f��m��ܕ[Y����b߅U�?3���9p�[6�`��!,];�%;v0s�N6�9��k��D�N�Z�(ٰ9	u"h�3���2�-�':1��|S�N��H�H�Q� Gc��ۋ�oھu⼅/���$��ƙ�.����N��'���n
^�:s���0�۵��؝�NH ���Pѧ�
i]*�1.�4;Q�l!qB�&b3�={%�������<30?�/��k4d���ff=�[�Դ/3����Tz�^�������OM+:	CA+���Si���gϸv�&.]�+�3���^_���)c�Wf�MV�3!�/C�������>���~��r&m4����^�����
T��C#o?{��3��o��CI� ��� ��xMܼi�* ��E[7��{ݻ-�\;�z�4� )R^�lҐf�Riܡ-�;t �U;ʥu�H�4�k7$o�FԪ�G��x$��/���8$T3�	xV��g�:����p�s�р�ZM��ۂ�)D7I���߾�лW'f���Q5�2�b=h�nϸ�I<�q��;�0�bC�������_��}�rl�&�mK�|�I���'�Þqi�f�����9���[����\�=�Ѭ��L �fF�?gU��	p	�K�{��:�ca媬��`w��h�¬I#�#�]�&��*a�T�r	�V��eBe��*o���,^�2q��k�D�	S�>m>}�,g���ݺ��'N����:ʹ��=u�5���v�.������ذ�0���e��l;x�������9|7���Y��Cy�SG�=�!o�w�Oaͺ��ܹ��+ֱi�q�.�A����6r<�G����[ع��2Z��Y[>���˽����kǐ=�?_GGcS�8!ŋӨ|S
�a_TI.��粍?�-�8+�v:�+'��ϙ�9���t��}k��e��b[���[1vUI��W������ؗ�ׂK����#�&�S�-z
t
x*#��y=����>N�Y���~��B^f)�e���t���]S��de����os���n����}
q:6.���V�S���{��Kׯ~v\�Y�z�s˿|1��6�x�9~����J��+I��߻͛̐����y7&O��_C��-�2���g�>�˝&�+�6g��Z;.�j��R%H��g0ͼi�D�w )���5w�1��鄋&�n4t�4���q�w�"hY�$m+%�!5�V]��ܾ�Z�$�v|���žz]�$U3���T�A����^�}��d��St97��:8Vi�CR]*��6�:���b�X�
�����u�^��r�M���ToB|Z3���s#ػ�	[�ff�JMNb�1��r�ׇ3�����������=z.II����.���͚�y������c�wa����bm�N�/˭В��f]����򌮷w�ӛ��׸�h3�+�Ct!����q#(���g�m�8\�UǹT%�N��BrŊǕ��u�DիGBZ�����Y��p[61�J�o����;Y�q'?.\��N]���̍ۘ�z��G���w�\F�Y��ً6m&#��`✅�^*��d=�7L���A<��9/^֓�k+o5��;1}ŏL�&.���E��a�6z������7o���=y�����_4�OF�z{���`鋕��M���)A�زt.Z�U����^ �ʏK߸p�['N�t�L.g2r�r���4	#�=W�;�3�h!��q�rnw��ŗS���YM�z�R�?�|*�MF�̉��<�+�X��h��}-�4~�5�!O��B����z��I���Y?�/�o3��������B\f�B6�^��Y�<�S��Y�j�ࣰ�ݙ�*�Ф�5~����h���[~+�oI1K�i^���7o�q�
g�_�J�U.\�̕k���]��ҧ�����Cq��L5b�?=����1A�e5�����e���r���K)�KZ,E�SiU��-^�9������=�����@�ĳ���k�`���s�7 @��_ɹp�+yGB�rΡ$�܊�\}�UkN_{?c}��������Js9���ًtk[�XY�$�M�=iE����,Z�z�j�8��S[S�Y*��5%�NS|�5�-�!�g6��3.Q �9�Uh�M����:�
�5��Z;�<j�3��U�b������|lc�43>�`�T�
�p�������=u�{�\�>�F��T=x��7c֜tFm���]X6f��������iܟ�U�sj���;ͫ�s��f�~���ȢZ��۾/�&������c8T'�ͅ���r=�8���Xټ\>'Iܜ�?6C��f*Z�����'<�8ř3Xѥ�z�f�`����1.�챵�,U��Ix�Vŵb2��$��X<�ɵ�һ3��/g��}L^���;w�`�
��Y�ҵ+ظcw�eҼ����!�W�l��ĥt�b۾48��=�S��j�Mb��B�=Di�g��-c�P�9��~�$^�����)��/��[�����Y�i�~����1}�a��8ʹ�5{*ۏ�����B��x���d�]�p��D�I��q�LZ�N&[�/��,��ŮpJ�.̰��,�(��H�gs1)�+gs���2,�9�͑�_�	:�;;�Ǥ��=��-�sn�8ܠ\��gB���sյ�����Z�;M��]sKGf��.[-�4Zq�����/���ife6z��d����k~N�c�5w����T�/D(�Q�f�+�o5�g�������
y�t�i���'\�q�3.q6�
W���ҵ��� @s��͛�y���Q �ZT��!��������j���w��|�	�>@�3��Z�����U��y�F�S��yZ4����Ԛ��YZ�=78�n<{��rݭW-#��^���Xᓟq�A��gxp>&�bb@Ac��`�@&�31"���х�U�	�ZP�aK�7L%�F=�*�l�8V��k���8��š|m9�k|\�9�:�e�)�[�jx׭#`W�h��S�6qհ)_�r5�B��}p�od�e�K�U3���Y�,���i��X�ñr�J�ѰME֮K�̙F8ـ�?�%!�"�ۦ1z�8f����f�Y���1!_]�������S�iaU����%X]�Y��YS����R���`Gp.�����eS�uQ���� OB��h�!��r��/f�I�;���m��H�UP<�\#����/%�ɝ�(pW�ڤ�H�n<C��eͱ�9{��;����LY���k61q��_��)���j�XbS;ת����R�6.	�l���m�m��F�pHJ��R*��S)֪�FN�������G���`�^��)��f(C$S���#H�;���5�Xw����R�[8���s��y�a�0���Fͭ�NM���qb��l�ՙ��n�	ºp_�Gc�?���h]� [s�2��}���gs�sD ︍'�s9s�k' ���X)����y%8ڠ�@�sSJ��s&�I�j̓+��W���i�0A���ԙ/^I�`���ά���;�����������3\����,�gU���at6�v�fdd|��J�s�,��C����Fӄ�S�9��[!��k�7<��'Rúy��n���뜻,�啛�V���U��l}����Q������pά��}\���}�<�Ѕ��i��T\��A�O�ywM�w��G��=���`���׼_�����s�XS��{]����߱ӷ2g\�p�.�c�a��ZXΆ�s"� ���^�8�F��zh	9_�s볫Ns~�Q�>u�P�Z]
%��3���V"[��|U:�oK�aQ�"�I}	�p,'�V��e�`Y<�b�(P�.�4'�m=��t���^�--�5�;]gL��܅4�7���V���qF/]B��M)�<��v�(�2ͰC'l����\�V���P$]�U���v\�Z��'��jx5��c�oڜ���ߥ'#�e��L�Q���2�-��~��a�_~��F�"*��E�Y,����6���
s8_�E�+0��-[H8]��W��i�(����ׯyt�V-g��ɔ��ǲu��x5���I����*Z��DܫUïjuʥ�a��MLټ�Qf1h��L^���V�v�8�����iKI:��=��ԩ;u��`��W�iI��u�������� �B�^�ZP�QM:S�iW�5�I��!4�;�U�G������"�+z�GΌ'�_;�����X�n'S%�FϚƨ��X�e�.}��?�[�����Y�@8�#�{���勡t�MvWr�#O�xr�%O�|*��r�l�*�y�p.���LNW��t會7'-��.�6��9KwNY�[�]{�1�=��p�x�?���\��������_�&41�!�hze�<3�}��߯�%�6g�U���*�}Y��0
L
0��=�Uz����<s�4����[�ά��Q}֧@�o���/%�	�)�)��y��r��-N\�,����W$�����ȸtM���ǘ��QV7������h8gVV�>���_��L��y��c��T�9K�g�<�{ڒg��7��������9�ءQfoh���*�������W8�v{B*��.�c�����m ��ݸ$�:���q�w �6�[��x�ԈÍ�3�Q[:V�G���W�*6��KX���D,G���Fk�}��X�ñT^	5	�{"k7�J�>T�ԃ�k�q��=foYΨE�l}�����Lپ�Y;1a�&߸��=�2m�&�l���}��i�/���Tiݒf��R�eJ֏cڂV<z2�����DU��L¾\9��X�o�ꓷns��mK�a��8��;6g~|)f�
��*8�eA^�qe]�'[���K@oox^v���h�Fs3� �"Xդ)\</������Z��g̬�@:z�$=G�"�E�1��.�V���S��ؗ��|�ִ9�^'Ҵ�R�g��LZ���Fдc���cfͧi�Q$�@ljoʤ�$�^K\��rm��_Y�Q�;���[��FD�oE�V���m�z�}���j�8:��Dk��i3h�����q��y��Dfp��\j�O%e�w��>�~#�1z�|��F����86l����o�\{6?�4��}����Ɂ<|:Z"oWlNƥt>��S�BI�,Ox/BT�R�ec���s�dןrs�O���{`�����m�+7Ni˞�3�r�s)�'�"�[v��C���=y���ό�D+n��
M�*#C��uh�f����.���4DY�?�LO������d�OMÙe�V� #�?��[֬�c�i�Дy���Y�!K�.�t2��;������~-�ݴ
w�������Wu�aވ�gV�iM�܋W����ç/��
xw�<�?�����9'3Lp�:|��N��ԙ��;{����p�|7o�6fɫ�B7�����z�~��d����kTY��g҇�Ԩ;t��κ6�G5�t����xej����R�=�P���o� �/��;׌O����\+�]�o%��}a:֞!)H���ٛW<~����W=����Nξ�$v:r�=��y9�"���IkO�rgONOX�p ���WcK��tmޞ�:)���Rq�
�*V��p��+��Cb9��c�
DVoBB��4<�N�g2a�:�����;o%���`��54��СՄ_���D�6Hl?����t����G�Yu�,K�a͑3�ٲ���v
$neʚU�u�y{�1d� -�1F|�5��T�V������n�sRK���%6��zu�ګ3����a}��$��������)X�]��"$��ؙ7�}a���d�_(���+���i��!����_�,���8��_����{L����xn�Up(_�r��7d�)\�z����6:�ą��;i6m��a��3�G}?�c�%o� VB�!�HǷz
^5��'�
v�qL��K�$�6&�S7���+��u�_d�+��>s�n�5t��S�I&v��E�:�Σ�f��חs��b��[�qt>qM���ڃ��ө�0ƍ��eS�|`%�6�g��q,X2�W�K���W?p��.�����xE:'nw�\��|��7����UL)rDE��`8E�3�zU�&V�B�r����[p%��r�������NX;rT���Ý�a�/U6���Ӂ������H�$Dsa����iH~�O����jS���~�&���eտ�1�������ܺf�g���Vݚ�oq����T��0���-#��������O<|��ۏ�z��'<{͍{�8s���T'Ngp��eΜ�ȩ��d{�ӧ�
�]���FZ�y?o>���K�>!Sl�,�����O��)�[��州3�{�ʏұ��V��h^���ޫݵ�Ԏwy������8ݵƸ�Wb�K�VnW�/����+�[��W���v�;¾��9T�'[u}X�@v�;	�yp�ʏ=�8��k7v��g�[AGWfo��L�۔�-RɗT���iΒ�1q9��'WQ�//`�ht�:��#�F}*w���e��� �Vn���3�d%��,�F۞D%5�p�tB+� �j:~UZ�U����Q����#)�6�J���~�b��ZK�né�a �; �YJ�mAŴ��ڛ���0.`��ĭ����h�s;��`*6�ýdE����5�9N�Mq�ڔ�kbS�6))4Ѓ��F�npV5�eA� �G�gwL��+Ɋ���ED�+� {B"���B
��y�@�S��#�3����fbS/�j�Nx$)�	�%�Ųt%Bj6�J�>�\��;��k�ju�O��f�~��t;�A�'0y�2��>����?mU� �yg<��
�50f��W��w��l�B�	㘻V���)���z��aj�
����0Gh��Z����.�o_�僋<~x���WѨ� J4�Lն}h�+�k��� �a�f�I�Ӈ:i�X�v�Ԓ��)<|;���Ry���<5�3׻�c�J�@�bI��@)���&WX��Q�,F�E^����&�zKv;����Zs�k;��t�rN�v昍#�s�r�cv��*�����%�����[蹜�,3�i�U�ө��-�*s��k%V������d�Ϭ�g|�}
�2+��Y�9�K��O���y}<3�e��[W[�tvm�ʈ��Z�i��kO���|J�����܊���s��x)����/^�@�{_�Q+dO$��4{��.\��i��=w�˗�s��%Ξ��;o���_�v���O��|l������yf鄄���W�?Z������G�X��j�P{�|4��2W��=4fwj�]��i{�����M����y�|�����5/��G����� �^{Ņ�pJ��]�g_sq�-.-<��׳u�V6�_�ֲ)lu*�^� �[�p�֓#�l��;��ÿ$[�VeM�fL��Bݸ$õTIlK�Ʈpilc��Z"�b��*UK�.1��P�GoRG�#}�4:�^D괹������p��׊�	����\oU�6�*�^���V�ʵ�Z���M��+޲a��X�%���ߜ��䭚&�f����glm9_�",W�#r��\��?�S��8�5k6��J�j�=�&9j���	TZV��׬A���9s,�f�aa�,)^�Q��Q�-��_�B��^��w�C�_��޼\��k O/�b��3޾|Ŏ}i�{�1�¢\ecZ�U\l�V����?{E�ve�	'T�X�6ThՕ����m��sc�d従��2�شv�u�M��k�&��_���ZQ�wfl�(�$�g�����L���"�6�L *�7��_��n���Q�1e��-/�>��������6м��ЍK7��]8|�;�&6�V�:�КQ?6d��N\��=�ϣ�%�q�i7f/o��e��� !5���|�X.�e����>,���
/���x6�G����&� ��Ł���\��e���u䠅�}�m��#J�j�2q� �8]_�T4h�d�/��������(X���|�A��tܝ�yZ j��	��I[�>�˚�},5�]`6Y�����k�����S�~���S���u���|�L��ͼ3��Z�~7$C�с�f}y�����u�\�[�b�m�]�ׯi��5�Hf�U3�.^���{Fk�p*�����u#�ܹg<Ku��¥Nv���>1u���V�������G�d(-c5�tF��E�_�P��I�w������?'P{�6�����ū�)��:w�k�nv�-���<9֍YF�kd�s2�}gt?����f;V����e5���|�nҼU��l�ָ\�S��%�ȯ�^�Y��&�$:}�{_����J�����ך���z י�H��ޣ������g\�tW��}�]{µO�u�5�����ҏ�ye����8'�9{�m���c�M6n;˺���n�N_�];�x����]7O���KϹ�4k/���D����3}�&�a�k8n	=��H���3��dVw���=�sb�.��ζ���Z�ݎ�촵�w^����:��aq�oª��U�&��W!�D<K�Ʀ��*�s�Ҹ���X ��q�SK�ʢ��X{����l��n�G�:�lY��&�I��E\���^@�!.�.�U���1]�S{���XEا&���X��q�p)�@�Nإ\K��]�ɵ	���_��r��h�!�4�gF�x�f��Z���f��5�m�\���s���l�%�(Y����,Y2��K��u"�
x�.2��1%������g�~.�b`!��V��%�h����
a���<7��ܵ��;��*�p�Ԁ��%a_�h-*Ըp�I���I����ш��Q*�%[�R�o_Z�F���{S�>y�{�&�X�o�����*ԧp�TF̙��};�sbg3IvWj�O��9S
���Yo$9���w������X��ǒbO]9��}K8e>��e��T������s��`��4�-{0{IG�����9�d
�/�B���4�2��;γ`�>"*T W�0l���/�7�a|U(��4�+��2���֟3-ſ|C�����|8��%;�����V���ƾl�lq��r�a�:u�k����?=���O$�<���>�N�a�~e.�%�E�1:NB�3���L�k}M��z����Kkx�=���:^ϋ�	X�pZ�{�J[VM�߈��5�L����l_�s�0���r�2��,���fh�Ij�R��Vik���j�SM�x��]��k��z���cG^�$���z��ó�=_����{���%N�4ƌ(� V?����<;��!gtI #,��+_�h׈Y&��B����Ib�IrN�ab*V�/%l����OҼs�Y&�2���w��^���6Sc;u�Q/+���8dT��w�[�O�CPO�4|���#I'O��6�%yKy�[5��)�@���z�>J��ٟMiXm�������|�[M����Җ������t.�ًWܸu�ݤ�;�{F�q���	�+�.^���wy�P*��L�Ɯ�2Ýr�(��5��铗ܺyO`�!m�z�!�Woc�.^�%Lt�MW��j)�������g���I	��Ռ{ub�H_K�Ը�F+e:���7<���K�:���d��]#C��ԕ�\{t�{�VH{*׿Tw� Fwh��b���<��oLߑ�w��nI�Db�������>���[�\��3���D{�d%�i�K�쮾�J�D�~�F�7��*�]��3�W�� 1�\����o����P_D��}y��8��{Ͽb��7���/<a硋�>p��/�y�q�o8���Wٲ�K֞a���L������1k��8fl'��aH���$��
�|����e���l�ɲu�Y����]��:;<c�;�����c�2z����B�����w.��-fܴ��v�}'_3k�)�Z��q�;}fd���������n�2��.!��l���ǀ�K��Z�^@Ǯ?�Z@�}�)�l�=��N�ǰ��n+�G��M�E�}5R�Ww �*w�Db+�ƦU>���T���s���[򞆆�\�1��GYu(1Ն�[o4>uS�^�7�N��m��Q`p
���d�u����sc���Lv��c G=9���2[Ox�cI�8f������ѥT2���#�L�EK�]S��áP,�x���U�<U۶g��u�t���{�2"��z���%�X��ڸU�o�=��U�⤟VM�cHa�W��7�2^	�x���_A���NHƫ\5��Vç\Mc�#V�����n�8.I�~����6\�דыې6}>?b�ᫌY���~ T��+Yմ�K�d+U��JcW���4`��ݔƂN�L/��ʘvE�dgޢl��.��<)��lNKȻ 	A�tSzȬL�'��d �=f��%�Mi�m�$�kc[�o�%P�e[��<�����k؊Iu)Z�)ś�S<�1Q�&��P�sbS;�خ/E[�&�Q\+�V�4�Y�q��֬����?�$5�F��QHI!�չ��=�ySN�[���>*m�ւ�Ԝ����/p��q.^?�?�@���Y��'�ߎ��ܸۖU��Ү{%�wH�R���Y��2�mЖ�}�0n�&�\Lb��oWr�Ƕ\q��S�hꕈ�SDq���x�N\�ԅ����ҕS6>�p`矲q�ʝٜ��m ���fߴ��x���Ru�Q����������k��������U/_J���z>��b��{#�F�$���)A�X��t�- �#��z�ʸW���}Y�5�W{�3Y���ޫ�r�J3o]��p��W���ou�s	W٪���[�b�f#�F��v�y}���YrJ�'r�L�/���m��{�٘�?�~�5�>����
�
:o�!���r���k�wR�=��7
/�\n��r��<-z���j�:�/���^�v���U�'��z(ר�F+���9�O��S��=���~�jL ��#�gzsZU|*��� P�Sխ���Ms|ͪ�qY�3�w��k,�q�C�ϰq�.�.[ς��ظa'������;S[�=zb�Ofh�,�ڒ�F����F��ٳ�9v�����c�<v������j�s8x�0��3֭�qu:�A��|��)ϟ��� ���O�Iz�.p|Z�>u�ѽ���5����u\�������۳�R��{�sf�Q���̆�}�*���IƮ�<�{.����#^\�ϐ0� �!atA��T`D�/�{d{����x*�����r��}9w�K{�r��Y�m�����8�rg����\�v�s;�pv�9����S�����g8����ʃZ��#k�v������y&m^��C�N���/��^9wt��/?�������/���\��=Kv�m�V�����f�`�������W�j�j�LZ.ZɊiY�pK�mgά-����a�ѡ�,��̢A��4�>�f}�R���7�F��~8�&�;ߌ2�[R�rg�U�H��iD�hD��M)P�˥S�9a����Eʷ"�@C�lb�`�֔I�J�2��,"�lD��M���]ԓ�����CDLb��!�p*E�^��H��@�j��,��kPM<B��Հ�-�.ז��m���Ϙ��F6�9�.I䍮M�F}i�6�
U�]���Z��M�;�:!E�%�*��Otc<�ᜯ.�A���L�'�"~���*� ��-��+�}�ݵ�I(^�:#	�1��J�pH�W|w�W�N�*�L�X�9U갣}?vvʒ��,��β"5�k��-�>��o-e����>�&�*�aT�Z�-_��R��nE�]�lQ��S��XD�"[h�+�`��m,?z�ik�3i�2FX�����
�д���z��p������[Ru�+70�Y����S���^*	�U���\[7�:�b�Mk�V2~s tN��[B���>��ͻݤ�ށ='�Q�MI<j5'�����w�ְ��iz�X@�6��ϪY�+��1S�_�$,�ç����Tv��cY��̎/������������-�^�|lh�\j0�%�4-yVV}�<9�|��c$��,/P������\����2m�A�vH��ɔm�Fl�6��ۄ��Z�XV"�xTH�F䭕BP�T���$�~ʶ�D���|�Q���M��H�Q�_ںa�K���eq�o��̅�ާ�a����e��X5~ˎ,�8�Y�jp�tuynW3ѾKN�`S����DVʯ��[\�қ0f�&,_L�����$gD(���s����)���x6�6ԩǩn]XY�Y�c�Yp�9�u.kˉo���Q����qn�V��<���׸wU
�y>~(�8��ݏ�B�M����~��k���ͤ�Xj�Z�k������&9>��^��z�\�v�����{C
a��K٭��oj��ލ��y��6�X�}t�t^�{(n�K����#���=���]�p�3w8u�Ԫ��y$���RX]���p�S��ܧ�g�޽���Gn�w�q�>ξ5&��y��nq��S�۞���ſ�]xEƩ�ܼn��M۫p�ܺW.¹��ɐ���?q��Od�x�u)o]|ml��������ݹ�����SZ/�Жw?��;w^��S��r�9���u~2�f���d�ug��|�񼳇��r���>W��5t��].��ս׸��&7��ʱ�\>.�ͤK�^r���y�ѽ9���<���g�8�X ��~���GY��{v]��q˅7�9�3g�rA������y�-ۮ�w�m�+��A�?��&;7f�}��=Ǎ����.O^�P����{׹}�
3�r��q.]>��+�(����q���p�?{`l����<xx�8~"&�^I�ɼ�5ʡC:?�o����]Þs�O�}�F�,����c����fL����شa���ȡÜ9u���.��t���ns]�u9s��1���e�\�$�u�]�w�a�Z֯]#~��5�V�z�R6o\˾�;9q���6m^�֭ٻo��w��g�~qZ��_Ο=i���m�7�}�v��7�5�;}�$�2N�s�vC�O������Ο9υ繴�GfoaQ�(���2�S��ś��b'6�ġ���O�̞Sٝ2���'���xv4ǎF߱��(�5͖FcY�l}���.p�"�R����Z�؜<������NwVTiŊ��WMcK��l�Չ-����� V7��ƴAll?�u���vg�ULcj\S�KlN�2�i[��r�I�m��t�wÈ�)S��%0�tSC}J6�k��ƹ^e�гl��l@�RhW�-�W�e�*���D%R7�,5��Q)��ա{�^4�ݖĸĖo@��;�fw�T�K��nK�G\���/ג�B5(�؄��݈O�Nh�x��/�,�yc�
.�s@q��~�|q���7�y��=����/_q�O�28��տ(!��c�w�+�{@������;�H���O`dyBc�Ο�k@)��J���_Y���`�Zи�'���\yBb��=e��(�[hi����}1,�H�zM��RK@��<+Jޡ�<?�����[ϰ�8�)�(�yK�Y���,�t1|��%2�?G$P�9�Ǟ��{��O\����,�ԝ���?�S#�+��[�5�2'��p̫�܋�ί[�K��>��d��<�����������UE�XW�	�6�w���*�� �����.���p.�@���S��h��,:z�A��S�I��c�r`���{R5�5mɫ-�K@����)Ĺ'T5�ȹW�����{�����!�>��u��?��ZF#�])�U�{9N�f|��=�
N��O(!�S��4�؜�W�	�Leٚ���C		�
Mq+W���Z�g�lfn���=��2c"����"��pVc��+A�fU����7e��$֬�����+[�=a%9�7��Q\���6�p65n� ���Wd�zyZ��x�	�G�HPr=�*�T��el�B�M��`���m՞��d�'קD�
�nJ����\�j��hŃbk�^�.�U]�R2�;��m6�1����i��s!
�;���:��g�ǐg���}5����#t�nS7��q�t?�L���rU��n�Q��8���MlL�@�s|�qqؔ+K��T�o���;)V�����"E���?�{����+2ǯ��b��"���c^xI6�v�X6����#�oNN�ɍCy�ֿ��cZ��o7��}f0��F���=�g��iL0��N$��g3c�j��3�����3���2~�f�_Ŭ	+�4d.c�L5��s"úO`h�q��#{�gL�	��>�]��}�),���U��3���Ў���j0m�w�m�^�HƠ�bG�Ɍ�9�aݦ0����o?�q�fʳ�ɳ���S�u"c��04H�۫�H&N���9�7a���gP�Qti?����n8�;�b`���4���ܼ/���Y�tJF�X2|ݪ�%���܎΍{�+m0�[�c����L��mdە�Х��7�Oz��tl�_��O��=IM�D��δ�.���F�J��Q�;���k�n�k6�A-�0 u�[��OZ���Eϴ��<��Naloy����TK�E�tҫ��M�Nt�ՕV�6�ԝm�t��6+��qB�UhN���5OhJ�
�IIhHKQZ|C��Aj�:�/ۀ��i]>�����eyyO)��ƦS�H}*���jB���T.ۘ�Ek�X���P�U��Ԑk�jS+1��[Q96��	m��܍�5{�T.���M�T���4�J������M(X����hӤKf.���}�9���vs��~��˞[�&��ڳg�a������r��Ξ?����'Ǉ���=�qVe\8����ۗ�y#��W�0�P:h�v��NÎ�{7�a�RV��Ϻu�X�~	[6�`۶��v�����vn���m�8|x�{;"��N�����?zP��wX/ �ڸwͪ%�v떵b�v�X/��e�lڸB��r��.N���_N����[龞۽K��ؿ�];7�o�6����;ع{#��lbρmƱB��M�7	쉛W�^ƪŋY7k1����o���W�!�I�˛�ؠ���������H������ڌ�[��!UP��~��`��7��r>�� E,�S�&�*NE[�k*teS���,Ԙ�%뱢T-V��Ϊ�Y_��`ڒ���JmX'itu�tVTKg� ��&}�Q��K֡DyZF����I���4 j&���n#��[ -���X�E-rx��g!I��0��}
�$�M��hK#�yKS?���*8���E9Q���n;��5[Q�H2Ŋ�$�b:EZQ@�z����oK����GU�)AD�8
.CxX4��yqr	��-{���p���3@~���??�^�x�F����O>|众�({W?l�|p�͋�O(�~a��{���勭����`�zw0{�@�M�gػ�biDn� �<�����k�r�`!�nA��{=��w�7�W�+R6���Hl��ecel�<�Y^�����p���-�����58ʐ����%�=���\����C�w�k��B�/%�J�M���mB��6�U�Ȁ�X�]�C�A����o8�M��p:w'�ys�ҏ�l����<�l�dK�
���_�!c*7�Q���/�E�"�
�*���bS�h�&�~�&8L�^C����}�F�.Z�<%�aS��� �������)�<شʧRm���s\5��VaϻR#��6!�ZSc�E`�&�'7�K��Y�1���j��B�]b��`��^%|���P�"���}[�/�D��5�W����I��bk�܀��Q�����-�0cQ����LL����цCgz��P���cݡ,�ֆEj��L2�
��XP4��<#�,l��˟�<!� m7�~�F�5.W�D�*W�*��eb��چ�	=O¥Ln��T?�ļ����+V7�<�ý�!��ţ�V;�c����t��1�C��^�Rғ�k��X�G�Oen���;�����vj���bt��1�IS�S鸦�����l^�����](^� v����W���K�� M��4cVM���~f��38ܘik��B���Dh$�bX/5�%���u �{�cm�8���؟�p�+��5�s{q�>�C^���"��֡Y1l�<��b�XJ2��4�ZV��x��+K���$�b@1����d����P�P	�(��DRλ��Q��.`��W��1���O�W��m���Ԓ�aE�p5Ηs�G�t
ZR�.����v��B`�+�2������r�K��V�����6^��S�"�����S��:H �
�v�Y�P�;�8�߲>(,~PL2l�_����A�
 Z2��V>�
��(�]�)�BaW��9���~�[y�(��RD2�'?"�(��Li�����!�ӟ�^�T����եvY�=����T�񠚳/�\�����}�,	��S^CI�/5��\;��ĭ����w�����P��'q����:P�ƞ��v�wp�D+���CK[b��(�Ӓ���$��oV������Htv1~�`�@e[�m]�l�$ry�dk�Z��,Ϯd�E+'"���MN���$ {6|�+~�HӸR�L*O��P�3B�����'�����OBd	����$�şH;"m\�g�L����݈�?w	�]�L1��ߍdΔ	̜2��?���y�Y�t)Ӧ����c�1m*[6�3�k׮5DK�7g������ؾe9�m����?��6
��g��m���}�*CG	(�ɡ�ٺykW�c�������X�����n�����mټ�8^�f�n۷�c��E�d�8�G`s�<W��w3�w�7�d��E�Z>�Kg�r�<���l޼�p�n�x۶�,[6�~������;���������c���m�ٽR�0���p`�zy�M9��â}7�U~߹o���a��լZ3��+g�r��φE,_;�)�G1i�H&OA�vi��I����	�Qx���R7(��>yI�º����R $����CO*�y�,�������$I�//i����#0�Nc6�����XӶK����y��9�Z4gI�4��l���,kڑm���>�k[vcW��������ڴ)H��E$�*&@W����$Ĕ`T�ahݝ�~Q�˹ʑ��(�����΂#��)F?bĭłC%_���_����×hO?�z���C�|����#�[K��߷4�~�	I�^��ʻ �>��6GIön�;~8x���掣�#v���=q�|�Eҁ��G/����ܰ�v!��#6�&2���Q�s7�ϝ�'G��\Mv�3�]�L��ya+����{{�&���o.��"_�����M���$os�|��+o� ��7W_<$�s ut���]@P��&��#_g�CN���a���l�w�g�vZ��`e�KNorZ�b�$�J.K/,�}���.�I�7���]rr#B�q�"5����R�Y��2���r�-�C9�8��-��#W�����9��3�s��-�k,�����|	ù�K��R=�'���j)T*Z��E��^�(vQ��\H�Ԣ���3���it�~�����q��<(�|2�	�񩒆c|}��ĹL���ͪ]��,�m��On�SՆ�wg�kZ�Śu�z���=F|πI�={>��[Ș9�>}����nǞ$��FՎ�(�։�z)�9��=m�s���W�����ílY�+�#�Z��K�+_�M�Ԇ"]�/�!_EW�E*�:���w㘸l:�'tg�>;֒3g��u�kU��umhۿ	���z��W���/�#˳�7�9���E��@��  ]w���8W�N��ȝX��.PDH�g�e费��nDx�B�U�k��t��W��B��p�P����&7�˔9���G��Λg O��6����u��ˢ�v�ǐ�A���L��U�A�_���%4�Ԃ<!�8-B`R$�����S�2�)�m�
�X���e�-����p/Q����$g���Wt��gyd��W���l�֏ݺ3[~ߖ͎3_�q$����q2�3gr�q�.��dC�BI�ZW3�P����H`��S����#5�ꁒ)�ER�7�؏�̠�S���.A���`.
�t����q\�)Д��{S(�@��� ����N���B�Hng�[�R�3�$qG	k7
�v0T �����Xȱ�ʊٹ��P(��<G�M2ݖ+e�OTnW�r��Z�PO������e7�׌.M����&2�=ѹ�)d�FW
[yȱ#Q9�	���P�7&��}A���e������|���Mn"�
�9K�oO���l	�6~�?D��3E��S*ON*�ِlgOuQeK���CM��V$����f'!W.���I�l�(%�TZ�KU2��$�*����-�ÖٲS<�W��}�g
}�����ƾ�|�o�d����9�Q曯(�՟(%ۂ���B9�Dq��)��[J���r���;r� )G @�*�3̪�+7UrX�N��C��%�-ɟ�+"���|��H�o��"��hZ4��C��o�-!�{hο�/����@jP0�mț37��m)`m#`m)�`A��y����pWn[�)���è��a4���g޴�,�5�%�g�l�l��0��F3s�d�m_��=+��d�d/�ĚU3:�o-�o��=���Ƿ�o�Z��X��m�Wp��F�Ο�é����{w�o�nx[#�X'ׯeӖU�i�ڮ���3�][�"�n]n���=��p��Ny�fî�{�+�޹�8>zL@p�zq�*C��Z�������N&��Nƅ=R�>�������s��y�w�4�]8����s��Q�q�\?��+8wy/�r��A�_���s�9vrGOl��)���k�t{O�e����ۗ�Po�]�(�)��ߙR�Δ�t�aG1OW���Q�ӗ�~�p�H�3%�܈��
 )�/e��)�dC��/��})��I� o��)��ƍX٬	+6dC�VH���~]7n��ƍYT�1�k5eiͦ,�ٌ%��Dʀ��M�^+�u՚1�hy҃#���!4���b����5��i]��J��;|�RB��kB�I���(�!y���57��z�փRe�$�
RI�Ur���T����n#�V�)�����)�W`9��#�t��%�h���q���wO�\]�����:��R���㌝���Tt%?��
�Mn�H���[,���H�Rar�q�E��.��!�\���<R�w7:�	�IeP!���S��N���vR��瘯U9ظ�]��J���i+ϲ�}�6^XY��]�#�7�X��<��}+n���<d�aǟ�lI.ɷr�p����['��l���mn�[z�u���)��ǃ��|�����G?�8d���>ބ��bW��k�bJ��L�[�eUX�����.�.)c��Zw^E�"��5RN-���D��YX�SJĳ�I;5�D�b�(R���B�p�,nL��,P��J�(�ږ�CG�j�0R�d���Q�Ȫp)]���p��#US�$����&��9��*c�LP�f�jݕ���g�"fm9��K���'��~ă�O���/���ƾ�N?r�b��,�w��6�a�\j�KL�.�>-����X	l�Y����	5�CޜV-�%r	��ׂ
��mh#������V��ՓT^�h±�����۔!�R9Z��ac�ܪ�JT�Zhᄂ,KI���+r����YFw����]��"�\����c�,�%�Қ�B��:��M�G�o�o��8�M0��3+B(3�V#���d����:���/-xO^�x8n��<Y�Jg�d�a,� �2;�x斺��?�<�E�DC�2���M3��{�����5S�Y�4��#ƥk�YL޷L8~e�(\-�BɅ�*]H�>��s��;'�#,Q�e[�?��=4Hj��4��dzpa~��΢�Y�Ҋ�i�,	�d��d�7���ƨ�����<����f��/���:�#���Q�u���/u�|��De� �%SN�n�_ ��@\\�o�X�
i��L�W�r���A����rO!��<���mA��������|���_qwww%�@HHBHBpwwwwki�K��;�+�
mi��Z�����|g/.=�����^�����avgwgg�ڝy�wL��m����� E�������v-??j
(eػ`����M��Z��zkeO��=}ڷa��d���3�����M�Zu�&	���477;�$�,o_��m	66%��NS��^!��Y��oi���	!�D�ې��F��'�ǇD7��	��#L��ɾ� ��J%�,w��އ�V��w��L��:r����
��tv!�Q �҆4;gMI�v�H\��,�3� I��l���"�Ԝ(���W��r�D{�E	r_�Җl�*�8�l%�Z8�`�Ε��M�fc.�$�Z�4�5Q���ac�Z���NdۺR��U`�[�އ��+�FW������)hˑ�&���d;w�^7�]�����H��u"�Hw�s�$Kª.Z� n�<�;;b���`�{�{�+�]��[��q��<}t�'�/h�S>}������on��l����ܿw���Ν�d�7������r�:�����{����m�����>|pQ;NI�-�t���v�47��;�~���r���t�k�?�)g8�A�_}���>�������C�;{�˿�=��^�/~��O���4�4@���S�����ws?��ڕ����E����ϯ��ٯ��xq��O~����/��U����{������n�;��<C%����Oܑg���3�y�+�)8���ؾ�9�)	�,J@H`�8&V�.F�.��0)��Q�}�����Տ��Q\��%�&1Y�
	�� S��22�n�̍��`j1���E|�%��HJ���?�GkUr8��c�8Y�1f�����(�@j'�q�F1[j��~n>��1)�3r��M��B6O�ͺ��ϰ�d&ŧ25%��iՙ(@8�Z*�S_���=�Z:3�R�,i��d���2#,����xG��1�
+X3j��[��M�j��P@`LB�8�O�W!~!�J��!iY�oAR���W
�^.
��4�
����)\�����n��7y8x(`����:V@P�n����{�C�������l炃�Jζn�y:��b�m�[�bma���9�f�8JZic낕�6.X۹�\4k[{,�m��q�s�c\�wp�F�bi㎅��&s)4�K�g)邭�	�.�9�b,i��5P�h��ļ��G	��f�ۋ����*�D�(�t��Ʋm�.|�����˷rv�¦����e�X��}��`���/hʆzm��{4��w &-�`<��d�Ҳ𫞏w^1���hޞ�^��iѕزV���&�i7R��Ӛ��jٔV�5���w�PղAU���L|�N��܋ޓg�`�&N|��6��ְ��/�>~�u�g�(�M�����3��?�rO8A遰Ǐ�ns��9V8����1�j���}$	=��]Օ��	h�\�O��mGTIj6-���b��О�_�����'���A�~��G/�9��_�jx)E����&��@:N�����r�sO�*K^|mN�$r�y"~�r�~��ܴ>����7ħ�1���R4|�CFi��	�^%��א�(�Ko�Y�~���(���fo����j6;��K�
�cqz�)K�a�.`oZ����(+�yʚh�)�&���g�[�,O_����s),!��>�y��u�b�֎l=<��r��_O{��{� �kBK�⑝�ezM,$�2���$�iiLΨ�Ѭz�H�=)����i��,��S������s'�p�C ��QJs'�Y��ۡ�L�Rh��:Hɲeh�������r s����!~�����y����� _�
Ԅ��?���T�t%?�_�̇/6��8�u���M��-�N%�
Np\pD�.N�j�y����e��
8
�X�jkK��rR cK�$��V�lӜ��M��)��@Q�&�DH��!`Y# �0KsB-̨�⬹�:�MM4���#a������y�V�x���??s3�J[�g���1^�&���J�$�՝��\���a�F�����t%X�giO�Θ0�8/��@33Mj�W��16��T�-�2���56�Kg��N�#���n�z[�eb���%β�!	���-�&����
��XS���ziב{�p01�Ps+BL�	5��`dN�������ݔ(+���Ĉ�Nd�H���.rO��[9�ofE�@pf`0i��DHfhf/�����0[-��TD�I<b|l9�u�|)�x�T`���_��_�:�����A
�y��{n�����׶�=z$`�X�M���|�������ܼ��H
���_A����Ww0E��� �����۝ܸ}^��s��:��G|���~��Qm���c��MIYה�M��N�rն���p�$�?��
����Qӽ����_>/	���=����?K�~%�J
`�	�*�T=j7o��x���_��o����&�~]���o_i��S�E�q��q���5Ƕ��C^�@Y�fk$�D��(ڇ��^
���b�(�^
ZJ�¢������%2,8��Q�V��O�d��[c��X�U�}��""�Ϝ�9��I�tm���1�R��P@&'�r�&��#	�8�^��j��M�HD&�T�ž�Z��� =��X�Q�2ф�E?�='35�.+�
Y�Z�)5x?�:K�&��RX���Y�V��2�&��j�>9�Չ9����Z�����L�c�\�~#i�[�Y���^=Bp���� �S�)X ���/w|}�|�w��%w;���p�� �M ����Wr�tԀ�U����)��IA�]��U
[v�8XZ�" �b��H�_�^�7�J��N����[�1sԶ��q�������R��V�����s
�k,�L[)P��	��qƒn�K<�������ɵ-���d&�[;h��YZa-i�N��Y:k�����א��Z�i��+��C��7X�g���6ZFf�y��1�.��ß�ɡӜ��[�o��O���]��o�r��u���67����=���v		�J~� �F-�j��WPJD��$�5&��a�M��\�??�a"���a�4�����6�+lH�Xގ�v��Rv?��KW�6��E�@����&SC7��L뽮��/�4��je�6�����C�^ȟ��f�ҳ�R���{�;s�	6S�b�aM{ܨ��'o�v5'�����H:4��O�u� ���i[q{I��/�^N��+��>]k^�tžn}��oøys�3�=.��q���]�����]�����M{��s��ѿ\bU+M��f���	�j�OqC��DU�'�Q���'�m
z���`�[u#ZH���hn�Ǖ���A��� �E�y�����_�Ph L��PK5ԅj�'����#qw~r��.��*
���ݜ'N�ʃ5�u�'4�D�:D���_jɱ�r1I��1� ��\$����q��pvf��7����XՎ��^̲�rvK"pF>�c�����)�/u��f"X:�%1�a��D����t󋢩g y�ex
�
���<��u�s��rӬieJ	OYe�[�Ń|I�r���v�ֶk��c\����fk�)�ޞ$G�b��z����E��� (+�R��WJ��"U�S��[�=<�ܸC{�#=*J@(K������E���^�#	��PG��:#MmJA��yI�#s�m��:WJ�F&8�)�HX���yJx^"w���^�Q���lߐ�+�و��XK��������+)?�l��u��d.�&��\���ò���a/�(9*W�`#��d'�k/�Q��"2<'����?�Y�W��"�H�o��g�����;yf��k��3S���b����`tYR�+<y�3��	���Q��Ǐ~Ѥ`FYخ^��K�O�{���ՠG�%/�X���fSR����U�Bv��	�7�	 �����Z�
��������뢀�O�)����լw+޹�pV NY�~��K�WZ;��gO�M�/�'@w��)Ν;ŷ�ʹ�^���o�$pz�����a[�G���g�Tu��[7�>n�u[����z�������_W����?qS�!P{]`��O�r��q�����f�����T�F%�4&����| ��;�:�e{{X<��8����F_$�r2�G���\ֿJ����g�ڼ��dds�Z&�|c���G	|����,���ax:$]R:(a|���Q��(�����cs9����|v��O�aSf���-�6{��h�+[���(���۵�.���RX-��\��k�4Q�E�o}V.�ꔲ����Y���{��3s5�M�ɬ�,f�3�q7V�A��x;`o�7�z����� �+�n�~o� �J4�3T�<g<��p��Ҏur������7)pRr�u���啜�xr���}68I��,�A
�쬕ߐ3����le]���A2K)xd8���;�'g���|�o�ZI����3��$�U�������lL�k�Z���F�>�J:ca)��!�K3�
� �NJi9=�՛�u�2l�W��ڎY�ZRZ,d���l���5��杍,���USװq�*֏]̻���P��9��^���i8�`���î���!u�T�B�
"�*+jHPa3��_REXESm���6�6�(l�^�6��-~u��i�J:�c��}\�qOc7%Us���}��k)��f2�+��)�z�O_/���_�~��U{2��E42����U3m�d��ed�_�
��Hd:��yka��<|6�ۏ's������9�h6�?�:� ��)�����0��6���ߍ�����El-n��F��ᅂ�]t?\�H��ߴ�6t`���4�DLӎ��=���S�ی��fx�,;נѕ���jC���ԗ�杩�m8�m��O������\���T=���EY��w�*�#kd�B�U/���Ŏ���t�p>�u8�_����B�ʣ�]���/�������A���,�*�&5�qJ��*$�_�>��MO�7�-~���ò^C�;v<�er��I$�;Id�v��3�'���y��a�PF��$	K��>��!�yQ�CU��hV;U]���U�e:{����Zi�n�HIO)U�t'2�u\���vL�$XI�0U��GU/FJ�3��B�f�J"lj�ImG��I9&�ҖX�8)M* TЗ�(a�	��X�d/�'��6?3+��g@׾yq��I�ce�Uɾ<��H)�[*ȳ"��?�2_�%�.�\�)p{S�QR@�`*�b�����^G��r����tX�a!�
�,$\����Z�1�R�m!a*�����s s,��c! e)���H\	��â^o��' S��rm-��*(S@� �^�`�Fd'�*�{W�C��haF� �A�8Ja�J�K�o��/a��D�=�mظq!/��Ɠg?�-L��40��ϥT��TӃڃK�X�sW�K ��cUuyE��i��GJ?k`v��9M�:�t뷋w�y]��7�q˙��T�/<y��o���o<������9���^�_r����x�K�W���3�W����5���W��×��]��{��6Ϟ����-MO����^��%i�M�xqM>g�{���_���kܗ�<���O�iz��*O�K������=���{���ϸz�+��x��T0(:�)��4���T)@
�lI�aGJ6;�2�����:���j\-�!)hK��t8��6����,f�`VMve䲻F��J�]���9�ȩ��Z��̫Ǯ�2�H�5��-�)�ȯd_��씌vgIv���`UWv7�̖F��ܤ#;�gwö|آ;w`]U'�I����$V���f�$���m�A���ӡ���b{�V�kۍ�����P�v�ͲV�XФ+�ug]�>�ח����D�����Si[؂T��`)h�������Wh:n)x����p�SU��Zu�����z��{��A�ms��I�G����U�'P&@���&I��,-Df�eom�����@���y���h��ϐ>X��X����
Skl�%L�������䛴���\�O)�)�3������s+̌͵0�Ll0�0�Lĵ���S�5F:L$�2�8I|�S't&�R0��<3��LN&�� t�W`�`-���5؋Y�f2۬`��]l|W�n�;,������إ,W�E�����=8X���	4��FPH���'�T��|�S�\����J��}��-��J�~{�%��+÷�D�N�O /�~G�k����
�:����Ӫ����45ڷ�ʒ����7k���O�����D�����8}�k>��k����Y���|�\B�:��4�ۄ����^L�����l'|ޙ���0Ꝇ�XNY�F4��_�*�~����jG[�r�8�-kKB�Z4ۓ󗰹����o��8��[{`�=�Ը�6�FHeS��ub�N����lчЂ��iNtim
35^\X�FķhOL�|��^����a'o����M3u�����]��Ð*��V>U�LU�<��/	����:����-%�֎�Y����ON.!%Ed�mMv�����ᒛ�sV-��2��HD����#�X�>�V�G2 CJ�������l������s0_�qY��=����U>�L�xg72]|�)	R��ٮd{8S�Ǖt78WO�]<4i�,_)Q .��I��&��M[O�d5'M����7۾�[�la�UG�%ՕaR�S�+	Z��X��9��x)��9.J�U�����5�T4a`��D�j`$@!a�K��@Π@�HUM��JuJj�G�� o0e�sS`����� yN- � =��e��)i�9��;+����%� e�3H��=S	�X��w256���~��rm�����l��^�B��<�LEƚ��R�S���u��+9ɳQ2X)R�(����`wO͒�jf+Ph&q��dl���ձ�8+3S�����c��E<~��V��S=�<y���|5�D�z$ߔ��w�' ��H��������Y�n��Q��;��챂�뚫�Ͱ������� �e_�!��\����v̳�7e�!�%N
/��5������_I���i͊���o�����7���r��Z�yKU1_��T�����HZ��./_�������ڇ�e[��L�?�ǋ�z=~t�'�o���-��;=�)�{*P�쏛����%��Ʒ�]䇫��v��|v�I��0��.��*S����1�Ikf5j���f�(mʜ��kҁy-:�V�v�ۺK��eM���c �:���N�Xгs�wc~�,�އ彆���q��~������~#X;`���X�t�B)�/�=����1����>�wz�eٰ�,>��C�1g�x��!��;r,��&Wv������X2x6�{Nb^����<��]�1��@�4��Ȇ]��z cZ�gl�!�� �����=�1��X��H��}�q��v�s�FT&զ,�y�E$�-�^��uz��ו����&��$験�%���Z���JN6�ث�nVN\6b�r��H��Z��^ҷ�x{S�i��Fd#H[)`�p%�t�����&W{<����J��.�niNR0v?�4�����rݍmp6���68�����b%��*�"y��{ N�!�{�c�W*v����4�z'c界�o�>zY�󫇇Mwb��S��JI':w�@�:L*7c]�]�~���Z�`�ml�������<��cVɻ0��G���x�u�9M�EB`>>8�F᚜"���G�:��	��k����s��|�����:exܹj�eN�Kq+nF@Y[|�ʨ+��՛9sI�����'�$-��W����FyS����Η��	P^8�#_��
5;����Gp���p=�m���igN����z{-�����C�V$V6"��m��f�t��LI���nӒc�r��T~�9�iۊ�<�&3'�g��	웿�'�����4c"�	j�R0�mwr�$�eww$�~��!��A�@�+��X OܰF-�ߘ�]�6k�Y����yk^>�C��,yjQ#ǫW���b���Ч��O��C��T�TU����6p��d�_M��ͨl݁����PLpa>	�_՘��zxժ�[V.^�5p���.:[?
E��'p�7��~1��dN����r-[��O(��{r�Ɲ�� �[(=uF$H���B� \�f��$K�)�͉TwG���I�3(Q��+%�;k�"�Ժ�4�&JJ��SD���;�'�u���0���5#���p�������B��3�\\�&��X[{=����
O�a���I����5�5n��5q��Z��8g"0�T���
Q�ieM���&o�N%���[��NU�*iP�
nR~�S�� ��X � ���C�����NUe*WUc� H/e=�����A�1T�*롣������T�����$��$����&sUm��@����2����Kk|$��z%w+�<4I&�ll���!�??�Լ�p�w#�х yW������;[S���8��z��vF�?��nz��DU5�x�P��>O�����A��Mz��.]VU�����s���4)k��w^� �����M)p�'	��אǟz�{��f���2	`�s����� xW.}-:��ˆ���s/qߐ����W9N����I2�X<����Iӿ��:�Ͽ��Q���j̭o�����MI=�'��t�ޖB�]9G@P�_�)0+�+�*\Um{��~��=ߜ:¢q�������
|)��4x���aÀ	l0��#gsp�6�{�5�f�e������d�ۋ�6�v̜ˎ��c���l��6�f�c����=s�e}��Yr޻�7�}3s���5m=��çj���^����X#��0m1[g���W�q��O|�S�e�Elzk!s��b�@���Ù�U�a�,V�����X�o
���Č�۪?�Z�gN�QLm5����N�1��m,�z����X�3�������-{1�YW:�UR;�&i���v%����𪚅s�Lm����=�q�|����G�����zڻ���ݝ�p�o���������	7Mʲgo�鵅�D.��V��8:�bk�)��dg鉳���jd����G��S��7�m�q����qv���-�DmL=��xMj��<�r	H� (C�6���=������j��_�?~����KS@N?�k�B�7���v�K�� Oo�� *w��-����ێ�b/��7��x)#�od�;[�0�V�X��Q0��FVug͈��6��u�P���*�CCq��j�֞�3���R�
�4�)�\��m��[�s�̪�uv>���)З_�:��r�~�>�|^�$�W�w�P3	��S�]+x�D��o@���t���H���)�����ߜ�����>5�Х;O���%���W�ǂD�w�m�gQ{j�K���n͆΢�ؙ4�Q})p�oKہ�xkn#N|Տ�#m�2�S����G����}�Ы����=�
Y��ħv;B�u!K�;�Q7��[P����[L@�RBK�YVEl��6h�uƈ�Rc��38xN��U��aR9?ѻ)b��W�o,��U?���N^��
���ߧ��H\U���9�����<��o�}w!��X��]=�^?��M�ӡq�+).�g�H+mx��GS�gFu�bb0�	�:��x7W��Ʊ/1��a�,
�glbu�L���s�'.������ݓ�����?g<�x�ƃ�ч
|�8:b� �fK��%���GX�j��HId��E�Z�g������ӫ*P�(K�T�h��C%Ue���)ȋ�K��"�ӝhg�%����'�x���C5w�n��N����#���DI � �H��'-�7�Jj\
�����.�Z�؅) |%�^)H@DI��[Xj`�!���_@%P����N���?Þ��Q����L��Tղ�ZUY�U���VY�,�� OY�Ե\L�q53��B����:3����bV�ڪ�H��^�Z���X+�jp���RdN���	qf���Ȅj��ȵ�%�hSk����D~6�x�*Hs���zۙ[�"Ǹ�{�)����+�n�9;
�Y���+�jr�0|��514���h|l���L)��O����������ņ�� ����/����Z��*I*z����;�_�ƍ��zEM�u��U��|�_� x)��'���Ѫm�%OY��iz���?h=[�����֪̾UA
l�,n/�T{����Zz�~�J�˿�}�]��uw�	p���PR�}[�-����M�g7��h��NI��HY�T5�_	���u_H��S��/��}͊�Zr_/��x
�����]�~Gt[�����U~{p�_�\ಀ�����s/�6��Ѫ^���hy>�ߑC�9Rу#zr�� N���f}�D@�T�����j3���j���y�~�n1�3m�M�a|�y(����~�D#8�{'zO��i�ɚ�a�|�y��L�A�8�w���L��K�~��H��3�/{O��Y�4`':ck�~��.�&�˖^c��Eo�5�8����΃9ض�6�G�zpT�O;�����4�}G����V=8(@w����t�Dyo���cަ[Q�@�]SH,�Cl�8��&b]���U�6X�o�x��K���"�՟po�\�	q��O�.8o'W|�<p�w�E
֮ξ������GN8������k�6���} N!�y��%a商�_6��y8����'W$��)W���U@MlB�+�>���r<������v����1�V)�J�Mfwjt�-����G��oͮ�����S���-��b�e`Sw)V�����zKq����˰+yG��žd>F�Wj �3��)5��'i���$L]�6Mu�`\���u$Ţ��U,���eCf�p�f��A��jЉ�f2��0�R�gg�Yb�))8'�▕�OA=|��Q���r�+5�3�߼\j��<5���8�*D���g�Rjw�Ɏ'��H
���h����Z�+��y��2X�����������sZ͝}��%��.�����PIM� �>������SҨ��V'"*:ܨ�6������@�D�A(�ߋ���)0��^�(�Й��ڲdg_�\�ƺ�L����Ms�K�G���f<u=�	�T]T@reC2��"����|�,�[Wpi}��*�j�T랬>�jNdejw���=$9��������f��$^���ey�G1���QR~zU�����I�U'm]�vs��r��2�ƽè�Ҝ�ޣ����jR�DJ�����W+Ϭlb����&8�@� :%���f������x����w�r�Y;6IsH2��%�=o�&��m��WW>�$�UU꣪P��		`Q�wH0}-wZէ�fU�A
씴ޘ*��&��A�&����"��B뭪z|��ZU}�����YZi�bb����i��jKghS�klI��`[5h���cH�M�W]�Z²��_��'�e��i��t�W�zm��U���\�u���)ޛp��ՓoJ_M���RemS���)+��nM�:/�
�)�Tm�|d_��N�IG��N�Y'������c
M�w0����\�+r�Qꥣ�CG��9��M(�2����z�_᧣*HG�c*|d[T_��uի�QG��S[��dDu�����fI���7'�\�#WYUG���o��h��0����&U�+p�*���G|h�Vu���U���@�����:N5 ��0" ���{�km���P�*��T��{W�}��]�|N<e3H��|�y�-�r��n
�?��Eϟ^���)K������:7o�ת�)�z��@��]=�U��?9���=P
���������uQ���Pa����+�3X��jjͲ'�&�F��U�j�8�M��-������װ����?�ģW��Ʒ\��5��v��wncj��,��cOL	��
����Xَ���ĺ�+b_|1�K�����T�mч���">J(�XR)G��$����&��Y�]љl�IcSD[�����Z{br4wkh{�k�?"S딡��}�����Z����T2�
9�R��RKّ^��ڕ��0��C'�^Qc6%I������ٞ��Ƥ꬏�`KL;b�������E$�!*����j���@P&��3x?S��?��y��J!��5��΄֙�C�w1+Y�� �Y���ԙ-it���q����?������䓌�w���x�f�R��Z�E��=���2�J�c�D��Hl�%��5��������g�5g�y��.�W�8���&�!�N���ƫ�D�w��]o&����h��\�[�8W.ġ�Bl,®�2���Xg,���p&A���\�v�˱��ӊ}���Ĵ�Vtf�����EW�]��*tE`\��B N�+�)�8�+���Z����ך"�����o����� ��;����bb���8�nM��M
c:�gΈItl�A���<0ӘXl�%g�&�wP���y��[��+y��[��\l��q�-B'y�EBe=����#�}�D
Gȷ'`%��2�hy���p`�ڧ=Jj��[����������⏗�0*ܣXH������&(B���;�9GϹ+�l7�����۶ǫ����F��ҍ�}�����A�@^���:A��5iO~���o�����6��%���r���M���i���-Z\��Y��O�q5i�3���h�G���Wv}�k�©z�q��2D���Q��6iŠY����e�iÓ�G�K�ת@a���P���b�i�C0H�S�O��x����VO�xyd뚸'��l3WӸW�$1�hԗ��V��ȫS%%�R|j�ƣfN)	�%'a���/پ����� ��T�-�D:����p�����R8d��Ys����7�,C���#w�X��lj��d��ffZ�5��%�S
��,u
�����O��+H���-��6\��O(�� �X�N���0%T䯮���j;`bI����z���q�]��6���t���d&�@�l+�zSZ�WRPg ;ö�+�(W�����o�����) T�9�G���ʚkՙD?N]��9���q2���H@͌�~f40�E�	"��m j:�$�*�c2u�(��V��i�u�+7b~�1������Hǲ�F�hiƊ6,j�cas�62bV���E:����ct����D#���=҄.������՘�v��8z���!T�3U��R��jG��NoJkC(�����DEDjm�L�<���*����=3�sl�Y��,�~�/F���edTg��TYѴ*O'����Bo��\%�����L��U=h_<�.	�0aD�G�҆���m�=U�����#�w��X���8ߟ9�w��췧����?��O'5)�w�gԔT'
UE��R/��7 O�⁤'������8�s��K�N`ؠ]Ӥ���럥��y��@������v���ĝ�x�Hͷ{���}����͌���]�8�J�>0�������iSh*��cY��A�������+2�=���@x&��8&�15���>�$�Gq�>�S�����;K/��rᴵ���l\���][���^�7�nR8�⼭��o,�8m���^����4�W+���0$��r�n���θд:�4��6�ų!2�u�ql�c[h낢Y�
��"y�7\s������7���N�`��ɴ(n��c0�A)$ToC@�,�
�cV���W�^��1�;]�(l�&�7E�h�ugc_8ۂ)�Nũh>��	(����+��%���`1.U���`�h-n�_i#��p�؊k�ٷ����7ڂC�m�84�%��J�pi*~7i�85݃M�n�^��b��0��E;�j��*���mr[1����58��ƣ�J<ʖcUg	fu����߁���q�M�l��HA��]��^m9Fd\{%��*iX���s��Y�^Uצe*�HWW O�1)\�q���[DX�v�ǀ����y Mv���]�tbʀ��5���8�&b�Ml4�I�xg�ܸI�;�]X�k�b�K*|�j��W�s�l�j`�Q��|,3�qLϥ�S6��/�'Z��DQ�[�o�[��V��ʸ�&�(=j��[�<O�M��������������m,`}S5%>�8=���~�z�$���C��ԭ$�c
{t��g*��`�P�F'�oO�;Ka���*2���d��~�:�Tk����������&�:S���s�R�k��u��4��N��QԦ�j%%�*��Y�ED:���kߍe;wj7���On\��&��IPz��gy�!��=���O�$��yQ�J��X^����h����q���ҝ��<�eUU�j2beb��]�Kv-��Tc�X�L  ��IDAT�E��$�œQ��Zu�f�`{���1��������[��?��͝��1�����ͣ��|����xHf�`e�u|�,n�F��-ro*H�KU�ƨ�]q��?� ��|�*'���)�.у��6~\����Q�΂p#�uP����\_�be���
�,�$׎�c����W�(a��~Y7�]s�����ueYs5�3H��C�@��<t�-�
�xz�&�����MIw1&�Ü"�� K�[�!�R�ʌAIfM7f\�kY1��U��j���>�����|�߇OG�pnV5�,���¬8~[���+rx������`w%�)���R��,���
� @俨ˍU9��$�_g���T�LO��Qq�Þ��lj��
/��0>ӊ	�t�q�I�.���k�ZԽ*�S=cM�ޕ�� �W��M��CtX8j�,�#��%e�TǪq������}k�@ǯ�x~��&4�ص�?p����t��ޢ���s\�����p�^��w�����.� �Q���K��Qm�]>���W^�rUÑ���{����f�SV;�Uv|�/_I?\���9|h�6eپݛ�i�>�d?��ܯ�`�f�PS��^�7��Ľ��y��6/�����㥪�y�Jj���RZW%��<y|G�W�ۯ?Ѫ�U�������;Q�;R��5�@�j����u�����~S�N_m}��|}�'��O��e�lZG���ڃ�v���򠧭;����MO��&6���VoK;��q�d����qn�w`�[ S<�����d'��z�I��#KN��_ٹr�х/_鬷/�zxp�ٙ��|����n�|m��)3>�R��s�э=n^L)�v񧧳/�}"94j&��̦]T:d�9f��;C\����N_[YK�m��g�,�n�zZ8��̞n��r���#-��h��J��꬘9��z��p!>"������a?�64�Ǥ�>ƍwa�j��vb�d���a�dVM������`�|7�`v6��@�M ̱�v�	h5ڍI��79�I��1kxD�I�O0mt
ӆ�cR�9�N���]�>t�����W$���Ww��=�.~�G��(�2Q�qt�����j2k���{��{0����bQg��0+X�� �Q�z	C��b'�b<�;�,K�kխ&%��6ȹ�.܄��?U[�1a%�������Fj*�� ��g\gFuWjU�a��)＄~�gѿ�h�u���%}:�c҈I4l���j	�[EW�6:
��Bj��j�۔�Q\j\���Uڶg^]��Y���إբ��0�~ZrjɿU��Ӈ���!�_��o��_a��WL��|_������n�ǹ�HM����>yί��r�ǟx,p�C��;`�E��U�/$v�.ܡ�{;In7��&=�k܆��}�<��CG�@��4U@�ޭ�ѻ���^މ�MJ2�뷏�ϖ���u�x��^*�30����"N~S�_o6���*�>m��뵸x��o����Y���Q�kS�<��ZD�4�/���L��7�K�0gx�������a[��p���<��>�^��/��e����iق�����;��ʕ��8��jߠ����ˬ��f^�%����rt��$��Bc��;�]1L񌠉$Գ��e�a��X�w�}�HJ�����f��Gȓ�$��dbX�$f�$�k�Zc�m�s���Lo��K��3H��M��+�L��`I��^Z[1s�Fs3M�f�t&�EOI�]�HU����a1�6���z�׫�媪RU�9C��a b_�GǦ�>z	�	����x(�T�d��P�}$qR���{�#��P�fl)0g!pf.2�=9�]�\g�iB"%��&�!��H��W)��Z��dA��%�>Tx�(؁�1F����5Q��ck����ұ��:�����&�s�X�������[_��Kx���Ǜ�x��OV��v�y�5/�7�ɎFp�3/?���=x�W�{��rkK#M������<;Й?v�ٞ��Ә���#�D�xW�:�F�Y��e|;��h��aZ=+��X2��=]l)�5"��D��z���3�ɳT�U~_թCU���z�&G�-@�!��C������F��c�=vu4-�õ��p[`��[ؾi�׮�ӃG���I~��,���ų?h:�ݷ|����}�O�|�ş�r�� ����|y��?��oN�������_s��Y.�;����q��ל:�9�e��=r�-lݰ�-�6�i�:�l����ظz%�6�e��u�޺���W��J6�^���[���K�j�"�7���F0z� f����ә7s2o͜Ȍ���;�]�͙��w��a�vl����ٵu'G��#'9q�SN���?��3_}�7_�N���Y�d9�v���O�q��q�����;�c�.v����{ٵ};��eǖ=��v�M�v�f�֬\Ǌ�W�h�R/Xƺ�+Y9ok�g��{����n�\��$P~�hI'T;\ծU��}�*�EYX+����I�:Y�o\�k�fQ��շ�`lK��������X�c�o4��X��Z)�UMM�*1�UI�l����8GF�(6��y5�P���r���ƨdf�/%C�ΕLy�b-�)�)�
�sa��,zk	a.�Rೠ����q%V�)EY:Hz#i�����D	��Y�Q�4�.R(���{P{;�5R������t�>��t�ÓI�ٚ�ʥj{1�8$���z&��^ˢ� 凴�f>¸���:f����X`ʲ� ֕R�wbZ!p%ۺ*������5�ms��]q�r�U ;�o\�`m��i�	��9�/�<��=Z��*UX�m@jʂV& X�M��I=�[���P;�y��	����-������l�ނ�i&�|�o�dRg�u6`^g���]��k��Fګ6y���՜����*��U���*]N�h�km;���n[7�I�#hݬ3�9y�`��gZ>�qI��ȡɰa������o�Gf]k5�?����r|k��Z����d��$&�ƃF��O��H�B0NI��z�5^�ݯ O��y�?�?/*x�T�.�F����y��K7x����s���zK��Ժj����W�w��ot��>)-�R�I�Aǩ���-�C�^)�1�F|���v�.d��In�^�VVP�I	='�d�Gk��ܗ<�B���RxEb��;x,�OO��˵R���˃�9ܺ�ē���`�	�4�ųܺ=�C�:�lsO���O���x!??~�UȪ@7�����!�o-*�o�8/�a[/��L��%��Av:���h:����C�|k0��v��Fd6�G|��8��`�El�ɉ���o[)پ�f�`m����40w��$�ˇOa~�^4�pg�$zch�K��G4�āA�Nt�r���YRzU��EYYi���M�A�R���`Ū1��nKM�#�J�#--����Af&���()���@O2�p#3"M$c`2H��SC��v{j��`+K.Ժa~�Z�f옉$�&kU�a�ڠƪ�Y��:+�m��0c���5�Ӄ��l(�3HU��A�ԩ�����ʒ�f�5ӑjgN��5�!�t�t���g�%ò����rk7�c[/���95��n.)����Y�����y��Xӓ-�<�P�{k˸��>�g�Ÿx>�>і�Al����ެh���fN�o�̻ܘS���2W�[3�؄�u�x��3�{2�ʕU�,mbê�l��ɾ�!���·o��ƪ
�������_[8ؔ������u846�ڸ3�Ԗ��6tO���ϒXS�f}6��@W����+�dmG��AaK!@e���?\~c���Pm5U�@se���N\<�O�ƼI�շ�`��q�=v&c�f��ь:�aF
D�ḛ�Tc?bÇ��~���C�ޢn=�ա��uaX���2�>}�[�Ԗ�}{3�wt�E����յ;=:u�g�v�hߚ��[ѱm:�mJ���ܣ3c�aD���Ws'�ԱØ2~������0q�0��N��޿#e}x����ݑn=��@o���ð���$#����3�O?�:`�f��a�1�a��Ч��cOڷlK�&-hѬ%M�4�Q���5������а�9ʛPUޜƕmiҠ��M�(mI��VTʱ%������2o�<�O��{&�}�_��4N�-߶���|�:YZ����M�uO)�y�|��4��8��jsi���|��NZ{L/k)��a�F���֓Z�?��d���.��;K�a�l~4���N��~c9?`���7���u���4|,�O��!���� .σ�s�9n�K+ic��=�:1Ļx�{f��Q���;L�1/� m(�`wo�<�qu���/��A��o�D��]��yAv�	(H:���[����iC�ؙXIڒ����{8�5
��Z�����-@��8�A�i� ]�A���y��
�*�`\%P��]���gcY%Ǖ@L�Q�P�A���u�:��i�@�@�r���DV���=��O��q� ^�MXU�Ʋl'��vbS������=kr~�_?�e~ݝ���Ģd���x�U�U�<�b=��٢�By���>�����x�7ȫ�Ay�rn����Q��*z�A�(.jN���hߦ/5��p
OЬx֑��V��Mt
՛��ǌit�2�xy������R�@<��ܳ�q�Y���w��7�rGu��P�g��uɠ���=�V;�_�?/��<�t�V�w��-)��ʯ?����?^YUX���bxʢ�Y_>դ���|��5�OѠ�X�ȷ�Q��6c�Q�w8%ͩ�s�6,�jwXٿ��^�n��u�CV�v$V5$�S+�͚ȶ�;y��V��`Rߔt�NT��75�t���.����R�������<z�P�T2����&�v�_�؇��r��ͨ�vjQ=Q��I��G��z�'5���T����i�!��gz����\����`3���`Zw˦M����Z��I.��!�]�?�^���;1�ǏI����uq���M@̗q�F3�;��J$J>�����K�[�ȉl�-�:3)m[�a�8��J��UM2dza���e�٩e-`g���ة�B$��6!��D��oi�I�G�I�Y'0&�$�Q
`���"Z�ySQrN��&��AјP�� 9_U��iё�cf�*��)�PC��AƄ������9
U�������5�EI��$��������^Y�U5l��N�dz[��ߌN��K3g\m[f��2��%��qh�'�&rO@���*�k���Mx����n�/���[���ϱ�����Ǝ�,�
�ݒP��2!Ջ�鞌��ch�9"M�fB�`#z���壣��H�5W��_G_��c`�(T� ��pCd{D��!:���0��D&'��v�+��}��#�O&�p��r����Ϗ:���V<�Y��)����-,��mD�H3�=a���
����Tj��\�?��Cf` �V����Q�N��7�M��*@Xk��TVK�IV6�++�ط/�GNbD�!�ϫKz\*I�Ո��Z|
�	Y��d��F�W8�n�����O��/���$�{��ObL �񁤥�Q��J��\�ɦi�Z4)�I���hY���J�ݾ��*ܫ3F���I]Y��0V�ͦ�3����|�e%Gv����|zb�N�����[طg5;��ώ-�ؾa;6-d��9,}���wF0w�H�3��s���;cy��L�:�)��k�0��\zгWSZ�*�ae��Zm�呛S�������F\T�f�N��DBB��T-��LR�e��RC�EjR��B�<�&�0�� �$���v�iy��y�œiᢵ�TV:5�y�@\�@[�����X�k�k�F�����ڠ�j��8+Դ�j]͡�hbGu+wҭ]���	:����إܞ�>�u�7e=�X�?W��F���j6�_J:q�^'���N��شߕt�b��<�7G�dGQ#ZI�*�
w� �֓jV�d�F1��N}���H��X�Չg{��\ĵ��z�'�{�݇ps$�˶u'��YS��#q�G�6���AL6���QQ���+�wh�O�<�EK Ψ�1���
\U�T`δJ��� ���k�<寬~���,gfU�O N�� ����;�*�3��i���3�w3����;]��Z��޵hxLG�AB<�|}8�����Ҧ�v�+vb_���M8
���݁k�.�d]U���ۢ��3R#T5n�̋�m׬~&~Jzȓ��	�T;����q�?���`�����>}���^�|���y ��-��IC��EH<N���	�'�PұmF�'�~��aѷv]mȔ��UU�S��|�jc.iH�������/�L@��ο�t�N�yy�f�{����x�"_��^��i��Z��z��W۪�[U�C'	������۰��#��c�lZ��H���
��J{ _
u�]�P�Ww�{��N���v�Kf��ķhAM)���5�_�^�[%�ז�c_��չ:\�+ w�	�����ܼ�X ���u受y��������@��i\�vJ끪����ބ��',���x�'���@�H{��,Xޒ{�gr�Nw-������te"�h���s��.=�Όy�Hȓ��X2�0W�<=i��NS'��$�rq��ܕ���7m-�ӬV�*R�3��K�{ђP��aj�%�jnR5���~ժZ�R�.R��S�
�EAV&R:6��(k3MsA�mc��E�>�fM�[�����'@�ϊ�����5�)�W���%���_�����yj�7�s7�ށ Ke	4����Zu���&๊��d����R��=iu��,�:K�^St��:ڌ�����i�{]Y�5��2�0���V��hK�V��˂~�[����8<(��m�X�ЍY��K� ��f���&���AoA���b@�c��i͸X[���03˃�5<y7ǋ�y�|PύՕnlj�϶�!���}8�ŉ��vњ��M;�E��I �����؇5e�,���{�&3 F�P�6*W��::�w����H������� �#�y��-�R��.�+�PD�f�Pm���	 9$U-�߯�h�v���y��p5�}Td�E��Τ��S��AU�|��ԥ^~1�Q�D�GdH����GV#>0�H�X�j.�͋�@}�L��`jEz��F���4+�{��v�d|�LҎ��3nPKޙ؍�s��c�v��ĮSػy
[Wgǚ1?0�������'xt㜤v���~���H��z�jS�]=Ï?����_r��i~�x�ӧwr��j�XĞ]sr��JN}��/���'�����Kطo���d��1�_4��c�ҪE>��3()̦�N.�j�R=;��Yd�����DzZ�ɤ�&���LRR���$'&�����"��DfF
5��Ȯ. ��DZl"�1���I!"�����E0"4���ǄF36,�	a�Zӎ)r��FD3Q~�Qa����`xp�(�q�������i�D�w�.��4�H>�i���r6��e]B���::��q�ٗR�\v��dr��!���9�؜QΖ�|��gkR>�=�H��v��t���+�S�6�=��X@��Lz��iqN�`)�Ƚ���7��>A��c����2�-�ގ^�u����/����K#'w�ƥ�b�T���Iǲft�Ә��V���R.�@	�5:�yc�F^��k(��HI ��a,�,�L��)+\��R���5:����1eu�,߃� �U���}$����� OY�`]�clJ�ze�1)߫Y��nǧY��:�Dj�'�(ߥu�p�y��YX���&yv��qJ��S����[�Y�J,�6b^�V媪l-lU��������i�W���Tյ)���'��mDWg%FyK��Ĵ�B�jO�u�yt�֛zy�tiݕ^�FP����8�c�qK��*"E�mT���}Io�N ��:%���ڳ�vx��x��Q��,�3�xo�n�`M�3��İ<�7���5�6�������t��Ξ=ϯ�\}u���u[�!�O��:e���?�?��OP����ۯ�Y�����|�@�@^�#i4t���׾٭[Sй+���#��@
��"[`/�mgmX;�?`��S<y5���{T��}�E%~m­�y�-Wo6���ܺמ{{���py�c����~k��w�r��D��\+�s���l�?{"�sWO��<���C8�W�����}��������3n߻̦�3����}�v�3�����#�ٹ����Zn��/7����HJ[fa���S)�z8�ekI��1a����m̉�f�Թ��7�� �:;�gmJ�����-f�ZOV}�ѢX���f�oCg��o�<��z�*�R���i��7�a���)e)3T��ɶ�ߛ2t�0l�X�iǩ�[*<�*O�>u-5�{OyY'M�E��d������\�\�����pa&��uؘ�js,Z�����6n��W�R�&9XR�L�t'��X�v�[�qxx,�/����\�Дs��99���}�x�*�YyA��pbP�}��Bu���O�!Q:�%똢z���1�@Ǽc�UZ���3�;��g�;z���'���A����1Q|7%��N��..����Y\����g�ۚ<n�)���|nm,��z��u�\Y���5����6?.�ͅ����\�ͨ�g�9�/�]]�Y�ȕyu�x;Ǌ�)�LL�gfmv���ܼ*.�j"�׈곢]8�j:Q�/N��M'�f!�FB�Tlm1�gjel!�U\�1f�\�޵f�^�j[���7[���z�zy��G��_� a�aKF�D��H�dđn�Ts� ��j�6�z��bOU����P��A���]�?�%�����UX��h�.���S���2.����v��۸pn3����_��3;�r�3��t��X�r��7�f�Tj�$��T���=n޸*��bEt�;~���~�>��_�s��'\��ׯ~ʃ�_˹?��ᗚ�]=�W�l`ǮYL�љ��Kh٬6�Q+�:qI����Ed@0���E�@Hh �[^������g�AA~y���'��=�}I�����5����j�	��PpDp�?�C~���X�^��G�yH5>L���8��M�ۘ$�ŧ���'5�)2y���֎��N�qp� ��H>ʩŮn]�ޤ�����kD0��C�M���$��3'�%Crl�$�ԩ���NFd�G(��彪��aBv	�L]���P �HD_z��w
'��8����Nd��o2'C�8���F��3�]�^�l�	e�_�"�Y `pl�[��q ��cF��t��I`�L�vb�@���ZG	��`,�g��SM�?�R�q)�-`��="�w�������ױ|��6�]w5>�kp�_�kݽx4>�����Z��6er^�j,k|�Y���4jP��v"�͞fI�Ԭ��]��W�N�c�0 ��F8���1��>�q��s`]t�0��y���f�*wj�j�Y=v�{%�]�VtE��ֿ��u��?��v'է	�e���;�ل�L�܅�d�����.ì�\B�fR�z�+�Тn9���m���F�c)�]d�i��gj�Z$��D\Ӷ�9��L[��+	+�"��RB�3�n�^:f�\�փG�ͯW��a���K�� �������_�0M�������hC��q��._���'����BW|���z��C�)������_��3Lyo>-����P�����@M���)�ы�](�1�����c�]�С;q��iշӖ���s�F���x���������y_t�����y҉�O�r�I�������?�����v�]��m���O���v�O�<��w���ӷ�Su�
���|Ě0i��܋�7&��`�N�ž�����SE��>-	h�Z�F������'�ݜ���&�ņj��;K&������cY1�=FU�3�n�+J�P�cj2%��q��'%�&��4�����#m�\�4�����+�Q���2��D�/XXQ�ܒk[j��gkK-+M9���Z[hn��%�V��RK���I)߈T��SDi"�mb�5��(�njA����gCM�V��	r\gF����S���B����*�d�
S��ܤ�2�s�%cPC���b#�v��#A:k�WS6�lt��:�&ɕ���j�ú�����e�[ی3s�88>���x�̑1i��E�1&љ��nL�udV�#�����?�Z��C(zF�� �0G��@۷�9�N5ο��O��eq�Ves��t�-M����ؐ��9<ݖ˟{���P%|� �T�qY���h'[�Z�z38%��9|�J'E�[���My�QS^|ؘ'�rwc�k���e��Q����s�O6�&�V�cR��i̴bKv��ws�95�P�=�޵|�l���)�FXZ��HbR��t�����D�j�zᚙ��E��O�٩6]�^�{���fp���OW�==�����ח _?�<\��t2�f��юD�
�[�H�2aV�lɘk�<'��)��^��a��Z��u�1�5�F���I]ز|_|�����ʍK��҇{����}�p���|��"���'Z��#��L>o�I�+i߶�/^�ԬW�]���K\��{.�;�����wq��#�r�$��r���r��ܹ�57n|��[�r�=?�>�����u�ټn6[7.`Ҹa�!82���8|\<�wv��	�
�K�7<�9989���򆜴g�������� ������RId�W�̃9f�	{?N�y���;�X����U�)sW>7s�+k>7q�K#G�1s⌹3�~��dL�V�Za�_ O}��l�ɗAa�ϔ���c�~�?~�1�v����8�a1_�^ͷ7��޵��t?_�p����3*��|���4K�$MRU��R@k��͜���?��G���>wI��H�5�e$�-#4}e���|i ���1[O��zp�Γ���|���AGo��x��+�5���Ÿ�x�EOF���nt�ї��w1���k0g�Xy��}�I��1kz
��i�[��z��٘�Ǫ��f}SÚ8Vl±p�Y�0��qpg�B{��8��w�E�:]�z���s����E��(yV�+1���7��ޛ�'� o?vea�]���K`M��s��?��<��˰˙�e��-ZتzY��5��:��}��7��Y���C^�6���j�;���Q����vx���0��e��<k6�u�Q�x0�yh]�P���▸�E��u�'n�!DT'�Q}B��j`\ْ�f��/�Џ�Q����8g`�T��"j���᯾լT��iql�q��^}��aQG�'��E�#��BL�}���|�{w�ON���A-�R�i�%�Ke����j�'�Uo����t�AI�����S܁t�:���}�nߕ���(�7��N�H�؋j{�ۃ��9������Հк#�����\�߂�6��Ӗ��ޔ�/;��e/�$�d�=����vm%���H����L���Г�a�O7�?]�p������?����zjBߢ?�z�u��q��-���(���T+�EVE:�?�ã�V�q{?r��H�S�����a.	���{'
�#(s��������Q�ɝXWzIIh����ں;��嫒�|Q��JZ�sE'�/l�'I�쒒��X��&q�?����2(���1�����ŰKJ�ۂ���V�6�)(������W~j;Fs�����;�<�X���bg_����+��>᚟�:fSp�Y�%ǻ�h�$k[vaÐ1�IHg�[0s%�����X�Ԧ��3��]s'��D&�����X� G;81�ց~v��t����+e�1�:��(ؒ�&L�g��}961��7���˒����'�uN�1>Ø���,,0cU}sv�q���|:<����fj
?ͫͯKK����+k*�ms�w���`�W���&�f�y�5H��k�_
�l���2��-��*8$�|(:$�>j(���;�Q�;���������=�z�
 o+ (�|&����wC��`��}փ���s�`nl*��\����ǽ�Y�Е�j�0*U�9Ɉ���Y�>���t�𦆏�Ve�z�&�ŒS-?~e�U����uD�Y��)���%�e�US��
����fo�z�u'�';���b<V�=��rr���F ϔ�gjG�d���HG5o�v���N���R'Ď��6���ʥo����M�&E�kQ´~�Y:��O�����x�v�~��krp�j>�xW���Gw�oX�L� ��'I��uU@���!�\�ķ_��c��p�6������Y��l�/�˂wf�f��·�$���G�9vl{w-a�w�x�
�}}�S�>d����׮KhT2�1�{�!�A�_(a>�򼬱���E
?6�.��{���U䌓��&g7W\�<���:+���g`$�<"�+�v�ґ��v�h�m��g�;󡩛���L<8f鯹�����ԕ�{�l|8�á��Է�#R@��ƅD�}Y�r->�ϼb����#8s��e'T�K5L����?��磇ܽ���'N�oԉ�6|��w��4u&�̆k')$��X�sNn	�����Y�O��.� ��\9�sf��+;t��u��:����A�k��k$��\�
�*���f�lt	eEF���Ÿ�N��o��t���T[;y�FQJ��b��$M�b[����1k�ED[̳���h���~�\d�{b�F����ĳ�y8a����ؕ��������&N��й����$�;NE�w����Y�ހ<%�_qP��UC�XfM�9}nIm����#���ftí��K`Swfep����E�z�V�������
�lX�"0*��䙪����n���hc� �fFu�3&��%�k-���lt��`�9������$'��f��ܬur���zQ8yŎ4h�C���iܳ6Ie��P����7Pl�)(�
��B,��d���[�k�����O4�!J^H�M����9A���I+�T�j\�����G~8��j�5>�/�h0(�[����ý'wy$ߐ�B��o�`���t7�c�S�g(9�hé�w�Cf�n�[�g �;u#�MR�u$�[o��u�v��l>pDa��C�;�m?^o̕{��r���O�p�YSn>ḷ�]4���=y�G��^<z2��,��<\Tᨈ��������ly�p^�ky}}��*�S��=����V6$�nC���S�˞/Gr��Ey#(�_��ↄ�n�w���c�-%t';Z
hut`��fDB"��}I5��qb�MdO��,��{('C8��q����s�܅}:{N�y�Y �u^����$������1I��X�𑅣�� ��d��v��kõ|h���vq�⠍����|�ڝ�Vn����.�S�c��!)����Z?$�nu�Ƕ^��fI`��ek����Le�G8{�}Y�������qt���ɍ�.�/�K=X,�h�����gm���xG/=;:�Y�'Iy�m*�۰8�y�._N)em�Hf�vbh�1�R�x�ؕ�>l��ѡ595*C����T�]�ϓ-����.h��������@�PY�'�l�� ;�>m'��Aܮ�v�ɡ<�ӊ�ۚ�b[k�nlƽ5�mu7�Tq}�������-*�Ҽ��+�Ҝz\�Q�O�J���R.�[¥w
��72�o�C	�ޞ.<=,�����k�y�/��r%~g:����<�)���&\^Pʩ�٬n��Z���12Ӟ)E���i��lՠ�&���R�Z2�hq���[[i�4���H��"M�,��Bk�ok���VCߨ�NNڄ��sqr�U����]<z���8;8��S�r�� ғ��Z�ywk��3�mk�gShI��C��Yݳ(bv�"��*dT�&��׎e�����X0���b��w9�q	7��}�9yd'�~<ã�7�K��@�G-	����O�j3�ۭ����+�|.�vt[7/f��i�]4�Y�&2v�PF����9m4�/���ٻ[
u�w����,]8�6-ې�R���L�Ȓw>=$���0� cad���-�N�� �W������	{��eO����?n�T����W ��C�i$߮�5�L-�f�$����؞�Al�a�k;�q�\A������] ��T��k4�gP��B��0�ދ$�9�	4>�-�\x.�}�H�μ�k8��|����p�g~��7o���իܾ}��/�ʄ��iP��ޑ|!�vJ2}5�^�Q5�v� TmìE�:{�L{���I�v�t�CU�n�4sd�ܓ�3�7k/6Zx���C�Ν�	�*���a�����<)�Mf���Wo̔��t��_�ۯ!OY�4�� �^c�`7��1�큭oml����>�ƛ�ht�K1��}Xs��J<�*�Li�_z3��0v��(�=���h�J�kV�1�)Gg��%����/}y�bg���o �r�yj���Mx�.�C`�$�����ml3��'��x.�뱬�U�Q��"����=��<�R��+��:�1z�O�<�.��Z�n�e�!O
|��3�O%�䘚�jpg�������.����kQUP�z��-��}�HV��e߁bN~ՍM;2���tYA^��+k[�Elqa���^@`�z8�e�դ#�>ӌIj
���=փ����'xJ
C�眠A�?�?-�B���������ݸ~_�s�3������S�"+����5��x��謹$�R�=8��9F�����g�x�Tr:t#�]W�:�&�Mgr:����@r�� �m;�[��F�����M�d�&<�6��@������dx������r~Ғ��j����s?���v�=�����W����rn?|����1�"�Fv�"�����n_������Ɉ���^4W��S��� �N�EA��ڏ�S�����YU*��{|��xJ[��_P�wa|�jc�����6
`������N[Wj�,�����c8ԡ�y��R@�TrI�U·��Y���R��PJ�JIW+�Ji�M��J�����FV��YJ�؂��Ͳ�Qg�iÿȖ-�.l��s�*=;�Z t��5kL�Xkf�&+�[I)Z�k�dM5m�8*�3�e�\c���WX��W��go���f����e�
#�Zy�\�u��K%���s$�o�0[�Ċ��9�ma�x�����FG�w�\��1��3�pdT>�[�`Z�p�E�1%ӝ�U�l����a�|=)���r}e�����N ��gk���Y��zЉ΍��'�W7��{�t�]-x��w�n�h����\ZP��9圝Y�o&����|�����5��%�M�RY׺��$��U��/�U��X\β�hQ����bYZʲ��j��V�lh��N���'�j����ϩ����]@�C�d[�\��� ���}�yyv8������m�~q]�If^�#S,�:�T�y��AΤ��niGN@i���ZX�cdL��)�"��y'��`bJ�+7R��^���]@���w��p��w�:����ܽq��'@�2'ԕ�q����-y)ά�_��ZF��aD���3<��2M��3�ezVe0�k=�ڎ�S{�g�0���'[pt�N~��]���ȇ����8�c�_���/���]����Q��90�'Z�+����郻ܸr�+�|ͧ�vpp�vl[��ų?�F�c̈�L�П�g���7nx�=;װo�2>ڽ���>`���Ԫ���Y�F^�LꦤkC�T��O�W.mee���3�vnX�8km"��u���Q��@����g��\� F�$��E Ng�z��6��f+'��Z	�Yr�ő%)\�:���Vp�#�#V��й�ΉS�~e��Yk.�q6:�.��ZG�@W�u�,���Oq霍��[?
#�hܦ%�oa��m,|{�>X˱�������W�8t����&/$�y!	�N��@T�=C�0�#��C�6��(�֨��u)�M]�{�j��9X�0�4d���aRx�i��v'� �M�#-M2sc���,�X-��\�WJ�Ng�r[oU/��[Ԏ��MX�b-jtī�,�Ū�ItU'�佲�UŲ�'ڔg����
p�M��/��8��j�]�E���\} �y#�;�����+�Fn5х��N`�{�&��֯;�4�S�Y�a��������![*?�{u��D�C��YՇ8Vn�+�-���a�'��׊��6�&���ϴ��S��O�W��eZ���sj��L�b���X�DWc����'���d��fz�R��{��\�.e�)���c�8���x���[-���4���_��9.�]�8�s-n?n�czq�q��О�Kxki&}&�Q�A
�����'�&�	�L\��[��j-ߔ�� �)��hc���ԺAo�����_I���ff�"���i�_R���o�o˺��!˛�cXۯ$+NRղ����%}����n�~	�/U�'��>b��G�8�-jwJa�Az�몪j{Q�k8�{�"�WR;t"�E{�:��r��L�ķ�p��$��x��9���˹x�9W�6���Jy����������<y6�;Ozs��p��ô�Y�z1�>=]��<�������M�ghӣ�����O�2n���nӚ�6������O�����\�e�[��Hj�FD���1$ +?w���!�[�V���d���$��t�K3��c�>�
f��;L����$�S�i��� � D@���k��#���[@Ii�@��N��k�zw[���(���n��^�%l�l4���v�$��jd�@�*�[)��J l���ȑ��R�v�}I�׈֚�i��
c�\o�Έ���
aK���7�1�5�/��J�U��5S�码�{H8s�|y�	��0�`��-��jgA�0Sʜ�qjl�ڇ3��+�Sܘ���z������d�<�T�_���gpߍ����T�0I�G����8ޅ{{�h�3~�ܞk+[s��*��T��s�2��W"�;ǰ�]�[D����~s�0�V �3��,�2F�12ɕ�	N���w��6��ꑫ��G'���5a@���cW��:%�Bk382��	�vLH�g����b�����W�Ǧqv^~z����;�ǉ���t��Q���)��ǺruU9_N���6�L��J�H��S�gI��#�����ٓ,��klF�d��&:����cdNm#K�%�O62%U�%��(J�S��,w����y{{j����U�::�����cok���	�N%�b����Pgs������p�t���LteLI4o��aDU
]J�ѿy>�Z1�]!�n��1-Y<�7sG��q�Y4s ߟ���3Y�x+Mf��Ŝ8��sg���s���%��z�뗮q��+\����WN=�჻طs-���`ˆ�l\;������c�r��kH�V�hӢ.��VУkk����A}�;cKߝ��	�hڢ)�յaPjVK#?9�Ҍ4rb#��p�����@��+��-yгut���	gWr]X��z�Sp��mP[̭�'������CYӼ�+�:0����|����a|n�1{/>��lH�6�Y��-5\}��&C�����4������d��3j�N}�5�������g�i�޵�q��%�XA���$:��[8�jks���$U
n��ZG�
{g5���8;e1�$�� �SS)����rO���4�S5
���m6��z����,{�9�t�cY�
NN_z]�ߒ��Fӳ�?^y�4K�E��(�	�h�jQ��������)
k�$L�{cUg6U;1.]�Y��8�}������m�4�cR��o��Z�Q} �Q�1���ohm��q�LGg��]TK �ոw�ހ<w�
y�w�6,K���l���J�m�t-�?�vW`����_���Uc�)�q��A��Tg50�6w�ȸx���B�w�Q�|ts��-'8q ����J O@�vJ2A1=�e��.i���0��M�p�nD���LAl�S���S��=xgj ������,n?,���J���������hÍ����J�o,���Z�H��K��8���忯�˰�uU@3p�1��M*�V����W���?�<u��G�5�{p_��_4�Ӧ,��@��/��W�Ssت1�>y�﷮s��U�>TS$*�����Vﻟ~d���T�Oq��Z��:=��w!�� r��f�>du�A^\����ڞ��1v�XN~v��O��}|�	?\�ĕ�;�u� ���<z܋��{s�� �^ɑ�g0e�8�w���y�L O�m�YM#�=������� O�K��V�7�~k��lڂ��-�.m�[r"���p��*n>�@��1�&�h�KJ4���
����3g�H�7�ʆ��������s$C��l@����3�EI�,�a�d��"�@o���^���{
���n�@�nc;v�j�.Ц�U��Kx[%�-FJ� O2�u�z��7Ao�$�k��4����&z�[-��R`k�� �}��*��v�j�T��J2y�_Aގ�%�����@��$��H/(],��	�=y&
��ib�Hy�͌iaiL'+���b�t�gU�&�0.ۊy��)���q�2?�k�x���� ��_�������Hnm�������ggsbd6���s�{�D��nKJB�U;�I�A���˨4O�%83$ΑA1v􋰥G���n!V�:��1Ą��&t1�_�	C�M*~JC��1�ҘhK�G�3$̔Ar��P3YW���u����XKF%�3!ˍ�A,lϲ�q��^��Srym_~8��=?Y v0|ܒ���rvN:�{$�N�?��Y�F�������Q������=�!�K�<�LI�s�j
إKA#U 0���ȳ}y
�||�4)�SV<寪pmmm��x����ڄxrcI���فo7�����E��9y���Ȋ�Q�;m�9�&ٙ������~T%��8Ň�W�����GyB$����^R����۱3��dŴ�lY���+7�k�vl��G���ڶ��[�q`�N6�Z��X��-�_<��g��,v��v�U�2�5�K��B��J%+=�����L&-%���j�&��%PW��թ��B�j	T��">"���h|qq�gan���56��l���\��v���){y"[=K�.n�36(�5䭗���<Ͳ.�!e�?�̺�tf��0?��U��.�����Jf�G£�\��weM�4�I����p �)R��)=�}�t��aX׶:�9$-T��?���$���I�jҁ�ܦ��wH	Jf�}���8Q��:)HHZf�D��M�=� �7�,�z�ΈI������O O�+$m\l��R�N�˄�6ʬbE�A�(�O환T�9_�iS���P)�*��y��#�@�.u��1�fNq������U�Zm�E�>Lʶ`W��:K0N��_}�\31uK�>����xŷ��=+�4��JI�n��w&v	8�W�Sg,6�+�U�~w
6_�ݿ�<�sF��:�l���O� l�E�L_��U�V(W_����y�zܖm�C����`9�`�3��w��^�X�Gdn$����6y����B�0]���������z�S�+���I�'3"����DѲ�;�-���3yܼ����ly�GQ��Ւ5����C�Q��7�9t��O?.y�/���˥,a�z���3@޿���uʿ`���?���7���1佲�)W��}��.����у;��fr��g���尩t��Rث�:�ױ5��"�c7jv�FB˖�4jH���2i,#�Ob�]<y" *����?^�����n�����@^gm��+���_F�z� ���@�^�iѽ�?:���j8�#9�~����C���)�S�K�b.ڰ����DUVԐ��B2�����1���oǤi�8؆�kz�d���_�`��J&����������0[ �WgJ���l4�EٵxO2�UR�]kd���	��!�V ϖ�A;Eۤ4��U I�`�S`� �����<����@m�d$+W��@���U����Y��0q�;6+9�J\Mj]Y�VJ���V���۳��xF�e󎃳 �$�F�ߍ�y��zsNߕs��,y��lliN;#�x3�$���_`�"o�D�4���'��ss��6���k�d[m8$	ȇm��h7�<֟[�;���
������u��5�M-bY� ��u<����[���tbL���:�F�30҂�1�1�8km��!Q挈�bt��\���ƴ�����`J��
��Q��n|P����@�6�g}#H?65�fS3O64�E�I��(P��2oV����ԏyuܙ_�Ż��ʜ<) dJF����jN��6ez�3�E��k6�����6<��mZ��y��ח��qy,k��L�Q�oO��=Y�֚�.K~�tq3���.����T�;yoZ�����Q�)�S��OU�:
ZY[`fi���%�6���&D�y&����'0/a�
t�YF$U1dz�R?̈!�H	"�يZ�v��[�^�1���yѲF*o�nǌnֽ͘���G�r��.�>ƕ�����}��~��xq�1���?��!O������<�����č��p��A��^���X�`�,e���1�),�7��gM�z���݋��[k���FEJTl1q����;��l=�]�w����+++,-_A���6N���gc�A���)���A��^�m3�`�����a��r;?��iɕ	���b�����'pv���`S�F|=h0�N�����sy�V,|�f�e��jh����|_��Cq�L��������>�>���xt�)�/��o���wyq]� )�{�{�d�{5�g6�d\m���]MҊPk�7}''����6z1�'������������zI'>p�dan	Gƽ��¶N-gY�^t+��Lm�5��E����'RC��q�t�k�D8���%s0�iX���<}Nvh`��CQǨ����"��Q��s���q/$$�9����l#��H�7�߈:�\�YEb�[�����_�q�����i���Ų�~
�E�ˠz���\�IS9F<����z�� ��v������彏q�"t�3�N~��%�7��6�NLѷ�ݍO#"���z�1��IR�b��ۚ�zDF�J^^
��Һ�K�'�ٙZ���j�ݧ��;������y�>w�֕\��?�J���u ��P��Q$��w'3��L��!D�#b$H @p���������eY֗]v������a �w���}�s��v8tOKu�U��T�s&�H�-�����x��g�=�u��G�쿈ib��yL���/w���sbvS���&�eM�L��'��47��S<��.~��3���#W�E��K��i �[uCl�ֈk�
�ݬ�����e�n�aM��t� t Y�fo�&���\|s����Σ<��,O��������v?���]�wBja.J:dbƪA���st[����T�̙_5ooj�Y�X���n�y���=,3����k*����\_S�ݓi$^e���|Ǜso�!��L��YR#8&��;%yR��d<z�O^7�����@�,���Nj_t���~Z}�F4��B��'����Xڵ?U�嘮��J��Eb��j���$"^v2�#8�j)"���ED&��
z3A"��TIo$�\o!$���dU쟄���]�L�x��B�J�X/��c��-��b��ԝ[S��/�5y��v����_@4�*�XDy�C��Yc&A<��3C�]K�dݴ�E(�p�+���u��k�'Z�o-K��7`� \��{k���t�ܒ��JP�������8�e*v���չ�X�ꅙ�����eL�
B�1!T�сb�`l�I�����4����VX�!Ć6�l/Ucs�W:�x{g���s=�q�K\�낫�\qm�����D�������(��6/���m������%
?Ψ��fD��)�qml ��ƙ8՛��'��sÞ��X����$���	WcH��j�1��y�P�h����7������x�67�^��t��x��R��ˀz	�,y�c�M�x��j��_�k�y������Ύp�7i��r^��T�H��*$�)	�2v�<U+�
�F(��6Ju�g�B~�#b<�Vp(�cA�4tM�Fm�|_)�n�M�K1�W:�h����ۓ��ӕ����z�|s'n�t���_���/_>��V���M�������)}��h��xO~ͧ��%���9|��J�"���$�ـ�k���7v�0�i��	i������3?&Q&��.RXA �H���ALºj�(�q�h��A����A����׻�<fy�[��6j,�W�`e�4|�r��]�sŕ���K��۰m�Fl��7����f�X?_5n�뛶b�����
�g�R*����58|9��5��S��y��Ş�s���h�h6�[��a�qs�I�oTV^��٭q$ 	S��I��I�|Y&��%@M(�ݡsx��C�qN�C�N*SjB��od�O��1�۬p�z�=��x��V*,�2uf�����	��-8�*�>�.)&��!p:�k�>C3�8���Seo�:fv�8�@�0����87�咥��4}=��AUo,�tl�w���K�\�A�	�T�1B] 4z?HU>���M��\ +J�#`�J�V����3��!�����fV-<K��H�GbWX�/�0����wIx��(���I2�'h��)+�nY��B��CV�!������D��b���y�<��M�/㭄E>���j�1����N����� �eF ��݆8b�����[�7���ɳJ���7�h���I�W]����(}���o��z,^=ێ��L��3���V��62���|ڱ��+����f���~��;����bڝ��榉-�@�S���M5��p����xx�.޽1E�`��t�1�l?��C�#��p�7�Ze�Q�1�ݑX9�~wG@iGx��wq3�jZ��v�0b�l<xB�Fy�N\J��[�����~@��<�����E�;�g"�iC�螃��+���9x��"=�?x�a��?yO�<�����f1�>j�jʿw����&�3n<pn�ɼ7n��T���/-��(��u������X�3)�ސ��B�'�;:�l1V�D�/֨��.��x$h�s�Ōv����l['� �[/�"ȳ ȳ�n���T�2�N��d�ۦ��?�	�,M�g)$�c��#���c���b�V����w<�Q��A�R��7�ؘW�-b�4�׀�yb�<K%xfa�7��o�@��R1
4:�k1�U �v��wⰬ�.�O�ݵx�-���m����"\��m<���R���Q�\ǈ)u�iN�.��1���8�+s�<�[��cWO�ꇓ��pv�7����j��)upwv~��s��xQ��NËu�x�9U�)�syK]d��
��́��V��6�5,��$)�ߴ�
��f��]���QE3�;U�'�����}E��E�ߕT��K�����nd]����mB�<���:F֑aXm+��az����Ǚ�x�����U[r�ìX��ZcR�Q�@��qZ"���!�,�!���¤ͣ���-,�R× �A<6���<��c�<���Ff�J�C�\��E,%��Ʀ�E
H�RW��Hre����q���`D�:T�4W�b�&�[د!�vO��.yީ�O�#���ܡY�va5�_݆_�7?^�Ϸ�ǣg���wlj��Q�e*���_�o�SK���x��&��~�.��]��ڱK�M��53�e�Bl۾3�ü�c1�$8 �y�'�y;9��Q�'
��
�2�\��$4����3�3j����b��]`�A��*{̳��W�����\�yW+���`�7�T��8���;p���
��8���Q��3i&vlގH_�e2Az;�{b��K�N8ע6�2�cE|#,O��Z�X��%��R��p�����|ӸֆĢX(E]KO�;m�$��m�º�L�9�O���(��y�w� o�X�"��� �i�vR9�C´�6ئv�&���yM�*j/"�����#f`"A^��t�n�_�t�s�x���i�,�N�������,,��~�d1#�Y�gS��1P4�y�2�ڣ�L���ū1n�쓡���ܩ���K]P����M���B9�P�:] �Y	+a�E�(9�y5 �&�1��䭃*��f��K:\�Ø���s;�C�~�f����%{8fh����zV����xq��̂$f&8Ϯ�����@W�Y�bQ]�&�*�=��1%	�A�qN��W�~���̄�s��^~�Hl���N2�ۏ���wp�~#<~�/^��y���}�>��yWT��K��m%��黼�7�^R��ר����g��y=ciϟ��pD+UTw����!����h~�͏�w�!��y=?��c?L�ǟ���CMaG|�M����c|xk�Yv��^c��<��~1	�{�c��7)�%�E;�m\I�WI�W߲
���D����{}�q��%��7��N.A^6n?*�7����ѺsD&Ǡ��>���_�����x����C���=��/��?�>�T��佤'�����Uk���71�cΐ�PI>B�փ'����4���"0���P7�u"P;71eIp���6<�� Xz��(���=&�t|�H7�=�<P�w�V�%��|d��XU��\�j@G���1m�%/�v��#��	H,x�L�F��M�gi�' !�[%0˟!�i�؜��aݺ��zy&��?��Y6^ؖ����`�h�Ph����&��n����\�i�
��s'��!��܎ô�AX�.��� ��R��R�v[c�Xk��[�kKqm|*6NK�ŰP��j0��C�i02Z�11�I
,�Sc{s=����T?g\酯&��a�i~}�^���ɎB�ߑ�����X�9N v�#�ϴǻ3���rw���Ͽ�o~ꋪ_��o�Q}g���c���N/��Y���Tr�%�O��0{A�g��m�e�x}�H����ý1x����i ��o/wA�ٶ��r����w��β|?-	�����X��Ĩh��q����&��84/�T;����B�� ;z�bD�-�H��D��C}��`�&��^��������	N���5Z��wՒ0�c�T�ᅂi�TBH�*R������	�.e��X!���JxzHѬ�=���$�HЧE�ot�F�(/$��#��]&bL�L���©mKpz�\;�����w~�A�n8�+��_Pi��o��˻x��g���+������x;��êe1iBt�����i�b�k�]:�E���ѡ�-��J��S��a�����p�8{�Rtjk���Wҷ� ��Y���GBP'��sH-�)��;�Ԅ�6n��u�� ���:J�Ҁ0�6|"���s��v޸���IO���]p�r ������~���9e8�p-���{�Q��*29$��na8k���@\0R����|p��W�p��7�bq�7
Wu����3u�1�ɇ������!ע'�kt���Z��e�l�:����q�1��C"H�<���ym�<���El�6�ݟ4y��X��Tg�yq�87f&f����,lj��{�1io����q9�Q��1y�'a����GH��C�H	u��rW��Υ�ss�B��&�l�z@�b�8� �C�tHSgC�p4S�:���'u����6m�)�X�a�����;��	yb�AE�f���slJ��%i��VA�����4̐Gb�s��lJ#k��Fpi�x�`�+`��\�XE��ĳ�#21sH�.h����P�<>A��vq>f/MC�&>�t��!���so�]mHt�p�qDB<5[�`�L/9A�������	�!��/U�:���K�wū�x^�N���kxW�
��Se4������u5���k��*S�yl�ᛛ�(�ܜ|<���c+L�g>�'�3��wb>�ׯA�˧��?��N_BY�	H����+кwK|9�z/C�/KѬ[S��@BeSԪ��{as�W����|�1�wn���8y������������X��5*{� "�1`܊4�TՊ��R>2ƃ[(D��_�M|���P�t��X��d��l�w�g��:��|3���L�<z�
�
,�ʮ#�����1ii�L�AY�4u,FX�X��B!��!6�z�
�OGت$�e㈉rA�]�Z�wDKj���ˬ1��k*��J�ZXf%�k7Ї���i���T�&Ua�R��VQ��F��z�����6&
^kǴwl,?'�cb<�FϤ�cb�g��MbJ�J�wٲu5�yfkZ3�1W(�Lֳ&țn����7K��2�yT��'`̠��ﶵP`4�=%�Tr�Mp6�M�7rGk/�K��������ׂ�5n/)�����e��9zx
�?�எ�S��Yh�խ}��[Ό���3������d<ݛ�W����L	^�i���+��Z'�fO��^���^�IF�WO�z�	�^���z-�Q�D��]A����X�q�Qض����j���Q����)��v9-���e��\T?��wO�t�,�}�ѹ�7�����/�������t<#�}�:?�L��>~���	32)Ǵ4'�웂�ss�~G�v�������7F�iP��!�*�x�	�����%ap��8��6H��'<�ɒ�� �	<��i�X��\m�RK��DN$�P"�F�R��w���s���=A}�:�wD#7!s������o'G��*�꠾�����m���L7��ҳo����aň^�1wNo[�o/ţ;�����x��W�~vO���o]�ߜ�5�~��~\<���;��>�s'�������_tGFvBCC����dD��E�s �\�����`$FD!�?���$*h�{d�'��|d��J%jHe���g-�_!Od����yQؠw��	J�	T��I�16	������%X���Y�g����o��P�zo��1;O����-:Ы�L]C��HW٠A��ZO��DX��G��oS�u��)��5z~���p]*�M�����
Dd�]|f���F�	�Rʝ���N�q�#��nM���C&b�_]�R9�(��!� A���O��4y��Z7ZhxM���I�xM�z�-�ɛG�|rx��)����?K�B���7�F� .<	.�x|)��� /�� Յ �7�u48�XhS'öl'4%[!ϘQ��嬥s8�,p6	��u pʂ"�ty���M��큢x�(=����*�5\V�2}AX�!pY�2�#�}���/���Ý1��v�,�+���V8d΁�g��\�&��r	�>j������!���;if�g����ExS���uba�r*����_���~�h����M��Ĩ�Q�7W����F��7	�~�j�V��:��;#%��:�c� ?�o�+ƽ?���c����\���	5X�{����])�ѺWT6V����6}��=^�z�+w��V���<}���?��lbZ��~�Ç0c�ĺ@߾��x�s�����<J�_����1�����#�z�EP^KP�r�ʱ8uu.�_���ۇa�����p(������ݸ�y֪͐���W�ySn��?��kw�����&6#Y��]P��F�� W�|�h�'U_P>����[��P�`�>��,����T�Z�CzC�����5�䭋��؎�9��}f��J/���Q_�pw f��F\��Zz!��(�[b:��A�9��hDw�FQ�Տ�` �=|PbpF��>%��ºV���5�l�Jw�%��W �&�-6�`A������Y�X��~�XL���xa����Aa�;�B��v�[��^/Vb	��zK)͙0-�ꏐ��*�uB���%�d�������r����"=�Y�x�[N�26��XFк��g�����~�&b�ږ���&O�iB9&��l<�Jc��C�"$���zZaa�H�+�Fc��97�w>��T@lo�{˚bK� �JT�_	���0.�S3����?���ƅ�!�a~A]>^n�Wg���x��`���`�����rPUL�6���q��.�9A��%���2|���x�b
>0 �&�"`{L�>\DB�<�4SZO؜�	A�}��>�e��o�y��2�3���"���cZ�|*�|^�9�-6�$����騮��7OF����xq���  .ţ5���$��`[kwLI�aL�kZx���4Tm+v��y�q�Ŋ�Ȗ���uU�����i!��1�Vχ�K�� G'8���@�4yv���g��뵐��Zfx��j�HdR0#)��H���X��pvUZ���#�6B�X{�yX �*�([	��h��&)��e�pg-���Ո�.$Us(�%�ˎ��ͱwbo�X2����+q��n|}�.�9�G�8r`��\�]�W�஍ػuvmX��f`ьI�;i���������hD����'��]�gKb�g'4H�Fr\��XD	4������o�Y���;��������Ze��hfy<���`����XuP�Hs����$l�9�Y�o���N+5�)���k�6�!nM��m9M0���+�F��gu���R�h��ʇcEE�*���e�q��d|�����m�d+	��
8K���$:~��7���G]|o�{���ct�o��/n��ʻn�K��Z	ipE}�Ar9�d"~,^6]��0\t�i��G���Ta���Qحt�Y�
8(1�iya��"y��(L��Ej��?��[�p��vPy�Xi�	�����p�j��|㱺IGh�~�á��i���|)W���~9�`Yx����G�S�ĕ@�� 2�5� d�a�1����i��>o��M�b�r���F{y(�րK��v/HTIӠi����f� ����� ��0�/<��1�x��"U��q9�!�ZQ�F0ϲ�P����~9̯�ɍ
�C�{\
]{��R��7�DEc)T~C�Z���O���p`y�<_��ᕫ�#�	�����6��c��r����aR�Zh����d� X��nb$5�\ѧ�?�o�$X�����ݏe���'���g�:�Iu1E%��i��U��Ysb�&x��?ۉ7o�Py�U/��}�g�O���������^D3ر������ݺ�Nl��Lx���/��c���>:NX
�2�o\�I�f��98}}6�E�GcފI�=f8��u�OI�g7FN�/p��%^	�>U'/f��w�N��O��lwLY�m��@b�8du���3ұ�`|sg"�W�#�����F�����zȫ���
{,j�6v������Y�n3�ݱ�TG���~��M#p�z��	�v'�'��ub�V?J??]\�a�n�.-�F?K-�)эZ���

Jy���k[��\�0,��Q�;A�!���r#V8�J�/pk�$��7 Gzá�C��]/����t����p����6X���Q��]���Ɲ7��H�*Nȃ�9����Q���孅�)O먢b�C�	��!O��Z*�WZ� o�@�C�*��S�6���
Zac�a!Ϟ@�A���k0�J��V�J�m��l�}EB4Tqh��-b�ݟC��Nŋ��
�����k+B1*A�>�UcF�+�u���aq�/9��c!�p�-�}o����)MbL�VM��f��2(ZWE��q�K�)����h�P��,�{0�f���xyk�n���'��7����T<?5/N��c���X/<�Ӆ�g�:��t{<���7���-���;&�U��v���'����^xs�@�� T3�~���Υ�Sޞ1Y�W�o�͡r���l>|7�/v�˃M�tK6��ݚ���c���S�5X��W��v����~�^�[;�W�q
+�R�=��G*A�%�Ol���c�( ��A�0h���$|<V�=v�#d����ZA�'�u9&�ꖉD&�X���A�T[����5�pB�$7�M�@I�-�ꅈ�#3�9���`��Hwj;��� Bk�g�E��f%`@�,t.m����0�[gL6S����1l@O��_vn�^]+�E���ӹڔ��83ىQ����CCP;(A������a���뇤�p$��Ap�']��4Q)#ȓ����|�,�;zf�c�STJk�̀���Մ<ֵmi�e��ξ����:G�o��J�I�x����rVD&૑����ꉽ����~�8��?��ĭ%Kq`���*���x����%���v���g�M�>��4*d�4�t�tko��{a��'��p�;��#��?�#����ژE�P��ɋ�2f��'�����g��XVw�-��QS1#$�T.8��Y�qHĴxy��b���C�F��I�G���R��
{L�����&�u�A_�D�i�Ê{#��PXgm�����B�E)�w���j0\���L�.wd,�l����BWL��@=��A�'�t�i� ��
f�a��⼽��a����l� N�q�*��6A�A �u�:�e�w�~�<Q6��c�8fp���ʘ��:x���wz,Ȣ�����tml<���p�&�;�O�N�%��0~)��K 
�Nh^�K�eb��욝�����_m��⵽�#�qx�e������2�?����bq|^]L���/���P����Dk����;bp��B|�c���wt�����u9�V5���-������-����o����A���S�/�V�=��{�jN5���d�<�IdpǦ�Z��������T�Q¦�����?��/欃w^;���C���/�Djy$�ۧ!�u.�+[!�y+�k�~�[�+�����;�w�_䝮�c�Rp��Ƹ�M	~~X�ۯ���ݶ�|��O,AI�"d5+AaeS�1��Ow���L&DٔXMU�v����TSj^����0M��j��_���A�� �9>��Lƶ�hV��]����xH-��V���{�1�.$>�8�١�����%T���k��Da�:T��U���+�`�W-̧�`�J��L��1s��"�)���F`K�
|�w:.^���&��U8��tl(艭qj���
�g�¡N#1�5�TFJ�A�I�1�zln��A�i��3�3��3��[J�	�� o<��[�}����Et.�}*�=�B�w���0�*�nbK��H�7;C�<�уÆ�nx�.�ԏ]qwq'�nQ]B�'J�(����pfh~����+�����\T��xH��r�_MG���x�n^V/�[������C���h�y�S�g?L�#��f
�_�7�����x}t8����{��mpo^[ܙ�������M��-���9�88;������6;[��6z/v��Ʈ�~���l�Ɏ�1��%�z$�P��8�?����ܜ�
�-��r�p�A��u�L��O`JP�~	��F���`<���ϴC�1jx�-��u��ͤJ���5XX��B��s;��8����G@=�DK4�"� ���cc�X�-��0���ЩL���!��c�����V*�P(�!�	�>�T�$�`#����1�Pf��ho��@CG=Ԉ4J@�����HHd�eP#����^�Xo�n���F{�N��s���jy���L��}��7�z "�u}��z�W�6b�BE`������{z�ˉ���\+��HO�#��6�X�_�L[)W����?\��<�L,��pg3�{���E��ت5A�6N�=B%v�s�'�a�o-���?�͚���y��w��@����ʾ�<`<N�ގ��6aTV#̩Ukc0'� 7�N���|�4�S�,�i>"��ڣ��!62�z�Y�QB��R*�Q�3[kOkDP�s�5���D*����8��A�ə©���oS����ɘX�?@�>j42a~Lqy�!Oo�<���Lb��Yd��:w�K���1s����8,/逡E�>B����;Q�� +o��.�'3��*"����w�2���B���{Ƽp�^ۆk�%��1�+�.=�E�~ti�"L��5X��-��f�6:�	:?ˇi<��	s?j��r,/���E�D�&�ф�h'$�������E�2�c]�&M�gȓd�5���-�&m�E�T~^aa!�Lh��%��a	�ߍ���y>��]�w�'ȃ�O;��e�pnM�����([fD�8�J	�F�:���X_��}��ig$����om�~KŽG�x���`�����#
𦺄j�xU=���,Y�_�p��/�U3�N����|�_�f���&3�Pag`�����}L�AޯO^�ߢ��)����P�fA��4S�Рni����[ÿ��͐޶3��8��w/ؘ�`�=���3p��Ɣh)���o����/�>mA����E���i�nC������5A�"�O����Ck)Ԕ���n>�<��_/�ulx���Kа ��Wf��c�x^���g����H�S�m��ay����޶��a�q*�<����U�2�u8��*tM+��v}0էfm��'�]
l�
ǡ��1�y�����6~�����ݠ)6���ݽfcNVg�	����r,�r<vO\�}_L��HlS����� ϒ �9K�z-e<譡���fȫ�e��̳4A�N�՜˨�YB�,�y�[F�/��3�c~�6��a��X�6<2g�R�;w����y��Rk��Q%DKo5�g���S�pnT�m)D��fx��6W -@ҿƢ����PYR�sc��y9x�������_i��7{��O����axy,^<��7�g��3���K���槹xqc^_'�4	�N�¯[���-qvR#���7Į����)��aE�H��	��h[̎wƼޘ�����{crg�Kp��:�X�}���_���
5�O-zh޿�/�j��P{���C�u1bH�#FŸa|�?݇`,)���/������yUW���7�\������|�WO���1t�������\�5���M�|=5�F�`eg�ɱ��uP��p�.O���L[dH��8���D�*�ޓXz�l�3���yx2k��1�	fY�I��S�(��c�@�i��
y��y&ȓ��4Jz1�� B��i�6Hs�E������C�V��%"TR����uR	��,98ZYBE�Z�6r%���*^��Z猪�U�@(���@OD��P�,7.�qhܠ�$��8>	���H�]��cQ�����8�DG�]��z5��Y*��KD�*�H��hx�xf�cP�@����z&l���/3�}�jz���~&y��;c��O��Ij����c����K����8;y&���Ş�"�k5����O���#��dNS#��q�Kw�ز?-߀cu�{-��	�D*��F���p'�c�P*�����-�F���@��P[OU���~$��?�. �q]��\�5��Y�VE��I�qy�������r�� �z[i�&Lތ��[oeC��=*g̎m�SC�bvZ:;Fba~k�뎠��`���/����qE,~�������d��`6�豰J�i�:������,�m���DL 4V��@���|:.� �@�E���nWw����b����t�Ϯ\�8<���C��*{3,�'�Sg@����!|�/�f�%8]*8=m��
QÍ�c
�����e�D �N����@��/~,}���n�Z��k�aH3GT�r���������Q��r+@.�Kz����^c�<e��U0������n�1���`D?��[SK^+Y)1���R��j=��{C��{
�x����3I���u#T}(#����e���]��j�k7o���㗯�!��ޚ.�Z7���5�!�y�`�=����>?c��9�w���yn�R
���Ko	���&��b��pkT�C^@Q���m�����g���¡��q�|�GC�z��ߟ�෇x^����W�tĺ���z	R�ƠI�r����{���U�9��'S��>֤@�|�M��j��	�V�g�ZC�F�Jg��� �^�L�F��8���o?L������8ԋ �����a.��g��R-�[��Y��!��ЀZ�z��T򚼕����ƫ�%hb0�
��qq�L���A'O�!P�F�f�+F��bs�8��NN]��1)X�w�\��mAϳ�(�w�BR��T� �'b!��|�*�b%�XɱQ !�c#!f|����cQ1x+[��	3�XFǯ�c�q� o�������1"�>*�B,��]H�EP7݂��R�E�݄�h���5�	���)�ú��~N:p���TbC;/�bz�3v��3��ޚ4<ٝ��g��͹���R�g����}���t3	��4t�& rU;�Β/���.83�)����N)XV^�r|04��b0����8�o�ztu&hk�G3/%���Q�B+�ۢ]�3�	�J�4��S!�Y�d{9�"�Zm"�A�$'��HrT�Z�x;%�lh�#-��9���B�����sѠ�E��:t&`E���%���1�Ƶ���C��3���	b��ǻ�F������rG�?�
8�
o�4���R����d��K8^mk�}���҉��B)R�&��$	� T�G��Z�u-��U�}��1��<�A�˟�nkh�KF��b���R�%r��c��qmV��X��Z� -"�P���!-��i��{���]�j�oT4��"��)6�wv@]g'�::��gc�pWDz�"�����l>ȉ
B��t+Hƈ�Rh^��z(���ʴDt��F��\���AA|<CC���� {������-�������V�L�[�K؜]��e����^h�k�u�כÚ����X����^�BEH�'�b�ޑ�_)�f�����O�8`��ךw�é�h�j�8q>~�gZũ�8Ҩ��f�>x�l��9�?v���V}p�>?ɜpQኋ��0����j�3�����y��ﷁ�u��0:"�ֈ�t��]ɣ}'���?��qE뉳B��8'�`���"���>j
fE���-�qZj������!�*#�/��Y2m�D�ǆ���e~q%��b�#�G5���0�aKtw�������a;���>koxaQt��<a�a�N�OX���=7�η38�"�\���&���̙0m��d�ؼJ�p͆�6�@+.��ǆ�x��Vep�!l8�M#p��`9�; �9�k�,���j��f�� ��m���U�Zj��@��6t�Ű��Mhk��R��\_��c!��l��9P����DY�n�3��2u+�1�!����m�jz,��ʉ��$�<W��I�WE����(zc)�3���p�O�M�ƚɮX<��#����� F�Z�h�玩cka��P���{�`�۽<<z�O_eP-��߶��������P�>a��}d?�z�'|x��ʮ�Ur��Y7���5��\2-">����鯐Ǣh�y���l�W����-�sn#8��Eg�51�y��u����hԄ�<�FMѠ��؃�o�䝉ǡs1��S�y�[�c���D��(O_��t�T�)z��7]�`skL_�'.�{_�G}`�W3s�[&s~��n*S��a�?l�x��ʖ]�C���ۢ�`7ܯ��?������*�1?�6m{Ձ!�.�a+#dT�;:���	c�*�H�E�E7�+
��H`���yMޚv}yM�<���x�K��.�Ca��4x�$c��-ZIp�*�����]�&a��U��k�F��n�,v��Ѽ��Ц溄�.�ѹ�vp�DCs;i;�6K)��>LX��?C��
X�?�<)oP�B��.L��H$�4Ol+���v0�
��*k0��K�rZBiΓ(0G��e�0G�Ck!��ymC��,ơ��x��ovTbmt�xK�3C�x9�KW��KQu�	�\���k퀟�?���~�\����{��8�/;*�,/�b|0<�}�\�=�-\	�\�h�"E���h�m��>�(��
͞@�F�Hk+Ԣ.�BdR� Em�A��O'������������������Hs{)G�d�pV��$�����^b�%?wRJyKG�~Z1�u�R�J��B�^�|jq7qW��Q�Jw�������S*�.h�'������'L[Ip��0����N��{��wW�����ޤ$%�w��}��js[L˴F�%�=�,jddѻ�b!D��%yI�>h�����ө�<�0�c�`����b�5C�;�؊��R
�������ӻ Q�!�}�J�@�F�z5�J�P��M^ՍB���h��Z����ZbE�^�ԡJ�롶�j������ W;��Ez"3:���P��9	hK�*=�������<)9�QT�r��M
FL`B���eo'����:�--x�31��s�"W�p�`�-���h4̐�����g�<sW�L��k��ֵb�99;�8D���2KTF'	��XqH`��Z�NŎ�"l�-���EX���!�c�Mr;�𨅵	��լ36g��*�H|e�K�����}L��Eb]H]�s�G,�����5$�m����q��ֈ��'��J�9��8��o�p�)��68-��	j�����.k,���iqe�dL��CZ^�W�j��=B5v$n�ey�	�L1��XC�b����%����������1+��r:"�>���sy�!,&�+:k������ !@����S����Bj��@M��]to�eφS�Dp��vaZ1|��oC��Bb�"�n|	�B6&o-�)��>�	A�!o�'m��'d�6�xK��3�}���<Q�Jk��\F�Oh��aȁ�#*����v��>~,?&���\�W^����N�c���H�p��"rBz�Iq;l���b�$,����=��o��<��_
-�V@�,� ��3'o�5���|�;A�+�rGQnb���@�7̞VE��7I�~+�2�{��_6�Z�-��ݧ[��D7
GÖ��:�%��[�/n�_/��S�-�Z?�;'�9��=���9�آ&G�ǽWU�t��t�k�284́cB:B��Pѧ_�o��^.ʃoq~L�<���y��GM����(\�97��'���/�p�i�xZ�Woۑt���=����H>���;;t�T��}����c�_��=y��_<�۪���l�c`�|{����Щ����d�_S��z��6�T/Ş���U��k\���: �Z|zhl����@����R(AW��uNT��x���O_d4����ԯ�+����"d+DXet��N_`G�^����ؘ��uٍ1!1��e$V�����Lr�����T?�+��u�r��{,��@�M��C��pi��C6C���G^�� ��|!�C���1VZ�B�1YB��T{7l-,�!o�o�'�cnV�XQR$�<�l��,j�7% *t�}��rXP.�׳������Xt��fT�:)��#�;�o/tě=���wc�۳���a�eQo�����S0����n6ȲѠ�^�86�K�@4-�!�
Չ��Ï*i?��r%�DV���OK"'�1�� &���$�Reh	A���l���Ij��D%���DN-e��������~4"1�/��Υ&�[ �C��_e�p� 	:9Rm�h�f�6����sx.�_�@�;�Z��Puw�=;G��d7`O'<^�����2����Mqjp:z����g���!#��A^Fp�������6Fؘݨ|t����<&�u������ug�9��qx�Zyȓ�`%�C@�+R���bz��j#����*Tp��J沤�_ gd�wǎhӴ�>�P�;�g��z�Fz��:x{8��!��	��<��� �S;Y�I�C@���O{�i��ӹ��(�LXޙXY	 �bZI-������P�Z�)�2��?C���{��ٜ��cd�LKФ�����h�Aǈ�L/��-S�ů>$��A)A���D�F�~�N�ث��Q�;ND��@��-Nˍ8gp��/g�<p���U�����wš�68��_��`W��h��8w="����=�T�M��/�#�V�VA�X޲Gz��¦��c �e5�� ��Q#�P���N|w��pa�����?C�+=/�E�9���� O�k�6�|#y*�%x\MT�Be���!�1����. 32
0��B��:����A�iX��I�i^��"m��^��J��C����P�����A�^Ϩ^�	nN�!��.p�ǌ������M:_ .~��a��k���,q�Qy���[����rN~�<�&����Pgy�xȓd.� ��Q[�/4.ua�;�������Ň_�&��"���%��y��|��a�q�̡�X֛ ��^�ѱv.�Į��غ������%�s�
5�:�;�S��FB����[�'K�z��������X2��$��V ��#J���>5GO&��7ɸ�S��߈آ1�l�u���hѫ)BҢ��$�V��݉/��ͫ�	�^���3" 	���>O���'&v�
L�����l��z>�g��{�&��04lm�Lx6HDב8}y0�=��@V�n҄��e��A����'�e��;t*�ś4y��ֳ���<�=~�E���m��Y{�{߉Nܟ�p"��o��)K/>B�_���'��jʭ[?�޽;x�</�՘o�YL���Ǯw��Sp�C�>�q��1(��<���Mo��?N���!�����p�L���r�vb���Gk��"�$��1��҈8Nƻ��xH�J��2+���*y+i�N�
[�11׆O��/�cKeg\<�z���J|=b6�E�ؐQ�C��船�?jN����I�X���N+f]����JaU�l�����c�{[�Jl��@U��'P���7����*�c�O�?i�xg�{�V��pP�D%D66�!g� ���h�''�j�4P���x���ǚ��)zG�uǫ_���[|3���Īv�1� #���#�%vZ$hԓ��ӡ�V/��R	�$b��zW��@J-埁���ZDbE�K�YR#�3	G� G���53o]��c*-�lKXZZ�"�m�x�T(����u�zK:����QH���(/��"�>+�~2+��E<��Ӊ�� G���aZm�3����x������w��ć�]����|CK���6���pnD0n/�Ĝw�������@/�`?������t����лm�[�2M�9����S#Ы	yL�g���ݵ"(��1�*2	�,�9X�5	�V�1m��0�_���@@�ź29z&r%���d�@@�����mV�xa��R)�虊U]�N��\�0-����0��Xd����Hl`%���b�����wD�Q�2�j�Z�"���SCi���1pc>��]�JY�_!����[��yf�c>��#�;���j�n��/�ۥ��� }�e�p�8hi�I��r.(�8�cto��pU��%NA ��E���Vj�����%�G7I.Qz'9)v����܅��s ����T�\[8�m��-K0yp�\�Q]:bR���ٳ;�O������Xؽ/�S�4a�v����?'(�;�2�-���ǔE8;z<�����<��D����O����R���Y��&O��2%�D�é�c� �9��135�wG��0�⁊�=C�w��<+<&Ң�bg����5n�����x*\g��>>�!�i��P��Х�]]�d���C�R�#z@h��{>ĩc�,��C�#'�����yD_�m2���9�G'�fM3�5yyV�� m����q�QP;�C��s\�S���c(D�P%��<g�����1�������k�[�6< �t�S���!_��ᵹ8��[�����(OᮏUR�<z﫨����T���>H���l��p����5������F��Z�Y�
��CG�p�J,��������"����lMAF�;��' ���ה���D<�0?�O�S%��7���` �������=����gfsOb5��Ǉ��m�Zx�t�CvX�� 8#	7���w+q��t,�2 ��Ch�f��<�Fe����/\@U�+p{O�e���$�p/w�eᏗYx�2��6Ë�J���5W���o����Z7�8�e�)k��x���@�u2k�̐w���s�W<{μ��x��^�tS�ܲ�|1flBc����Xx���?-i�8v��W�F����k�Y�Q%��9���-*/Բ�D�n[����JQ I}�-e���NC���[����l�В/Ǻ(���`oJN����Ğ�f؟R�#�q��`\�<WzN��/��X����k*���3�'`���]��������W��N����<�l3�V*TY�y��s��Y��z&<���4=�Q2o�<�yU�Smݰ�����!o��4&o)��
�yT�,"p\H� J?[̡�����3��'��7���/�è+\���';�����=��_��Y��o' 7f����޹!&$�����z����9�I9�S�<	��hٙZ��P:Z��@=�;��DA"'��Q~M�'��`�w�B��
]?���2� �,��L0�Qx��P�	�&
k
�$V���7�F*�	����y�,�.�zv$;���K�u�X�5Ϗ������5��η����p;��&�{{bn�{��Ǝ�ih�&BAd�H�R�y)1���]�̍��^;k#l�Щ5ppp���=6F�/6��Y�*y1/3�1�7�8c�0����h+o���_�@Β��,�>���C��ƺ��aP�I��O�f�"/s^��ДR^>������?���e�"���u���97�-��|���Yv�ɱ��S���(ܙ�lY���b������
gk�IǞ�b�S9��G�;.��y�#��#N���ڣb;jqR��)��/�����i�iK��7{��ݓ5�H]���d%A!}����1e6���5aTFq�_�?�<������O����ܢ���K>z��U��o�Y/9n�qy�\l���qX����R�C�j��{���ȉ�T���J�wVB0�v���̀C}�Ez���6�I2����P��'�3Rc��<��s�pi�4,�k��v����ŕ#��=����Wt��$y�F'�(�"���	��������*�{�Qp�_���|�Zm�2���>�mQ�
,�<k:D�+a�d5,���Ș	�S!$	c��_e�jH�SEBlU�`��7�"s��d���,j��P�����O�N��b.\8�.�ua��G}p�a0�f��V#X����V�)�!�]1����5�\�n���G�e�r�.��f�;�-tm�3�ply�Ϋ���cp��;��8�P�*z��Y�H�WT��t���x��ك=1�?�N�����D���i�>  R��$�ڏi��a~{Q��wK0f^�f������ah[�8��/��׋���5T�z���̣�j�z�������*���3�w���Ŭh��S��(�%���:��*"S$16���O�r�|x��[vS8ƥ $%	S���+q��$,�<�GtD�V��Q����QF���_}C�ܮ#���p�]���?���߳q�q�(�S�����U;<x�/_���'��U��0�Շ��C<���j<�`H3��W&��a�?z���GM^�H���޾�����cĖ��><6ua����pmP�:������b���gF��v$}���]k5
m�QI-�No]�:h���A0�D(U��2;m�[��B�:�k��J�)J�&��6r2,�TXep�|L�q�Z�P���
�p���ҐX^�!�m����0�?}b0�����
�����@��Z��VS���*�T!2��6�ۨbXG��T�3�G��N��[ԫ�7k�L�' �S򐷳�v�H���J#VѶ%T�/�V�B��K���#z��Ȑp�t��O�9e>�fn�K�7�#���'[+����G:��q���� �M��qdp>&�����VȱU��Q	w6�� (@/G��a:;h�k��]cr�ʴwl,����T�;JDp ����A`	�Z(�����@�i�L´r�]4�\D�Ŵ��cPfI�d�4�/:���BJL�>�Y{' pc0ǎg�;�m)��ȭ>������)ᥖ�c��^�	�<t�꬐f-D'1�����P����~�Y��Y������P~]��m=���K�kaX��	�����e�������N]ć�B�o \���2+[-x������c����s7��P�}�r1�2��m�n�,&�jJ�}�������k��t��g��,5!ϜFM1iY�&�c��@�i��F���}ܗ���1z�wz��ZA���v�vu����⳰7��y�-Q�4#Y�����Y�)qN��y�g�NRc�}�'D�A�i���N�he��"#���ƸY��g86����!��CGO7��d���;xA�w��]<|z_�=���pTFf��1sq�Mw�q�%A(G@I�i��;S��A�:�Y��q�8���5x<�1��||޽�k�f��r�8�<����b�7�^"�3A^G�?�G�aQ���O�M�:�O�����<a�ݐ�·exXHɽ2a��\� X%/�,� ��X��� �����AM ɘG`��ҵ���ؘ�S.��'C�h-4Ytl�A�1��7���0ާ���y&M�A@�y��3�W�8��a~|�&����N[�t��Ka�UC�6p��

�Xh
�N�I�F�<�&J�i9���^!�Ƞ��2m/����]ڴÉ�8�&{֦`�H|=5���=�� }�υV �����;w�
prd.lj�ţ|�zJ(�O�@�F*,`��Tg��]��p�8��1�7����*��[b������� ��EE�|L]�	��Oŝ?n���.�R���y�X�82�N5����Yq��_�L��B�����~�}'�)�\��Ѡu���k&a���y`�홃��#�M%A^+�.j�Jj�}��m��۰�+Vl�ƾ��z3���r��1-^;<y����\%�xZ�_����&x�~0^�݁շ��W�LM���yf�c�ǀ�:����/������.����yfO���g��C��J�]\.�	�a�˂m\:��u�X���c:���
�͡��VF�J�0-�^�.9z@u�[���3��:S�<3�.��K��a��?f	Lݟ�{sgE���Z�*�g�fjղ�ӭJҌ�6[�6`�ʈ5ZGl �\�����I��*��*��c�T������U`�V�	Z%櫴��6�yUl��j�6Ht���]�&a˟�u�2�c!��x;&�ؙ ��5c�7��� p�B�K�R�>Sn��B9��:Z�"@�M]ppP}�p�0%O��k��jO9�l�w'�������'��i]T�Ȑ��I�J���pV��q���l9�#��!N�����Z{5�%|tb��%��!�V�Pk)�l�GmO��7�`��tn*�0%��dL���Ŗ�������
�('p�u�8>��w��w�\�yr:���3�����NBp)���JG�
.5܍*�ڨy@��e�g-G#���iP�~�x�A*��T�ZZ�5m�;J�$�Ã����(z�W��v_����V�����>!k[�cF�#&���)�r�i�����ϥ|7qvAI�H�թ�H=7'g��[L�� ���:�5ߥY��-��b��k��"f��	`5�m3˟������5�c�jjk������\���y.����,f�c�Ǻ~̱.e���Y�G���W�ʴ�=&l�i����`k���#�	�'��`f�?A�Q�-Z�q�����#G����)�)��q*#���YZ��S�q�����̈�r;�+{�a�k�w
4��>{�a���AzZ�l؏+'�a��5ؼn=�_>�����W/aڼ�HjP� �p�O)÷�f�LE{���yL�wX��'�c���j\�y����M$^�����e��
{,���4����B#6ZRYGe�B9�u�pf�$, �ko�����i����`���w�",�A�s����;a2|ht��uP����'�0p�`p�e��:q�>�J�A���k3p�HX�����py�!+^O��
�hظ��=sl
7C��
����ԑ�l���m�mq�`Yx��%��q��VŦ�d.g?�]d�"�w{p⺰�kM�H�A�4�Q�!���č��i��$���9�|:̨���K66�i�q+a���n�3?׶����X�]��=KSpsI~������2���?;q��+���aBs'|���l���~X2�r����.T��]ѫ�7�n���ͭ,ܺ�������%�8(Ž�%�}:�x"�S �G"���F����x�l�����1+ӖQ�Ou�?2���N�X3S00���;������1���zF���uG�GL�0�m�[v!:N�ۦaݦ~8xt N\��q�"������rD��B�Q����� o˞X�)G���|�m��E���1�?-����x���!�{@�����\<}�/ެ@������2.���Me����7{IX딹Ga/��e���L?Q��t��?GӾ�!�=A�wF!��>1�1Ip�ρ}T��Q�0>�	l!�P%��!M�BK�	�:YHP)ף��Q_�T�SE�m�Đ���e�4Gw� Pbc�Vќ��#f���@�K)	 9Z�a5�*J���[G���$,�-s|�ܬ�ط;-�|!�ƴ0�,c�:� P�i'�0[fX밖�ź_W�Tؤ��}�iy�[ȣ���@o��r�3�5y̺�A��X�%�e���rR,��`���
��rtJ���@��څ�v���dzGq856O�����XK�̗�:8gG4��z.��qH$��ҊL`Ǵt8�sRke	�H��7�e�U*h.�������̉���Zz^Az)/at_)-oJ�A^��ZJ�5s�J�@ h��NnI���7?���j���vPO�@E��� ��0A�Q)��R�I�bJ��"(�,؄�SK�\2�Q~j�Z�����<ڇi"ԩ$�WD�)�s��0�$����)NJ��ӡ�/=������8���~�������텸:*˛�b|�;��� ]$@������Uxx�iDR�"x#�J�������Z�&��][S �i=�-Oln_ln43H�!��D���U����	x��k�g����y1�ɟ�tR��sw-�6�Z��B��kךu�l`K冽�GG'��1�����8����/����,0⚕�*�q��OK��n��bZ/2�r���c�g���<�s�17�L��N�۷.A�5��w�����Ƒm'0z�ٸ�8v`7���:�|��M�������C�b|3fζ�5�A8�r����O�ĻPa�w�`���k�XW�!9���H�g�!1�5>wR���SQ���fK6��Y����U����<s��!%k$K�.Q��2�͋��.Lx�+8��%���B�H=R t˄�VOhR��*k%�����hA^cp�8���G�`Β��ka���9��� ѧ�r��&�Z��1�tu!���"j��:X�0��'�����j%g!(=����?i�rW�·8��0���u�J�s��:gt�#�B`�y�tX샸�,�)�J	�(M�Ϫ䔩��Ti����H���3Z���L\۝��p�p)�>�8����c����r�KwƉ�`,�싊4euh���v��7���A��oɏFNCt��ekbp�\
A^~���_I��M��7����4����.�cʪVhҡ ��u���Ǩ^u��?�z�z�M^��S��(lb<b�2.�W@�3�U�v��v��k.���6�M�BL�L���owf����(��u�Fd���-(G|��4q�=|b��k�-��#�`����K���V~�#�d���4���'o
� �^����p��$ ߤӭ���UG���@���?9��M��L����<�_�Oi�<��d�ik��f���H������e���&B[�>�N��x��6,�J�t5�Z��T�� �kEp�TeD���Tٳ��>e���\�S��0�
�����_��m���2�����,9�8*��Y\YZ쉰�~�������t	�7��v%���!�H ��V��N
�s�`�њ��]A ��k��+�_<�kD^�g�K=V�?�)�-s������ص�6U@?�H�Q���<�Q��D �5~�Ŕ���2<d����S�̓����}Ec���o��ۡ�@O�ꛁ
R�V�UKF��#��MΌ'X�*f���]�ll�!	�Re"!В-�|Y@/�@��Hy��cl�".�&KX'�5*��ML��{z�M*�cd^��m�����xh5pQ�aˠ�(n�L>slr-Bi�	(��k��y�꣈��VZFk%l�,������x3�ໃ��A�>]�K��c�^c<��o�Ѝ�ۺ�����x2~��g�'Z��4���!IjTjш�5��(������돞s�w�=��s%a�� �9�<��c@Ǆi���5?g�ŀɬ�c��1pb`e�/3X�����!�	�Ug���c���s��^3��ܷf��u��ln�K�� Ϭ�c�9y
��=�����j�Pku�1x�vt�Lbmg��3���0.�� ��	x�ѷ� �A�w���8=�sZ^�O��I�-�(<xM�Y�r��lp^��Iض���e�v�>���ӽGa�{��آ���������Op�����/����)^�y��O���1|����)*���ŉ�=��%'4��(������	�$���Ÿ4j���!OL�.��q*KN�	F�qT憃
P��ځ��`��s����yL��XfĜz�8=|*����2�ý����2rG�.k1�,��O��,=FtҲ�Ж�N��G����`.�y��M_.�K��Ӻ�!�t.��:>��a����{��d8�6഑���!w4��!-�E�xغէ��Σ��i|�0xw\�y�\���W4' e�=Z//;]�jp���I�;�!'�{�E� ��6��է�Yi��SZ\�����g�<DM.����S��,2v�]
���лg�������}�	.��ķ{����<Lk�B�
�0��C��ѻ\�Ƶ8�+p����8���ʼ`odc�e��
@F�/�t�â��}$7���w?5�����q.�?���T���4�ӧ-q�h./+�მ���i�߱�Y��ԙ@����5������P�����$]����Y5�P,,�Vs�{	���?r��y����n3v£�K�紃KV죂�oDK��kP�~%�_���;!�K/$v���
��h���V�SJ�� ��B9p�^H��	��m
z�ֽd�}��'U�xZ���/���e<>��+��%���ӱ��l<y���u�_o�e�|<1t5��+1�<�}|UUp���Q��#d�։�MB���yi�G&��qD4lSSִn)�aE��Hg�V�{׏5h��Ӡ�*�&
�NHR��U(�U�aVr�����J��J�D���T�.��H�-��{!���ؗS�δv,B���M�w�2?x,b�9L�
Z^L f���Э��`�H�QF�9���I�޶J����mL]�T(������"^(Mp'0���WQ�� q)�yA�D{l.j�m?C��a�<�Kb�<���yR�z�M�F+*dzEs8;!��7u .u����81:�B�Qp�������52h	�xw$218�������|��(Ol<��BL�gEpd��Y+A���/�,,(�mg`%dFτ�Ja�7��U��@����R)A��}
�WM1�_a ʖ�:��ʙ��,l)t.�L�s�z~�U^�1���1����;���uԠ6�}�^����u���ǻRrpk0�_�W��Ŵ|�H�o'C	�c����Uπ�.D�o\�6�4y��j�F��B�Y�1��:�f�	[g*R5ż��R�jB�9Ϳ�֙A��`Mȫ����Yj�����ք������1�3��=�� Wg��l��1k�B�Y�yj'G��z`ra9��6���U��� ��Mb�t���8���>G?lֻ��	g��N��k�jB�%��XJ�G�w� �Ix����Nű/�c���;R:+������fe�+Sy��9J���r�c�'m���_0�^h������B��X�Z� ���B�����`��rH�}*_l�	�V�Pl�;`�ґ7�8(1��=Vx$�T�)�\刹1�83r&�T�B��.�XP�	���ᒿ��?�`QzeyM�A\vr���p6�pL�K�H�^G`��ȱ�4�����V��P�d�)�%T1��o8�����K��fA��%��(=	Y�>XE�@K�8���g���!(�B�y�yͯ����O5�5I�	�r=:�S&A�����I��x��O��GS���U��,9����!l~V����^ �;i�s��p9��L?����h�����ѥxz�Ϯ�����6?�O4Ŋ�)H��P� ƨv^��O��_H�E��Eq���&e�n�=t6H��p�Db�Z7#0���bq�Z��%<�Ó'�H���uc�|������J��6�^�f�����pf>���3� $@ۿ~�|�%6�v��&�A�Y��.�ݬ����MwK�<����7�>s�By��3��M��>�e�����"��\�f��c^ا��;5C'�����P�m8pz0Z�i��֭�Ц3"J*Pҩ'���Ǉ���܃�7q��l;P�ç�ܥd|�C:~����f��<y��'o2��M%�/�ǮF�IРiG427��,N�'����u�����%�eSٙZ��B�<#�:k1�1P�6�.*N	�0��ҡ�H�1.�����/DpI$nԲ�
�
h6�����5���"R)E����FLcTG�A�z��դkc�7��Ϡ��\�&f����eZ;��*��$�����ɰ�JL�'�#V0g�,-�|e1iwZ*y�S+��������uJ�R�)|w�fNM�����J�I�X=��ũ]ByZN��TɬI�i;A����Ɯ3��D���� �!ț���!o�G�[H׳�*�	
=*��M�X�Q��"�ü2[|;+O76���m�b{����	���� ��A@�$��(C/CA�2�F%4t�Ye����1+V3}�"�|�je�O�dއ ��"�Gy��~st�9!-?Z�����WB�dVR���d]���3�`�"aV�,�����e&l��3��}�X?����yDV�<P^,���x��.��,L��4|Zτi��ላD�@�����+9t�b_��9��}8�����.x��!��u@�Hr%hJ��R$A)][��p�k�C�3A���j��h��@�;&f�&l�l���_�IMP�)5�	[���G�W󘿃<�o���1�y�9��;3��W6.���_!�zl�� O��AO�Ǵwfa����G��7���������N�7�v�<�P㉡7V�b��{i�q�#NН�������$�8+ ��8/��u#����Z�os�6��կOp��j���.n��WN|�3{/�������o�����U�o����CX�����ݰ�3 '��&M��@޴�:8a튫Z^۸K�%�5��cO	�@̤�o��c�̑��{E���F^�R�+�.��'�O��Ҷh�s�#��o���po�*WM.���	pM�Â�G��A�YX&.�Z���ep��Z�
Ka�\}�^|81U�8h��.��6�]��=Bh�m����ZM�Ӑ���u�~X0�ZY=p���O��pD�x�_�|Q�u�ː��i�+�*����Z]�u�.p��� W8�E��a��6���ο7��&@V�\���J	�蚄-�����(-6�]'K.�D�G�E͇M�4o7��N�ݳ���f/�>�W�f�#E8(K���]"������H\_sl�Ec��x��?�l}�A���3�G��Y#?���Gcp�j*�e�ۃB�����YuS<CK<���ߔ��������N�駑�uk;��>��G�y cU����{^Lݜ�u�c鲐e�ݐg^��@���<��c�/^�ˬ�d��Ǽ-�wu+�Ucf8���9.�Zt��p��n���0�Mz��~yK�4i�����|н�=��WW�Љ/��`N�K������<x�������E>\[<{��K#�i��K`���:��37�>gִd��d��f�W��W��S��el`'-1�c� ���o�R?�A1<�b���]�zj�j�AS/�z\T��LXz8�Q.�\M��	���R~��#U�aZbl����+|涣�L�/��01��=�0�J�)�~:'! �����Ŋ址Z��r>���]�k�|�XZ�Ňeݸ�;������ļ寣��H�K�����)T�N����k��;��̺D�B��� o����=�4�˨�^!0�Paˤ��� oca����^����	y�<1���S[�\$DC[)
Cm��K4��3�,l��m-�pU.�K���@��p�&�qQem�I�S���0L�:����#&0_l�Z� C<�����z<0���|	o�Js�3;(f��ͼ�V�g�ܚ��zgJ�UL*�����a�!��!��C��\1���$�J����D��qv�k�J���YlV�AJ�HsvN����i�q3�`�L�OO@�1`e�w���T�Yf�@����u�8:"���e �]Oz��ʸ��n�FvJ�B��%(!hR#�!�;�����l�l��5�{-3��&�!Q���hT�07���lx�}�Ie�o�Os*����_�ѽ��wM��E���b�;�c]��.�O�'��Yj��4���U)�=���?xL���� �w5�<ގ�G+79J6[Ѳ�wvF>��9jsE����@���E�{ �4k�E�����A�Ǝ�)pDc��RGt�o)��q���7J���	��'�c����z��	ly����67����!�<%/����70��H��w�)��o"������FcX��m2c+�c��8u� 6���c��|�6��慓�?A���$ܛ��GN���:8�s�y[	FGp:�٠��Ytc�vXCP���{h�����y�cc�V�]0�ۇ��Ҧ����0/�����2Q��4A�)���G��^#Ⱥ
M�1�"ƀ#��l�H�i���3 ����p*��&���Σ����.�"�����p	��M��Z3��^�xY��!��EӸ������\��K���A_�5XT\���7p�x�K	��A^��
T�8E�1��@����|�6��]�E��ϬɳjF`Wt� � ��
877� ��(���NoG�G��Yس�=��G�{��5*�Sc�qo)bj��v����l����/�FB�#��a�k��\� ��O�� 4J�E�~��s8_�T�o���w	�^����2<���	��W7�������!�_s��?�b��/��ӧx��%��+�1��Fl��q�g�cp�,EMӰݻ�oߚ��Mz����g����Z×/_���G�/�������~���>|�γ7»�7��t�svc޺�-)�9�n^��+����q��Ft��M��~��7v"n�~��#�y���t��7q��,�<�'NG���P|�m-��s8^����7����X��c����]���b�e��saQ����ay���)����>�&����v�5�����Nf��4���1����T��KDWÒzC��ͯ��Ѻ#�b�*0�:��=�%*61i��M�,���2Ԩ��/�
 =l<<�Z*#B�T�R�b���ij�"%J�l�\B�btr1�Feb��/������Yɮ��`y�Z-5b��e,e�Mhy�D�'�"%@���Z����B&�d�[e�Ժ�E�6��t���4.$N|ȣ��ۨp�he ���]�L���E�1wL���Ԗ�ָZ���u��<�.�c&;x}��>��x�[J�� o�POi��15�$
4["�(Fi-��s�nę����x<Z���gdcc�X4�S ����J�U�����I��)-`��E#�-o�`�h��Fǲ1o":�Xd4,� �J҂���ܱqz�gӪ�Pڎ4w#	��X�8%�d%B-<8����#�À�^�
��e��@�՘��������H�U%Z�-5`}[ll�-��XWjO��˪"�)uŲ'�+4bz���aH��Ch�F/
\$H1X ��F�	Rx?��b!6l� �P��z��W#��Fb�	�S�����Ѻ�xy������on��mC�%��H¡����*k���%-��W�2��K�&QB�Q�R-�$��+ �V@hP�#���yXꕼpr)8+��J��B1��Δ&�Cȉd���J5b��oF��J��f Ʈ��Y�Bδ�����X�[�s�)��gK� ���M!c��-����0s�lɺƅ"XY� ��J��AOyW�65A s�"�)M����5�l��!��3�&�rj�*X���z��E}��HG0j�|�F��:[�H��������"�������� �<A��*[�q�{G46�%ա%�C�Hғ�}��e8A@w�����$u���]���]��N�,u�e��ȼp�ETo>�������Y�8c)��]��nĭ��pw�^\��'����I�pt�b�>�g����[���c�c�\/l�7��9�w�ʄ԰]]7wf,µ��1/$��.�B�w����H��|*"��H*0���a���n���h���C���.V.Q9�V����8>`,��@G_�uÂ-�*g"
B��(,ʯA��2$�ס(��&?@\��-oB_���S�z�2��uGB5����6�Y�qț���6H3�C�`$Ic�ɚC�ؔ�maͮB��*���@����{a]z2fd�O�Uz�`��t~A��aU�=����MZ� Ȼ�W *?ek�m<�w�Z4?��e[^���G�_9-7�9���~�i,�y��/BX|�"��F��ga��C��	ʔ����>�!���tBw�9xwk^��������EGX�Cu�R��2~q�z���va�����B�|�����ܱjs".���͟s�ï9��i	�j�g���}.^6^<�n�����B��w�O��N��_���=�|����1��˪7x���#���-��L����c�����n?��ߟ}�:��XYMF�D,�?{��OMZJ� �������C�(k��<����)!��3����D��1��B��!m�1-+�l�F<}񀮎��^�c:�W/��w�ȉ68z"'��������b��X�9+�о$jeׂCl���%�&�)�J����-Bʺa�=�����Y̴w�L^�u�C��C�������_�����yU�H����U�<"V�;a&�v�!	�ip$T�c���7�ë�CT��c�������̂��8�vN�qB���JԒ��E��3`��b�	�Xec����B�,�Zݨ5�%��
��Jk��{������,�b�Ɩ�m�B�	MS(��2Ia��5Ɖ��D���a"��X�@&��&l- ��a�m��_K�2*\W5� �6��f0 \la2�`�4�+-U<�1�u!o��76� ��O��@�����)U��:
�hA�4����E㗹I�}v.M��DO�넼�J%Bni-�X%R�[�ϐgo��R��E�b�VTI[��,L��m��a��<���=-��Lڷ(k�l��q��]�� )z��0"� 6و�yvXZ�@� ��+wtǉ.8������վ��z�?~���P#jBm�0�:%�M����cV�ϮO�?f��ތ8ܛ��ߧ��׉��ӄh|;�n���K#�q�w(�+ ��`e��g{b\��G�Z�hA�/�C�[�F�k�(%���b��f����1��h�c�C�����"�"A޷}��|\��������S������r�TT�L�Z0
�p�XÙ�OQ�a$ȳV����	$�RM�::k��L��M��(S�V��S�*�	t�	J�\eI�*u�IT|�H�	a-�]іK,��F�D̟���v��/����	t^;Pw֚��-���"!�����imM�4p�7��֚���4rF��l��pT��n���ވ ����oG7���C���V���xy#�? 1�!���A]w��#�/ia�H�]��FrD-$ %  ��(��F����KC95 [��F��L��4��q�y9�����|�%�9A��Z�uj;��ﰒ��}_���ZO�5����䱱{�.(��μ��U�3n*�p\��ޑ8A������q������L��8۴�����8R�'�"ڗ��
Z�xiwj��Wb_v){��i�+���`e�k�]����{�����Ӱ 8
Ǵ�<�1.��6K�����r"1���[��c]ϻ-u�gi���Ke�����`A��zI85p�4j�.z�$8�U��NB�;�ڞ��`NP��H�}K��DM���wД_���(����v¦h?4�l��I�U\���9�+/A��l*O���a�+NB��<�-�B��+H��p1�ka�f$���y��l�5,	�p�_�kA�l������`ٚ ��*�� �~�ut�@v\�M~�����
ڏ�%��e����r�ќ��%�#�+:	���,&���q�*��VB;.�ˑ�^��:c�~8p|(Μ��+:�q�];�c��3�KD6̂4� ��Q�d$b2:!ȭ6|�q����A(m�Y��H
.~���~���?����ϪJ��]6Ue�	A�� ��yz�L�������u�}��6�U�[��O^3����c
����oO	M���X�,�!��4��^�}�k�X�޿{�*b�ߞ��^�[�(���;����g�	��L��щ��h�f�G!�U;��DV�/���a:#��G�ǬJ�q��u��8����������CgW��_�f'B�U�h��S�_��B��a����f��l��.ñ��7x����y�{�X�'�	��5��1S��ϟ�knc�Nf+6��_���1:$�3	����H�o�G�8Ep=^S����<�]}�tuy��G�c�Bra�SU�y��N�됫uB���^�
¨��F�o�+�U�L� ��� =[vAj$�N�͏$��� �&"�wK+DX|��6Acg�P��<�
K���1���i�"m�REZ��<�SE�Y�=B{�4��M
����"�[F��4z��
yL�g��Mw��V�6��������yx��
��P�2�
�kХ��u�WS�pkv2~���m���S���e�Ǭ]��b-A
?���3C���Fe[��:<B�uTQ�xk��U��P"H*A�N�����(t�x��"D�z���aN���})s®r'k�K=|�m�@�8<?�!�o�����8<\� �V��ɺL<ߔ�[��f{&��-��+���	Z>��ǚ��hTi��íP}����Cm�v�=�
o����Th�';K�ǆb��(�M����q8߯uÎ�X���=1���&ѱ�
���¦��O��X;�l�P�U�xG|3��5>\�
�0w6�B4w�@����։��&�(�E��J5���HPk��� ^�B,\}��b	E2��3O�����B	�����5
d�H�Y I.@C��Z	2�r�X�PC����B���Q��4'Gĸ���Ⱦ3�Tw{~�l�d_��uL}����qXJ�D�Y�8��N����W^17C߬Rtj��f)�h���&�%(��G��T�G��2�mh{��t���ٹ�K�z�����㚵��m0�yF�axQ)&���*��V�ǌ�=1�s/�����5��`���9�&��iÆ������l�LlY�g/ź���v�,2c[u��Yq��%v���{y���3J�J8/��$�Δ:b9͗Hl������%��e]��.��r�9���-�P��'�nX�ܫ����)�'.;ろ.�q�ړ�KF�Ѹ�x��я �gt�n�i�'������2|E���qYl�C�1�`e�<^�
?L����Ѽa�UN�sp�2��@�W8`���5�8���ki�����lp@d�����]\��6����	I !��@܅�$HpwwwwwwiK�R�E��w݅b�׷������9�s���Y��G�؞���e--��YC�8�!1����e_I3���c����.�(�L��}����N��h�K@���SӫZ��Y�{�ֽ�� �i�7������;���X �S��Ŭ����x�����Ӑw����ͯ����r�^�����mz����4�&��"=nӶ��Z��4���uJ��� ϛ��k�6��e�JW�Yέ�;-�' �D��k�|��4ݒ�;��e��oc���}n`����s������է�.;�m�A�)�=�M���F�3���q��M��Qk�HO-�CF-!��E�١�i}��Kf�p��6��Lix�(O����3������4n�Z��T��g���k_~��[@�?���������a�_����~z0���N⻟��˯wD=��ү��#�O�����/�O����Vp����u}�~�~��7����'{�==��VQ|�O�Z��G~�,/��K׿��Ug�(�KQ��q�*�5�H���Q�Gn�pW95Mt�7���z�&o������0
]��o�<u�{Bɷnmg��1�UFvS:��E��	��YG@i����Bѽ�P. w=����{�Q؃��w��}Չ����{�л��޿N�jg����ꫯ����M��vR��ں��o���W/@���I�ᾼ���o�V���el�y���!1ǤLy蝵&[U�gվ�Fܾ�٘��cc��@^��;��tncJ��OWC[�F���/a�&��Fm0��!]H��H@Z�~U�S� ���H-n4�h���>z��V�~�cmd𗨚�VQiZ���T��o�ExP�}E2�I�}�)\sRzP�T�f�S
S�E5�j1Ԉ6٦F�*gƭ�y�۪Q�-��d��+=�9^ՓC�'3)4�V�-�k�m�Bz��%�uM��(v��6ԊIƼ4��-��+��5-���$[��!�m#��jtTS���3�S}�4�3�{33�3���yh��>h�z�9���nE��-͡v���ef��J���͕��8<B�ק%���d�_��o�:�����ۑ
�H)-�g��9�K��F/xe �1��ҷ��>��`|:>��τ/E��_��_��S��e��yOd�����N�t&���&��o����Gs��`~:��W���lCW�^���ى\����11����@֕ٳ�ș�n�G�n�VkT}m�=8ʻ�icM���N�k����|xM�sq�LHbl�5�&:t34azl�*{R��C�3EbH��P.Ϲ�ʊj*��)71��Ι���;�1�ٛf�ٹi��ځ�~�J�gdH �]�͘�`���0�C:��H��IY�IHbPp3�
�ק7u�Y��dѫ������/-b���rX#൴����H�_2;��%5L�(`^V
��aV��,�0����0e�d&��ډ�Y>d,��f{���9�g�L���y����g�-���<3	������i<7w�����K��h���܌EZmܝUxq��;v<����<�t�/]ˋ�7��ڝ��d�6�,����+��<�7l�pE-',�eh�E�P5y�M-�!�~G׎;nJ.<��Ψ���U�V�k���Fn�4�� �%3Gn��F�Ա�-}{^@|]��C�5��.��m�4|[�A~��z^�uo���Ɩ�=������� �+b��cf��������j�~޲����gsxG�X�Iz��$F���qN�]3q���E5D�N��z�Z��6-�w^ OŴ��o�~s+��e�Ϊ�l�� �p����"�����t*݀}�K��|�6�ަm��^Ǽ�'6
�5�% �:����N��['p��9}?Ǹ���izW�L�o�X� �>���q�#���]�/p���b�Ғo̼��Z_��7�A�f��"/c��e����S�7p�&�C��o�x{������>w��-ج���u�H���?�g��8ם©�.Mg��<�M�\�Oc[u ��형lƼ`yk1�Z�e��a�qM��m�,�;/�+sAٳ��<��NC�o"0����b:%6Ӌ�qCI�FY��TW����/��դF�P�.�������WVr;�0hP{��s�N	�_�;��/���^?~y��O������p�h�q<|4��~o�_���k���K<x�3
RV�A�w�.����m�
O�?��o�o��^���w���=xе^��_�W��\����<r-�yMx��b�����xw��5���"�2J��A��Ѵ�ї��jR��c��SϿiM�
�T[��<�E>��]�lXFN]ay��SR�w�r\�
�혍cZ�]��̫�=?_������[�MN��F���E��E�T�Yҽ��wM��D�Xk�85��K��Nj���;��՟N��g���z·�����o�KZMot�a�>��̢���<yN�Yڲ�?U��-��'���;�h��T<�$Qn�6�HA\(@S�oM��+9n>J����T�}5"�3 ���rbcP�T�u�`i�#���!���1h�Gfj��A�
�D�%��)�oJԲj�zZT���i�"KՈ�ʹ(y굥�(�	������{tZ�M��Մ��N��-z�l30��j��V�_ ��{^�ʱ�^�;����%�4�)8�dl���5R�aCS�%�=ykY:/Oo��	<7"�������)v�9��H��\���F�*d��8[;��*PcA��!]<�h2el{3�g�q�3��\�í	~�� �O���͎4�ٓ�*��X-w��νK<�ڗ?���M��7�x	��'0��4��/Ⱦ�u�/���+y��)����5?t��R,����6If�*w�d��b\���-�G;$��y"����v9n�"i��Z�\ş_���{���|3_>Ӄ/N4����wT���Bn-����N�<6����(����iI}�)�-q|�?@�6Ƹ�kږyI�|��+�(�5�/���U�,��Bw���,���������P/��N�`eǴ��:���ʖ)��N�f��?#��[]ˎ�*f��Ȣ�tf�v�p�o����m�2)sVT����z�@���E��q ����C@l|rg7�eˌ�L4�AUݙ9x4Ų�;p�%=�Sn��6��e��/���Ɗ�
d���G��X�pv4p����`�������0����Ÿ�cZ��܂J����|�A�j����L��cZ�f&�����}ӫY�O�ه���L�mba�F�Uճ����y�������K�?����9յ��9��Z͙�rNg�r6����U�i�d��|��0{*�q�ރ��m�ѷ�u.H]��H�R�uwY׾������A=�BE�Jy��SkBU�^6�Xt�e=9�C�L��Ұ���]0;/F�y).��ߪ�O5��𔿾K|wں�'7�^(��c�1_�k�<U��
yZsmP�@>8�m*0g$�hSqu��1��qQז�z��{"�9i͵*��	I�9�����lH���5��?|"9����en^U�$:w9f�/���A���L���:M�3�s��D���զ����,�ɲ�@�No���o�>A�ϻ��P��o�4�#l����7q�.C�Ī׍���W�Į�
���p(?�S��"gq.;�k�	�
��½�(����K��g/�F`�>}>^]���uY�pϜ�_�L��F�>�讓hW8���I�L!>o
	��\5���)��O �h"]�P\:�sh.�F�ڱ��BUaj��0�a
k�2�b�J�0�~0�y5��1���3�R�xA���`��8���(�]��ە)��I�$%��"�������2~���6���Ume����
�\���b\�-���|��l^�p+���F��O��ص���=Y�M���;(&h�������{ksU���v�_O����	�*Q@���7��W��~^ħ�4��kͲv�8g��V�Kj�y�R&Dw�O�QT�Q[O��a���R����U�0OG;��o���<�̩��D{�}���K"��#���$����k�4<�*4���R&X����k��,#��dv]x�ճS����Z?��!O��u���E�w��'������o�s�������J��%򙫯�QӌIH�1q��Xĥ`%��j씨Z<��%���l�B�Y�&]w��4/�vvdX�QddE^[#�E1�����6�L)�S�ꛗ�!��մ���j�B�
Nuq&?8���!t	���1���Zۑ`�@��+�&fD�mdD��	q��36&LW�жm	�Q�%D�Nkꕹ�$�-s^KՆytv�5c��?�v��a������e̩�}K6뚰հ�6�5Ӝ���9k�Y����v���v�D�h铷���@�L�)���˔Q�.����+�xiZ$צ��ؠzG�i}��HR[[����=52��@UQ$T_�pG{2|������������� ��ʝ�|�0��V'���l�<�+@S���N3�6�/7�?�M��f�������
�-��h�Ծ��q5����o�X�$y��������yto�o���m�qD>H%{��)�[d���'r@r�A���l���w�a�����v�_ã�ūc��K���B>8ۛ����罽U|����Wd���xnL���AĊJ&tr�6�� }-���T��G��=#�j].���ա|���C��&���807>�ٝ+(w��؂fk��y33�#<��c��Đh���2"(�A��l(��+a\t{fwJgJ\"C#�����Z払:1.��Q)��Icjb.����ψ�d&'f2�C:�b�(�&;<��������"��B���_���	LO�eJb:�:�1_dN|� fc�"�߫��X�ѕEb�-�Jb�|��r��E71�b]|��	��ɑ`7g�}�%ײ8,�	^A�9��+FD�|s�66��Z�ii����7� �Ԓv���Z�S)�m_F;y��'�e^����3���1l��b�w[e�������+�-�������|��;�[�qY����x�̙��� e���m�WDn��qSk��Z䶩�6W봐f��\��憡7��4��
U
!�[��e��k&.�l��K��jV1r�	l��tu��2�s|"��ہ[��j�}��Kx���=�=w��:q�,�u\dIC߂[b�nd�#�Q��b���V��u��PgJ.�9�Z��=$�[Ӗs}�	��(�Q�҆��.�@��x6<�]�װ�y׾o�&����ml{��m��xy]��3�%�{�ǭ��z]���.5��S�,����Wv����x�<�k�	��8��ıx��7�Y���m�T��ʣ���D��'�bk�Rw�Ժ}���"��r�e^�Ud3�[��c����﵃ꁻ��ʦE��ZJ���2v�o������I�W3o�F�,�Ò%{�7o;3gld��u,���cW�u�Rv�^̾��90uG����������fq~�\��|ǐ�����rz�\�9�s����<;s&GGgNZ*K��sn�\Ig>{g-�[�,�l���)���y��EuJ��~L����~��F�۟���o�������IY��SE���.�b�~8��7�3cu3�~��P(5��w�{�)[j�>��������A�����7^O��S��Uw��ד��S��O�5�Bui�;U�>���M���x��{�L��kn9Y�w%��6��b�����w8qM���4�G/F,Z�����Z!x��N��:���	�Ƚ����OY�i]�T��-�^S"�v(��^Mg�n?j;��{B]��)�5�:v-����"܋��u�d�����o
��>�Ek
m�:%O��֗�"n]ւf�y���Ysl�De���4��[�U�c�����_9r�&]���ƿf1)ĵ��S0���=#G>�j�Kj�Z�{z��gOO
l=;7mT���Y��]M�(��m�O��yVZ�%�BEUk�/SS��鑕���
��kk�TG/v&�s�g_n���c4�WJ>;��_�������TV���ˏ���o�����D�X���Wo9{�M��Y���2QbK��af'j���0�����]~�@�H7�[yqP��:Vy*B�9[D��[k`�I,oy[-��
�=�_OA�bg�ֳ�iý��`�R��F�X��M�/��m�C7]T��
>^���)��89�]=C��lq���F��ii���
��j5�t��ץ��)�:�3=ۉ]������ɉ���3������<8_��k��A�������@��%S����5�m#��Y߮�`�։չ�G�s���۟{yxO�����������{�r����-����x��w������S@�O�?�I=.��V=Zϣ�E6k���@��R0m���'i�.����P��6�u��/?�Ǉw&��呼}q�>ן������M||��O�v������W��p}n:όnϞ^�,���G��;�`#ϰ�<����4�=�� �xt�'��$31��Z��<[O�$/�afI���%�X;S��M���֞d��.�q���H��'eE��.>Ի�ShfC��=�F��j�^!������;�n."N4l���Q+�N���m[򀓉v�m���*�܄F{7�;xk�9���Qn>�k*P��#����h_�8��>��p�c��;�|�A��n�m�6�Ӻ;�XQ�����P&2��[Kw��?Đ��0&�ʘP�6��Ǝf���rpb��?cD&K�3�Zd��(?���1S����>�ށ,c~@����¤�8v�+���������\�o񦡭�d�bԾ`�j��dY�L�U��ۺk�[���|cO��F2H��'��9G�%�v˰e��μ*���Q����We%��~���M9���{�@�LΥ~�ѓ�������}2�>y
�ƈb�:���c��m�yO���u,���R��2��DA�ۺ"mlyS�zU��.���␅W3��h�������PHMr�2Ɛڰ��WU�()(�DN���%3%���e�s	I�H����4���0�1�3�!�Ci�FQ�At�j&6����^���&3�'y�}�,A��i��5��s�>��,b��EL�Dd�Ǵ��q˘* �dք�̙�L m1Kf�d�,���3j:���f��e�����S��h�R�M^ʼ��Y>a!��.f��ٌ6��P֋���.�Ǚ�z�
 ��n�l��������:���q0���%x�|0GE�.��Ѯ=9����΍O��Tz=SX��W?vt���)l6�mS0�� }���`je)��UӐ�E������n�Z�{��ٗ����F��[Ž?
����K����_���g}Y}�'��+	�Kg�����ٗ�����_�A��ڹy�O�wS#<�x�λ|�ɷ<P}�$ŧ]�<��_L���j [j![�n�i\"��Ӄ�l��9c7\6���a��k����q�sϩ�ZR]��j�S��W�WH���l?u�o~��uy$I����S�����<���^��������gJ��j
��?s�f!sV�R�{\;t�!���R��j��U!�W܇��b\z��<��x_��C���Ç~r%r�Ч�i���B�ǲ�vU�d}�Km]�w�זQ�B��.5�R��j�kR��UZ&�5~�ݎ��*���E'�V�Il
��S��N�[(�xAe��t�cC/*�H�iq���G �S_GG���E�YQ* ���e�"�ŕ$��IH)�
41�8��:�W>�c�[8h!���
D��^�^�h�����~���O������|t�8w��<d�γ�>�wa���>G���k�b�*9`��kN�zp�ɛ�>a�%�q(���F��Y�c`N'C�z�	��Pg�A�V���
�)�$��?C���׮�&ow�Q��kV��C��$�MRXo��A��I&�p  ��IDATF���ҡ�G�u=��ao�[�ʕ��\ɖ�@Rd�`�/�Z�����6z�9����C�$G�{��9�g����L��E)|�����{��?�7���_L����m�/d����+��7�j���P���ot�m��]x[���~���Gl�}��1�%3�m�UM����m/��Y ~����.w����-� ��[���QD@��r���j�.�|��W��������|u:_�:��^��W�����\_>>уώ��s�Ot��M%�Y���93�=����F��r�� _��qb����� �{'jycI�J}��p��oZ�i+`Ն��h�W�T3;���L�*ez�j&g�17��9��L�ԙ�Y���)eqQ�YYV���)��R��(�beQ�ִ��XW�3';�%�y�+.������gjq�(�b*�h�VImi>�%y���`S�j~md���d������-�bUq���C�M��C��r���ZN���q��  @߿ۻ�bp�ni�����ܽ��5u�������<'���=p�g?���Q�90j���gk���0�S��sn�H�����C8�k �{���\6�+�e>z4/����	3�1v:�FL���sx}�t^�8�;Sf�/�����سlL��s*LX[{^�o�K�vK��S5m�i�~Ks�rp�w�k���Ut	x��9F5��2`{y���CW^�w�T�e�m=;Yo���B�[��UI�I����y*}0��~r���PAޛR~�l#c��۴�7�db����y(���c0��s8o�E��{8�x�{0o��s0�:��Y�r��Ik2�a���=�R����c��MN�T8��ܷ+�Qӛj�32��a���i�<�� �NX۶��97�P�"�nҁ��y�����t�xd�-(�9A94x���#e}������'�+�L�(:ƒ�KG1��O�"5 T���I�����|�P�����������M^d�i�ڻ���Az@0ib$z��+��o`E���r'�-���ѧ��)�����A�������Ͼp1��"����*s/֚��%�-��lpm��7;F��:�M��"����5�f���6>�o`g��L�����S�6s1�q��iZ�|���陛M~b(��>�\�Ƴ�2y�|>���/�)��_��Q���j1|{��O�9{���t&�&�4|�VЩ��3/^���j8�ZR��T�<�'<��M*����`��_{�_Q~��'��ը��������)�iiS�����G���}*�m��r�x�9�q�(�3���J\:W`���A^���b�N��i��:J��k�x��~S����܎�����ο/�G���ן~�g�������ΤU�p(�w�����ôN�Ǟ�`��xB���*D��޸���VR�WY�5C���������Q�&���J�Lݹ̟ܷ��.���o�Bu�rŏi�u�Mݐ&�~���Տ(�o�ժB�=�3?TaQT�P�:���q_�k�_�`��D�@�]�Ÿe�`������K��>5��y$�ܣ/�z_�Ǆ����q񦭽�6����ggڛ����K����MȲ%*�S�LN#��{��J��71�!�3�/� ]3��e|[�K>]�]`d��9m۲�@�պ�lP���T65WM��tԲ%�L�'il���ܜ��^�'+�m�t��b%�a�NI���=�<���J�\�=�\�V�o#2u�K��	P��jM��/���۬o�v�f��\���a�����L]��*h͵�QRp�k�:6��7�	�2�@�fsF����\��QǭY�46Tt����j���\���Zw==�����uaF,,��Đ�\�ϛ���|sg~�_ɽ�M��� a��ܽ6�o���W3�kX��,��O+%�����I���=ަ՞�"0��õ<x�Q��"��
��Q��H�7�o�����k����We�}�7�n,��+����<>7��'��롁�=ԟ_�5���|���ow���}}��� ~8��o�������ό�3cxt~2\��nχ�s����|{q�^�7���ŝ1|tk�_���{���*���8���g��7���2�.���I	��Ĵgj�	�ӡ����� >XٕwWw�}��zS�6���5�k��$O��_X���fV	�	�-�Z���F�t�ǲ�ZVwcsq��Y[T/ۺ�A��M5���8��=��F��q��c{��g��������lm�����l�9��'0�����h��Ç3��@���ɳ9;{9wn���eܘ����W���\���[�6���]��f/o���K��ss�nm�ǋ[�s�&��[�|Ic���l����3�ʱ��<v.�&,���\�6��d�-\͝�+�!�\����3���야5w�&�����kys�F16����-��p-o�Y�kӗ���M�1e�&��§�����g���̍�4o;�j��ը,NX]�1皑��+�%.�W�[B����JTөj2U}��xZs�]����i��oUh�&ΚϼF.�
�\��ח�T��?--�9h��Z��U�����]�����л*e�'�?y�qJ�o�l�Y���	�d��q�'�#�����e�gC����xh<'�c9"�tH��_�#���� ��{M`抡���yK7���{(������1\��}�9�.i8q�!������FO[7-���Ȃd)�&Z���>���8g�E�.�t�xD:\#H�	4u&�֛ s'�M��:�ƕP[W�m�5��6P� +�G�>_�#^��q�x�Z�-Ƶ��9��F8`�'e���ݖ�x�[�ad����&^R���8�-��N��]�G��,�����vk�Q[)m�8%��[���N��(>n��So���N_6Yx�E@n��{�|�! �d������,�����+���QsY<j&�FOe���LnBNH��,5�Q݋��I~gF���8ёw�O��O:��/���#�_��ӣ�\~c�'����D<s��-(&P�>�b�N\�'_|/*\�������?��婊��iR �����?�|�V6��[���?��4��1JZΣxF.W��<�U�X����2r�	B�P��������Y�sV�V��޵�9Z�����ߏ��*��J��׋�	׵���(�O�����&���[(룷op��"殩$�>��:)�W�p�\%��+��~���W�0#���tL��B�C�x��R\����.�KP��4,X�sw>�<9��q_hM�Pyt��p��(�C�c٧�4�~y��}�zh5�*�{�����V��*y��> y�����âgp��NB.Ɲ
��S5ynB�b5;'�XTD�޽h_[O��C�1c1%������C['<GW��q�s��@^����褛ؐf�M��Nm�[���ĚS�H��t�\"�'�`��!�mL[]�<C���E:GW�y��D����"��6�1�bҮoc̪��Z��ݲ�� �CsvIA���n��"�lP�ɾۨH�iۆ�������̆qR�(g�
���l�zB����urʹ��<�V�V����	ص,��zf�����l24i����y�����O�e��râ^�1��D�ɛ�f��e�|������qmR47��3'كh9F�P�J�;�P#���іm��\��5�~���_OVq�\�/5\���ypk<ޚ΃��k��x,p��T���]�c5��w�,���zm�ý/�q��9<���>_��gq������`~{a w :ݛ�D�i��������ۋ�4��+xnt!��������&Q6u���`_m$�+C�Q� �V���6����(fo��/�C��쮑yc<�������\�%�6��kKJ���������c}x�l?�;ۓ��6������x9�*��S�|�LO>=�̻����l^�ڞý�Y��Pi/0=���,(�U��kKG�ޘ�sC"��L��մ�"�+���Ň�N���q��H/sgz�A��΃����|��Cm�$�}l��g���`��`�93P���� '?��z����r	`��?���K��X��]q��բG8�8�&�*����p�Cc靘˰�"%�1 �};t�9�3CR��]���*M��W�/����<2c������{?�](sf�G���Y��Ҡ,	KbNTGf��gqhK�۳�G���X؁����%A�,�Ă�d����"2��Q���HbYp�������4M�E�5�3�C35������J�}��p�mK?�KzV��d��+�
䩹����5�;�9��j}ݮK�� 廬<�Q����[�S���IZ����
�T��j�U1p�)�S�{w=�����x�[�-������E��މ�&^���)��K����9���Ԟf1�ٸ1X�� �Z���ދ���,�	�@pW�\4o��w�L��T@�΋����܍=�����K��4�I9����W���"��+ƥ!qf��ۚcbD��)��ݹ* t�؃;L�	��k�/�,��8�ޅ8��8Cb��U�ǣ�l|Z��|�3��$V�#:�ii'Fn;1ңڈȾ�Rf��q"�|����D���ߒ^���R6G?���r�9a���֊���6�<���pN�����1��2�g��61�:rZ�X=5pe��#��]٧����ed������<��r����1�
8*��9+X3v��d;�����ޅz3������Ht���k�s�V
|���d��7���Y=�\��A@N6�i;Mx���WN@~%��/k���k����.evK����<Q��ä��������Mc�N�D��4������:F��+�5J�h<�Fw���������	,�M@I7�
k��U.R�s����h�"m�E`i	��$�n�}�iW]I�c���m�#9����S�'�M�;�_.@��?����Y�yɕ]��J�C}-�#��t<�o~�ý�y��LJE��5Q�U�SN��Kpk�#���u���;�Os������ 56�G?���B�#b�2��%j��4y:Oܱh�(X�=H���ӠQ�o����?�8M���e��P��z�pO�ه?þ�S8i	6YU���gVa�^�KV�V5�۵�0���Rb�kH��ABe7zϜO���Eơ#���/.�:8b#�jgG���V6thIjk@��#�p2��H��M$������!�!Q��5v���ڐ���9��.3� �!�T�=S�n���,i��R��R�-�tY%�V	�-��|�Xp��ڰYO P@q�l��F_B���]$i/ik�F9�.�g���OO�F6%<Q��P
#_I�AGO�9f��+{ĚS�xZh3�2E����o-������k��c���=O���̴ѵ
��
����ī���rO�����Qz�LN��|���N�m��hHm��yv�o/����i�|��_�5s��~�5n��)P��)<�t>�Zģ���/+$o�=�������/�I&Y �̈́�S��(85���{���&�Z[�KKxef/��ĥax�<gz�p�)F�U��,L�`a�?��{2�����ĸ30~�������φJ;*�l)�߅>����H��ͩ����ǎ�_��5=����0wƴ�`R/f���k�b9�7���xiV!n.��5�t��oNW�<�O�4��3}y_��������3�'%r�w{ƥ��o��@C����'k2�t]{���Q`;�	�Sd嬶���(`+����ܦ�� �`j�(c�1�Ą>�CA�)F�#c�0�POĀ�z��ۜђWF�a2@��k�QvJ���'
n���(WV	���J>����]���-�ƖX�9�d���+��K�{�7�%�{��[~�i�/O�����x�5�J���7�����'�,r�a����.��`��{>�X;��L��3��49h��1[Q�"��Ea
��UrH~�q� �1�RU��ܡ��cN�})y�ҝ3n�2u�䬬�h��%U���W<��g�R/�q亁�y
��	�T�1�O�wC@J���x��J4����ᓚ�����	t��iXA��+�S�Ts�۶�\0�8��=ѓ�����/\K����^tr"�=�S'ҕ1R-�ȴs�~gX{�a�M��w;{[:��.�pa�{��b����-TMǯI���|8i��IKy��<k����-s��V���Y��K�����)av�$�X�[���y ���ʳ���X�	�g��EFb�[,�w��)�Gʥ��& �(e��S]/� Ц�I��V�4K��G@�ii#W�W�[���Fv�Է��@|���'p5@׆�z���ױ�o��/$�A�y��M��`��1�P���qV�M��!�|[NʻQp�EεI_t�|'G�8.�8lf�KA���R�☉��K�ziQ���{�B�ȉ�&N�ZʮEk�4y.�'�a�ą���MuR&�j*�>�;kS(J��4Ӑ�#�9r0�W����;u�;]Ϝ�M�� �:ˌ4l� �(�.Q�SzW�;�W�]k�8o|�`A��y��0�/�C����|��g|��_���yOOA�y��O���>-Z:�4��4yt�w~�����Ѿi&>�#�)l� ϧ�Z�<5W5w�FOݷo^-Qݚi��D@i>!�](��̺�����-�{
���<z��4y����=�����{�"��O%���.��+.�hx�p��L��J`�]������8��'c�R,�T�mj���j
z����| �j�P1y1s����w?�����"���Z��:S��ةfW%
�Ժ?���X�@�C!{�4���)T�(њf��ӯq���]z��n�Љ�E_,}O�N��
�;��ݥ�ȪF"�눪�%������T��D��Q���ozg<gt�<1rq���Q�a�bYښ��m&��-�V"��;;�oh�53�fP/���V���F18)��b�B�I� ��\c�&hM�B`��1�LMYfd��mX`��3V��Lπ5F���L��"KkEyn�k��k�r�Y"� 
 n�7b��s��;#@�,�m�!�kcE�\��5��WNl�%�h�~�]�=���SA���ޓ���!o�gGk�����yEh}�Tmc+�m��V�}�@AOs��L'n�(��ռ8-��S�ya\G&���Ū��H��uQv,*��ٱ�|�!�ߏf���\�8ߓ?_���c���P������[�����Җ��ϖ�ǻs�{s
��O��G����|��ﯯ���<.�N���t^�ȑ�Hv��� ��]�X����tg��90*܆!�����9�v�Z���Δ}R�Dl�H�5%�L,pS#�s��!�<�"�&���x��ij�ŖU�8|�41&��T�q��,E̍�(�d�X�koC���nVtsP
r`l�S��pe���Κ<>�UƧ���x�V��ə&>;Q�ǻKxki6�%���=}���a����>[_��:��X��M`}a(�a`�$#+���w2PD�Қ 2Fd����"�a���'�&�L�!2K����Et'yo��ђO�����m,���G׉�c�D���&��&H��)��=P�S}]�d�����}��*�(qU��m[֩'��JC�sO�����"y�f��4�X�rH�D�H[�?��	�_�k���9"��8<&���,��G�>���G�أ���9)rZ��wA�WrQ}�"O��"F���y�;/�_�6U�R���A�h{򌬹%�� ��Z!�A�(ٖ��t� ��N��j�D��S�3�ur5��@���ƥ���89~*���8/z`�ED�c�u,P��@;C[R���lɐ򳃱����zw�w��څHs�+B�����4rb�s8/��sS�掩o��
X��@���Y�p�ʗ6<c�Y� ^�ㅀD�{PnkC��a�$����P��<�WLy�6�\#���O��QR��;a�D����<Y���6��y��=�nA�pU��%�������>����k�E���`� �W)kd�C���jռ|�=�Cn�Yc��Yw�=�g]�9g���f�s��Y��Rn����p�Wn7�~:���~8����vJ��cb�4{�Y�\g�y��ғuFά���DIM������x[&�g���kICzm���nŌ�Osi$�Y��W83qJ��1na��J.�y�V�t��å���F��H>�/�ƽ�ׂ*:�ʜ]��Q F���?C�j�������4��"_�G�V(��
��JC.M��-P�ۻ��u�$MC�*�O`�P<�ip�
xO��d�ߍ���w�k�,��J3n,�����>���?O�_��ׅ�=���?���������q�zjG�%���:<J��[Ƅ��<w'����k�1zq<Y~��f�ݬ��S/�!%��r\�p,l��L���7٣�3a����1�߽���oOE\SCAT�Ai�)Ώ�Ab��?�	�ɢ�o��^�^K߻�e.)=�����Ab����{|��N��������}<N�՘��c���[^%vIyx�� �ܮ���M��VҮ��.�FR?c.�g. �{Ol������?:..�����䤅s�20� ��cblIv� ��Nk�R۔�`)\}���M�(���S%�z��`Ж��p��5�i!s[F�3�%F6���o��S�-�k���Ź&�,7�a�Xd*r��r�J�@�[)�`��� �@��%�DI,��gQ[=���X!�@��	X))�j���\��ֹ�L ��̘d�����l7wf�(����ZS��o�4Us��!O�/ț�����l�)���jSk*W���Tǯ�t��uU����9�ʺ��V̥a\���	��T�:����X{f��܅����dg.��.���jxq\ɣ�Cx�|__RN}�ޙ�O��z�f����|��.h�홍\Z���x��5�22��Q���Ӧ �yr����r��9�^������'�� =<�5�68�zmq���(�F*�*v��(ly�J�����(��J��D#�����m�[�%���͍z/ʯ���.vF&8�Zj#��̈q�"N ,���LGc�=Lb��<΍J��%�|����w��ա">=X�WGj�|g�.����Df�82�S�e��y}U7V$���Pn-ObG�XF{[3Y��}s��M�k��o��vr�%����Ƌ�2��%�ۨZiC�Kޘ��@�I:F��tyNs��oh�\}�ѲH�Z$F�ܶ�̔oa����p��r{Wƈ���� �2W\ڋ��0*�����gj.���*y�]�o1&�\�Z�,�1��c���̣书����e�#��ݴ���y�����l���,��S�2��K�w˶V�%�CD�o�f�����߇d�C����Q�Ӳ��V9�c��m��A
�T|Z%/�[q����=/[r�Ȓ[���H�V�k���8j5pʵ�)nʱ�\�WP������Fݪѳzj���Vc�@NI��Zw�/�
K���V{�F��f�ϼ�s5:���W��ϰa�v68δ5똹h���*Ǧ,��9�R9���'R�5Ƚv��12�V���V�4HY���t��ֺĴ�����'�:�LH:��-�P^��⦝ϙ:���3�g���zqB����sV<��<goJ���]��C=�ܕ�v�\1��u�(N����Ȗ�?��6�эt�A.�	n�51^�	�]q
ⲽ?�����0��x󼬻(�w�%�]C����e��+N!�\u�e�0I+�K�a\p开�)���r�Zlq5h�U�m��U�*�{�`��+?.[��3<ڎ9���	�fIx�c�X�.����l������gQd6'��1�-f.����gzP{��$���Ct�7K��9�q���g/a�l���#��j�����ڞԥe�#/��#��\�Ca�(¢m��A���D�v�7�a�Pa�����������5	���\�����rB��!������%>�M�L���6�S�B+X==�m|��~����?@�:^������������+Q�hi
O��<�y�|�w^!�q"v=p/�}v
ꔴB�c��SV!E��7Y��Ϊo^gƍæ�s8�i���D.�yZE�cU������՛�X�y%����4�h�"�E�q��b~��̿����6+���X��g�]��� {�P���3��.ƶ��\E�#	(N��1lx� ����������|���ɵ������& '̮MZS����?�]��ب�]ܸ'�j��$������W^��դ��KZV��Z;��b-d�W�b�h_�LB]3�$6���TN�N��9���FHa5N)�1�K@?8'���󕹏�*҄(-5�P)�HO�(<U���{)��q�{l�V��gfN��NwQ܍��Y�E��B}�C 3"S�����'�B����2+2����)cE|:�"���D�k�PZ!���D
�u��1u�bȪ��J�*�[!Jn�@�"���r}{D���h}1��"R��p�{K�7e�";���.Jf������F� 5�V�j�՚rE��ں�F��w��@eo���0�v�2�a�<'y�Yi �' Y#033�]��w����`�M�������I�i�g^�7;��cG��I��Ce�{���g���� 89N���=��xp�'�h�e%\�����m��j�f�z1=ڏ�A.ԹZR�bA��)����#H������Mպ���ij��� �Q[�=-ʈ�<W�^G��&���ȻU84x�k۶-:��uڪmƲ���,�6}�6-�w����>�>:F���.:�m� ��?@�l_�Wi���j�{U�Vw�=?[s¬��hiA{j<-n�����+:��\��څ�/�}ռ���k�r��-�	�Ӓ\879��ӹ�"���;��9���V�06f��)ST��̗��D-O���j�T-��Vț,ۧ��"�p$�D5�Ċqf����M��1C��B�9���m�Z�i�m�)�.�r`�11�����-�&L@�B��oiK����rn�/AD��T��0�)Q�T�H�H�H�H?9�DICu!8`d'�f(b��q��U� P�E����eWS�D5w���&{d�=���5��A��<U��j��
�=�c���>wZ�;�u
�^00�b�*y^Ҹ(��e�SN�9{
��{i��k����yp7��۔њ<e�W]5y�@�.5�U�ow� ;m���S�sH^H�c���n�|ә���(�b��Y<s�:Ͽ�
�^���or~�$�Ʀ��;���8$`q,(�3	��`` �B�9���(��2�Ιb�+���Hp�"�Ԟ|3;�8�p9�o����@n�Q����y{N�6�ᰀ�Qg�7��9�0��ky'���re��f�\�5`zQ��qu֮D�;&P��Wo��6��+��ܴ���h>����T��ZF�aV�SW.	 _1���<�C��,�"{����h��y#W-jɳ��9sZ���\�<�1ii�o��n�;)�v�X�������z�⌙<3}���žc8?n*{�{�> �MA��=��f-�X���'��ޗS2xf�LN����v�Y����<N�Ċ�L��t�Ȝ�l����3��z�,֎���A��<�g5��i�΀�z��pt@O�Ws�]V��T7���2�u�v`%�K�P�Ip���v&H�.�����n����QT��Ih���'����;��0��T�U���_>�'p����� 
�Z�?�����W����I]��k|�G��v���ɸå�/>���W�����
�TS��Z�@DYm�Nr
Q�լ�>������t���S����nX�Iݾ�BYVA�_{��O�c��9���wiLSsi�=���x�ˎ|�U ��ޙ�^�a��N�g�b!��ӈm^�9��(T�6-��5��|�EG�l?���7>X̑��\������x��߸��=�}�K�|�#o|�+_��?���������?�������#y�����C.��;/}���(�N�`l���K��]�_Q�����SPO��^t��ILu7�U�׭����i��D��������i�-B�ѱv���?�e��Ɓ33<D)+���Z�/'W����a'�ݿ���I774�ڄt͹j�lS�u����>D
�Ǝn'��4���G�������,��ʺ��,o���A������2#-�R���zYh2�O����Tٗ�1�L�`�|xÂC����\V��X"0���B��S3��b�e�L�(Oym�hnM���[_v[�̙�Y�o٪��E�ڻ���I�[E���7
�)��W�o�[i�R�������6���t��R���09Ņ��ysK�y/ό���v	֣����-93��#Wdj�}w����T��L7�8܋;��Ӛ|�X����I<;"�u1���e@�=A�丘��hB�����1A�x�b+0�j֔ceU�f.@a.�k*ϫEt5_�J,佩�5՗�H�V�!֗�ї��F+�S!���UT�\�hQN�l7�3���D��D���X����l#��F�][]y�*��F*L� ��&;öx�liB���v{1$�Z={mf�����MyT����W�pr\��bȪ�p����kKҹ5?�C�:11О�vT?�"�D��sZ���B�F�;Y���?�LP���T��������t�u���D���k��jU?����>��w+Dao��c��${I^V��A�_��:��QQ�;��Y*J�(�e�v,7�c��,��2v�D�[nd/0i�-��yP���99)ǟ1u�yKvIڪ6n_[s��pަ�@Ϝ�m���e�U����_��^��p������G�z��!p\�j�wuJ��y���"W�V���]յ�@�U}n	T���&�P�UU�2LkR�/@�O�yj��j�}ٰ����U��o���I�q�����)W*���_�UT��P�0T�(�S������L���0��_4c
C�1v=�g{.��ȅ�י�Fq/1���r�.*�_$_�)e���$�K��qt�u���TnH��P�aOc[:Zؑ��K��5�g�8yp�/�<B�@��;M��{�,k�����y�//9D0��ODՅ&�|#���s�5�׬�c����Xz�A�h' #���k��\���­]�g���K���p
�YzpU��+殲�E٦��h�nd���+��=�xr�@�7��<�ݹ���53_�F�'/�z��B�9�k�sZ��1�ٳ�G��lW5�����?���=�����cyu�
��=�	��-���82h
3C�l����N\_���c�>8���9�:�g�mbqR)��zpr���^���K�0a>���� oՐ�Lm�GmvW�D���������X�;b��YX�i!�`Ǟ$��؉��Ø�̖�ᾤ5%SSEL�~�T�ĿKAO`�*�+Q����,׾��oW�d�c귂��Q��R��)��(�S ��i�?M����
�d�Y��f���X�Rj�.@@�F��RB���#sqJةfZU�����7��[�Ib&�Y9T����9XUZ��a���τ$ս�{�?B�v�����-w.��M�x�(��'��<;��d��9޼�VG>��o�Owky��FF/���S�wͦs6Y]qI�kr�։�1�ǔ
<R���ӗk��߇��o�y��(�/�Cqs_��N&k�Jfl�v�V&o>ľ�O�­�|��3|��q.]�ͺm�$c�e�]�L]G������&���nX�uýK>E5��VPZAxy5��U�)��7�b1d��E���[���Q��n����>&τ#:�����7���-�a�l]��w���O���vFF8��i���@�T�=�\��L�J�b]�*D	���Q�}�u$i���]I���
���F��DK�3³�s+�Sܝ��4�ɲA*�QJJ���cuZ9ۛ�0�c3�S8Xן�c&2�C2��i>�T�ە:m�al��P�]��ز��K �@p���������T�i��j��(�\A�v}���ӷ@9GV���Um�:ٮ�����r�#��^%V�J��~U:�u�*R!�4*ޖ����ޖ�\�" �����Ll���XΎ
��-�|����EZs�g[��fk>�m���ٹb����F !A�e�%n���t4�'��H�Θ@[<䷓q��S�V � JG@JW C��@���CpCy6
�LT���J4��7�S�j���~��f%jYI+�)Q5|��g�d[+��8�m��Eleb����- ���)QyL5�ʻT��t���W�=v27��Ɗ@ksb���d�C�@-
��	����3//����^Z��E���ތ�v�iL�ŉIܜ�Ʊ�L	�b���f�ƬxS�Z�k���ry�����6h+�'�'�E��_o��%�;����X��̢�ެȫdOM�s����`}s&{��G6��b�G�V[}�6��V�����H��.�$-�|{L�kO���N��tJ�愞�tm9c��iQ�g��9�Vդ8k�Q�
t��c���_�����8S�pژk�����W��Q~�0�u���.j�~��Cb���Q�N�ȳ:��"j���Ӳ�5�J��	p�����a��qN�AU�wM�U���3r p�
3��4������:ZV�9@6�c���X��Z���K�/�j�ZP�&Y�G�UIC��{E [5�ް��料@��o��M zD�<�w�Zx'z��ڱ*�`��3��møY;����ApG�	m�{����+�\w��-�P>�
�#�>�o�3��$�/}��]��\�[�ty�Q���%D������8q+�#��r�=�����w�5����n�\��h�Lm��2=^@)�؞�r�ϺGq]`��v\����U&�<Q��x����g�j�|7~q\����xYD��}�;���Ѽ�����G8Ϻ��<�g�Qn^.��s�/�����
��˾�\�i�w�#J�Gr�'�kj��G,/z�x��O�}� su�9� �c���7�|y�ڏ�u.��˙�Uȱ���Id�W���e����l�E�'�������Й�Ȼ�cyf�4�$��9��I��3�����>�l��ϙ��=w[�-g��l��P����ǰv�LTԑҞܸ�kHJ����y�f^��{��|�����j.U������Xw�����t�GRe%��ꉬh ��^s�f�Y�}�Z�����5ߪ._�5OM�_�Vs',��C�ާ@������G�"ȣg((|x����i.j9���߶��UQ&�}��3L��1�31����ax�u'0���"�;k����Vp!e��@�UTX�5�:��a��IP�:&/Xĕ�Y��Ŧ~}��/����yjjm��k�*?�5o\�ĥ�����n�p��۶1hJ?*=��Л˷Ry��6��ֻ<�_��w���P������5�A �D)㐞�UѺu�{F"����f��W��?��͏���@���*,�.�X½|��'0pޘ�OL��Ϻ����[�OnE
��q8g�a�^�ej!����%����Zٝ���У/i����ԗ���t��I���L^���[�R8d8�1���ĩC*!����V
c[<��	�K0w$E����I� A�X۪/��gd% g$ֻ� ��HR��3}��I���A�R ��åp.JY]C�U����vcTl�fn���b��{�S���x���U���/���\aj�F�D5zuw`<{�˙�ՁE���˪����L�Ka�\���? 
��j��kPеIDs�b�M_Qrj4��&C�+Q
�y����P����v�j�z�D)�����C o����V��dh�,� ��4s�yS;�V�o�t�� m�5�\ch�yf9�~X�g����\^���ql�waL;֕9���Z���7V���R�X��xo^'>����X_�Π0C���o�C;kC"�L�5U��:X�(���JΩŨ����
Z�ͦJT3����2y��)Q���S����g����Hc�6US�
tm�:�hM�2W1�ML$E,̍�8�{
U�<M��JT���?Υ֩{T�`��Ԙ{Qh6�$Z�!�72œ��S��4���;���T�,(���x�2"ԕI�>��Ks3�? ��Q&�-k��R���i=MTm�9�"9����"F�\�]n����؎m�#�)���(fxy�8&�C�F��i D�m-������8t,�}�<:�����t����@8���o��zC+H�S5g�����mU�eK͑�&:��@�+��z�2�`��A�=(�+��y"jy��S�P��+;-o�s�uc���f�f�ٱ_ ���G�;Q�w�8���V�e�n�F�hE�d�Qߔm��b09q�9�MV��p�b��{n�9z��ރC^�tf����� ��{�R��B U����<#��V֜y���\��゙W,�n��e�[�r] ��Ɨ�l��h�>�<ob�)Ϟ�v�I������f��kw�Hw�ʅ���B�عG}C8�s~Q��ᄣ�@Q�yG�|@{N�%0�ց2����d� �͑N�,f�@���1܉�e_xG��D2+$���>��0�/�)ޑLta��/#<���l{��Gs5*��	)\HU�E�H��#TπHK+"�� @���2�M��T��6�06���A g�g��ko����۹��T y&�fX�������v<�"�=�}Q�)�wh`D�<[�֤P����քD��7�Eެpf�@��pYׁU�Y#0��7��b�.�f�4���{���'�E�,�g��+R~G�L�m�W�6 d���G��ƲT@u�_{�	.�e�w3|Ù) <]��!y7j������ ���3��\���Uy��b����yy��ڸG`!G�.���z����,ɮb�� n^��	�Ew�W���8V�s|��%��k/��X��IK�2a9�'�dӘE,0�yͣY>ls��{v))���q�'�����o[K�K�x��^{���:��*�QͣG%��n&��ѥ[:1�5t�ޗЊF�*�j�U � �������<���ҧ_��O��XF&5x��wOo��-��|��W�:��1�㏇�QaY��Oj� *�-���,�[���&�ɲ_��NV�����`�[N<�z�S܈wN~���.�/�����Q��ev%�K�V���U��e���oi9��N���E�*�ű�����h�n�L�<�,Ԏ"Z�7�w�ןy���\�}��N_���os��%�\��=�9t��ݧ;3x�X�%�L[��'_u�{���E�6`�����t��.-���z]pȨ�?7��;��Ow>��+_�ڕ_u���8z��ʾ1ا$a%�kٹ/�`���Ys�����/@����ͷ#X�������d�i�<<$3����_Dhq�}�. ��w0q�	#��I��6y#�����r�j��1G���)���<��v�O>�H)�h�f�@�P�26%P@�Y,oK5##,ژd� V�35�ɚϮ*)p
�w���R0����̭��kmN+ꤰj�`\�2�ۥ3<*�E�e��2�0;G2N,�u���f�� �����d��{�%��k=��� )���*��y��������@��}�1���2Pb�(�]���X��p54��P��Rp�e�e(����NQV*n���
yJ�m62g��WJv���,� ����@��L�O�7�	lnPM�m-Yob�8Q6�~h;kNN����9K�(��L]f������Ęؔ��E�Z��[3�3U��a��Q��� �tho�җN��t40�N
hKVq
���mO��op$��UD�����VDO��%- �ַ����i����j�����alf����_`�z�p�*�t��DΡD�����j�y��bbF���6z�����������Ď��Ё�S�908��)z�,,����D��	fj;#m�Œ�,�����h�'�D����|���b1%
U�<}c&���g�r+& 0�H�	��*�98a�D�,�T̚��X�g�6�B�u{V���w��թЀ�FfD�M��i������P��:����w�ٮ+�'��Gφzv6�{�w��������t�J�<hn��Gk]\� ���WA��̉5b�m�g�(�^��O e�(t5?��IQ��E��N�|n1/��~�S>7�깜_��U����iy\{Yʻ�r+�!�흚�\����n=�\P���.$�p�c/$�r==���2�.�s+5�Ii\OL�vR:o&g�Fb&7�u��*J�Rt2c�x5+�׳�x%%K�͔�:�Rzg��u�Fbwb$?�u�fL"��y%&�Kq��/cs^)kS�؜^��b6t�dWfqK���J��t��$z$��3�3M��I�az�Μ˪����<�/F��Ԡ�,�ه%}�x�P�Ê��X�<��=�	0�g����2��=Gpn�$n���؛]R��9�����+�`P^9�R
Y�_���n��)dY�b�ɶ�l�.�b�KHcpj�{�>����
���d�(ܳ�l_�R�u��#����կ���5�)����7����$g�DtΊ�j�v�evZ!�Ҋ��Y�U���bv�cII����̫anQwf�Ti�aF��3!��ɢ�gv)g�\�����3W�U��3�K󻱨��9��۹�	��Ȧ��C���!��͇�iΠ�u���	K�4w3WM���yv�J�M^¾^�Y �x����Q�����=�!�r|�N��T�1]�Y���1��frr	s�z�o�V-���)��0y5�&,a��iL�5�'0w�$&�IqZ>�b����":N��kGi��g$R�ǖ�!�L]�ω+�|�M-�<�-�?,e��"��T]HlU=�eMT�ƻ�{y�ziXw@����}��?�S���	V���ܮɲ�S����!|�����������ʮ?d/��2M�oq��X�P�Z�W0�'��qW﷖c�n��K�<K���x �x8^��	*j"��FI�¢�T��}u_B�[|ze�*��;�+n�:c�>�a��4��ǜ���޻'7:r̻����7߷��?L��&O�TM�,knL���{W�r|�n~�/_���>��[������ҭ��;4���t���BS���=�~Q����cֆdꒉmT>`J��1#׬\�H�
��K��T#�j�|ۋ�����_K��~)'�$�]�7)<RK�/�������j(����z	K���o�2zf!]��l&�����J:��0�Kr��v�Eduw�j�����)�<��)��*��]
6Ә8���J�QD4�~�y`nㆋX�^Vn��9&p�kJ�@L��J�XIv�L���� ���l���3�q�q�cd������0��C��
lmfN���bIF=�7geJ��	ف���G� F��̔�a���X��mhIW�D'W61��7���Rb�G��!}㒘ٽ���X�rm�+{�<���X�[Rke�@O�˽��-�/�e=�z��Cml*�9@��4�"��(��_ O�C5�*ũ@ME�بk�z=�ɽ�����V�+w}��M��/��3�3��:ޗ�zմz`D:�-�µ)q��el��@������D�,K���p�����QQ<�7�%]����#\��C`FvQ�δ~s���� rb0	���	\��_�+��oQ�u䘧����&
��wA���o�����׾j��[��	�[��ጝ�&Fz��\{�!O_������lo=F����O[y."~�W�uH��ej�?�Ƨi0���0?�fs]
������}X���hk&,Γ��D��2�em5i��k��r\,׮j���W����m����$pr�6fh�+�����̌�q	�7��I�u	bm�Al���v��/Z�r�?�a�gU��5������:z,���j�v����V�+w�X9~�`�쯜⪚<������6W��Z��b����o{��!;����5�I~��K��F���j˛������1t6�{M�V�ɼ=r>�O\Ƈ�r��X^8�3cgru�F�\��[S�ʈ�| J�����q�J~����'�Ꮕ;�}�~�|w�v����E1�j?z��O��͵��f�f~[������;�F䗵�b�&�]������ś�n�R>�:���n��-Gxc�!^ٰ��6n嫕��r'?���g�������l8ΟK����|�l+?o��Kw���\?~�c�O�i��n>�%��o�6����s;Oqj�Av����9{�<g����ͼ�d_�ߪE���m>�p���Nqn�	���ĉ�{����v���棜��:�� ��f׾���u��뷱c�Vn��ȿ.����g��|����_���7p|�n�n;���kٵx='7�d���l[��K�˵md�\��'�#׻v�Z�O]��e[زbGW��Ĵ��VQ&/��ey>�f,���}l^���S�2n�֮���5[Y�`9+�`�ةL2���ǳb�d����!SX2q� �ZVN]����X>c5��|�f�l�����;g)�nbÂ��������x��M[Ī��%���~%筓4T�ۙ,���=;3��7��@�)�r��ƉRSƦrz�Q6,�Δ�8��0�^��Frl�p
"Y��S'Ȼ�8{=
�Y4f=�V�oK���l�$�dϊ�T��ѫkw֮���%Y�d�ma���̐k7|*�'���Dտ}��S��p���5�.�ad��уv]��
��"<����4N�͉��y��Yz�J���we�?M��N�US؛���Z���W I�\��\Mp����z�[_?R�kڤ*�Բ̩F�
����?���_d����&��s��N-�D�R���R��T��Q��o�Z/����u|�����!�fm ��x
��[؋�
뿚�2��*��nDY7bTj�U�@��M`V��\�r1m��^�D��Il�c���Z�uI��	��N�J�y|����dR���˥+�%o�p�]�f���N�����=�X�������I,]6��>5�fWa-/�/ߎ�"��V5[Ov!�oi�y�0��4����9� �!�2�ث�k���	L[�ؕr쇵r�|�m;v瓜�}\$n��g�L���ҍY�������?�@F}�nw}��֓��~t��L����;U�W8v
�僯��X�=�.EXvH�N�1�N�Ŵ�M`:�>��`����+�DY�ih%��(#�dڋ$�Y�hgO��� �.�\U�R�Ƣ��B���0&�#�f$��bid$��b#�c��X��14��X �R�clP�k��-l���/�%��@��N$�օ����V����I�bn(�tH�M�G]#~.�8ʾ�>��4�Ĥi7�ˉ 9w�(�
)�{j11o�q�č1r_J����NF���}&����T}�;	U[�@os[3-�ښ6��h�<5D_A޾�c�&�u�6A�:]c��5��7e���y~�����++4�x�3�Y�e�K���P3wV%qyF/��šQ�bJ��@������[��H+S��u�Z�� K�������^̵����H�z�p���e5xBk�<�]˓&[W"�pq��j[��� �Vi��	�)y��^�
x����@��/������Nos��:s��U�s�;���H�t����ҙ�I�0gzA0Kj���kstY,����ȳl��F����3�'r����k��J>��ȱ��c���k������b�\��d���(3|�y�����!���Ss�K r�l�'��iCg���֠=t�ٯc�!]�QͶF���{�S}�N.bTL�֚��of}z	;rj9&���a����_�̡���ʾ��lʫgo��o�1)s^;r�#�&�<�X�{��c���ؕT®�R�dU�+����I�}��Y��������꜍|~�*�G�`u3�+z��~ k+{�^���h!�����~�ndK��UX�~1�
��s�2W6b��Q�� m�=u}�XR��������C8�4�=ս��g[{e��	��6a6#>Ob���=�")_�k�?d���k�i���:pS��]�g����r�0^:��W�e�Ťv)#).�!�tIȠ"���|�:S�Y���Y�@�t:%$Cpd��M���+���M�x���˚ץ�ʤ.T��,�*&?#�ƪZ*
K�مN2�N.��b ��d��T5P�R@aF	yIy���::���%��,e�����МQH���1�Ď��8����0s�6:�
�dѡC:I�Hiׁ�h�b:Ց����l�r�yl�T�;f� �`ֆ��N̢SJ)�]H�{WҩCq��bӈ�I%+�������J",$���"�����)��5w&Pל03Ua`���j�Z��m�H��b�ĠQ�Y�j?����o��������	M���6�P�m�����ҙ{�$ݞ�S��^BLH"9�7W���������b�~���Ŭ9k�;w5S'�g҄9��<��RXQA�P
�<(w��&:��1x���2(��NX��{�����sؼ	�^�Ο�gr�|>�1���K�32�N�y$��	,o �[�U�8��a������_ź�W���w|�KK=y�|�=�|��U� �j�U�v-��󶠡""���D�DS�T�6�Y�����S�߾�|�Տ���%�
k �r QU}���	���pOE�V�Ծ�A����^"�t��O��^�
G�w�M����Ѕ�0v�h���ήE�v�Z6�Gq��@�V O]�?L�<E��h�X.���[/�eSc#{b�9����|����+��Wɳuu�8����	*K���3�<Y{(���H��Jh~w2'��@�L�K����4���X��d�<�*.^�I�.fĔ����`>���?�(�ǟ䦶D�닥��]R	�R3f��st�n(>j��O��62�����$�Ij�F��6�m�,
�L���i�2��ֿ���\,��픁�|���Qw�Z$}7m���H��;�ƶD���^�LI��	&V�[��䌓�~��3#� Q�J1����N|b*���1����-#"[kY�D��2�e�'��|�*+{����\��'f&&-�N��\I�P�8g����ձz�'��ܳ/�nb%	@	���9��y
z��6�(�ZD)Ɏ�L�����>1�E�-��?cC:1��S����y��U#�yzymd��@�s���׽?{z�՚�ט�@�:�N�j�\׀�&��������k��8�'�	�tx~t_��Ç[��27�sc}�0$��Ձ4�ڐ�d��<;Ukg. ���)��`[D��3�U�dY�N5]�>g٦#׬�V��U�zZ!�iPj��çD�?�����lk]V��Lt�vu�It�/.v�Z�k\��`��kh=�UԺ�fZ%���4�.jD�lS��'�b,�]�����g����<Ȍ-�"�8������HMcQY4�\���Ĝh��1άů��y��V91^(�R�XTS�
ɧ�k��w�쐉.�d���Ky��%��zn�vG��͛���:v3���K�����X�i�W�A(�gmp�>IK5����gt57'TX'�����pR׎���oc�i#{J��UH�U�Z�%b�7Ht	��q�x��H�2�ٓ���LNeqtk�P^����(���!�����X&�3�ǟ	���+,�i��.��z���0'#���1̎�bRxc��π /�E1>%�%��,��c]j������l��bcp�	�(��|�U尣(���,��PY*{���ڵۺf�.-�E�ɼ?~)/Tb�(��YY��̆�T�îl.OeCa�JS�U��Ϊ\�����"�j�Ý�I8���@S1p�	r����F�ba/ƃj�0����s39ݻ'��bor.����0q&�ȎP3��-�l��|�Z5�l72#��\[�6������^��R�>��c��'�i�1l�����E���Ky�&p�oI��!�FDؘd."y���z��<��˷&�
�hbG��(CG
Ch����ڇ�A4EiQ6|l1s��Ѝ�Ў�q�=F�c�I��Q���[�gF��%A�&8I~u#�E_D�w]#M���Ɏ�gޤD���gI��^�x���i`��\����<Pb�}�j�c팛|+.֮�Y���#��a�(p�@��b��(0Eb�\��(Fs���T&�[��y�	MI���gs\�L�@[ɞg/�[�1����+ t�{����ȉ�p���!W]I7�5����46����/%e=�����]*)-�#�����|�FB��R+y�KT� o0���X�b�Gf.�U͢�G���!�-<zܛ?���9xNʞ)	dvϦ��Rl�@��k5�aU~�5?{6���+B���17���7?}�_�͗�}�o?�Dk�ǿ�ݿ�:����?x��Z_=5��e�rh�0�.���~+����.'�|���(�������U&��/�b|�Ч��y�FyV�г���H��ALu=q�uD�TS6t�u�Ȩ�&.�6�:�&6a��}�97}6/�4q*����z�O$Ӝ�Y߫��} ��J����<u���a�rO �G޽t�}Mul�qg��[�9���I��̍�t���7q ��WS�3��a�؛Ō��+�CB�6B$������H:H^`:/��,g+��X��S݉�&����1�,ڜ��*��|�U�צR;"��}2H��%�{7ͷΠi���ˁ<�ם/�if�2�J��?���s�62M˧и`��<�=d�V��j���J5���	@�[�?��^�	�9ٹ�+�<��
��H��N�P�X�����X��θ��a��/���K�U�*7WGb�"	�t�Mi���(�P���h�V9Qn�qR�VZ]v�G����`���kk��(IU�g!J���T����&�aCg��Y����@�.N~u)��K	^R�(�	��c���Tc�
Q�ZZ�\z�Zd5*m���c�cl���V�z���h>Ô��)�b�\�&��D�̩Ѳ��ڕ"W9TD���!��ޗ���0V
eyj���[)���W�7K�����F����8��u�~bE����|���W�puF,�F�s�)�q	Nt�2њ��}���-��<���;�3001�Z Jͭu1�V�&�$���6L���"U+��T�o����B�����m���jU����	qA�f�P�%���x����`���P5+�U��l�*j���ElL�q���A�����E��Ӡg)�����e&y ՚��4'��}��?�eU1�s�{���^ ��6���
y�O�?A�29�29�r��D��R9�U=C�����4�m]���$�N�k'���ic�k�V[�������3�ˏ.rl�-�7"���Y�+[�Z9�����B�#u't�8%�wB����������m-8*r�@ �)��'�S�1�y��ư�lʭbyp8�O���簤�����L��crD�6��1�e�l��ȱ�#8?g2KK�X����UM
L�TBgn.���Y��ّ1�E��P�t#++�E��lݟOo���;7�t�*v���n�p6��rm#<w�������~8��_�o����x��f��޸����G8]Ճ�N���RN�O�����k�����p�Y�?��������w�/?�^����l��L���8)������%�5c�2R�EvL9�At��#�ۗ4oS;1���7�l�gβ<)�,yo��'rm�(exy��S�.�$7g��Hr�%�ÕLwOr�)
l���2�ۧ10����'�/P����k+���l�2�>Ed��#�/�L�@2�(J��*=�!�U���'�ڃQR�n���K)C<��L��ls#�џ|�`���(�� 4�g/�}��VL�g4����Z��ɍÈ2�"�+��$::�*@�D���" f���1>�VY�.�������~��r!�ƃ��8b|�7q�M�B`�oS{<�l�0o�+?��!Q�:z�p�jF+PiM��	ɺ��Cp)dtMo��:IU^7b�
���׳�;/޼͡3'�--&Lާ��N�����w�.�⳴�����E'�����F�i�VJ�K�q�`M��IV��Y�	�;a�H��+��D
ǚ:*@�'�!R�C��ݽ�(s�!�Ӎ�h�b�v������:t�F���5���������G� _
?����j�$�.=H��'��?r�u��u#����f��ôc^�
Y�g_�t���N��W�y�݋\�]n���~�%?��@>�o���6r��o���O��_����_r�Ox���8��;,>t��7�y�4B���m8��d>��n}�na1e�D�խ��^�$��T�(�&����CP<|8I5�dUa�E1 u����ͥr@3�Ǝ�bY�c��ʗ������s_ի��_������Eo���Zڠ�n��RA��+�ѕ3�ӝMb��pg�}0�=�q�+���ø��-)�.'�p�_�,������~������q|!�)]��.�U�[i�C"��~w�x�)�\��Ã�1�?�g/�f�$�-������Qr5���"n��ʉK�^�L�����r��d�x��~�]=��ACH0����9��������k)�j��)�ӏl��|$:���y�b�≩�bq���,G��Ta� /Z���hQ&!VNxY�kҕ�M��Q
��؀pOO�C���Ѭ6U�j̔�~UC�'0 �\�|H!2e���Ɗ��QY��:��o���'?:�2�ʅ�y��/�JS/�g3w�f��NsA-����+�ɸ�>���TW9��1�1gһyin>�Yh����j!�Zj+Cf����IY���������]m�P�T��<��"��y���l�ˎ�c���L����1W�Q��,u������������?���j�9-�[3S9>0��9��9k~Ҭ�:Tm���� �!f- ��ʲ��.��8����F��4Ԗ�d�ZF�*�R��@�W���JTM��@��ϧ]�֐�'��5�ῑ����bE9@�߲]���s�,'���d�;��)��_|
jLe?5�C�ڰ6�3f%:����rxۙ�go���."�֦Z�VPT���k���
�2]�}4�sinGFĲ�)�U��Mp��ǔ�`z8X0�Čyb�/S"�^9�^�V����.+ڶ�ޯ��FQ��|��OA�L&�&sr�L6U2�΅�����a�������k��ɜ�!�W��X�]�V�W91�Q)�p��E����ѵ��,8�kǑ�Jl��j��6s6Ъ�*,�n=S��w�O��~=�:��� �����<�xe�l�&%����e�[3�����.eG� E�X�i������ܓ�+q���۹��b���rg��Dd2���������Ifp;rBc�O��cC
jӣs�/���˼�� [J��֠�,�Ne�a���KlZ�A�"�c���ǱC�E��ܩ�\z�4��>����X�xv�l��������ʖ��$m۶m�vI#vl۶m�v2���Xgt�x���y��~����U���l�V�]U̭�Hq���O>���;ܾ��.������q�];����]:�˯>䫏�f����!Zj-3�'�����L�2��"�S��T�'Q�LMJ.��ZɌI��w#�/�:0L�?��.��xy�U]͚YSY>{�62a���-��Ig�FJK�IM�'������w�<a*�>��d�ܙ�<w���gҷo�%T���HZj��d��1x�Hf��F��,��w�"m]H�
�_�@jV6�^�xy��H�O8n�8�����MlL2�խd���������6L셀����r�
�����'���bd� �h�|���"�;�h7q�{80<��C����Wʌ�?�>a�������"y	Xz9���M��`O
H�)O`��UZ(�QN�̵qb���T�+�o�]x��=���ú�4�x3/>��v僃��PP�R;o�J��/0y"����Y���� 6��1�Ο�)�=����h�}\R��I�����T}��0g\O3Ƌ�4Jl��ڤb���g�0S[F9x1�.�6�oW7b=��ǆ�"�Ap��� �Bb�K/"8��3[������K+�������{�s�z&�(�lP�b�R;��2�`��Pq��:q��}Ae��1��÷?7��?��Mb����_��	������'���W����_��.���{x��?��Q��Q9j1Y]��l�Gp�1x��#����Fh�e�Dzk��ܦ���Iʠ.;��"g�p�O�k�:N�G��R ���)��4|J�i�Ț��9�џ��x�/��Q�w�w*�D/"��,�?~��_}ÿ���p������Y��[?�ȩ��q�昙�}�&��E�f^v��"z?a��C� �Er�,���C��μ�}(�hů�ۜB,
�0-k�GBQ����ģ�������d ��S4r��mf��=�^5��7���?g��B���Bo<�����|�[�{���%�>�#�۩�DҀ��M��h�:�ӸtmL�Cz��1���������=��䎥�+vw���S�d%�
�j�x�:&Zs}��Q���bd��zj�4T�����Z�����oV)=c�z�(���(F:M "SHv�eb�j��Ű�4>�r���4E'1���q�$�gհ .���]��
amHӍ��"'0�/�1��,ŷ���9y�LMc��F��ųF
צ�X=b<K�����h3{�ʰ[)hP��Ы��*��GO]��Mp5��Z�X
�9�_�J�~�/�'��Md�<�yׇ��@�D&K�T/����b����Z=��uC���>�T���h�..��5�������7!�-5�t��(�c%��Dޣ�\Wk�47�o�B��.Z�z�f�#`׃ GK�lM��r���oo���)&�ؘckb���kbf���G����o���*��Rf��H�Q-x�1P׍��!'>���@b}��4�S����+�V��8�	��}��3x;X�)����x:�o�������z�v��8Y��b����OA�j9��7�Z�շW����lw�M����B�wD��w<cR���D��=�}M7R�g�J]cV���2� O˦�A^7��xS��Qʊ��ꛋ#�6���n��	̍LeCnwGO����X_�zS�79���j/'����Ob��a�� �HΣR�]p⬁�UaJ,����jBEKN��	�Ys�̖uvṈ�g��9sP7H]S)��!:(rD���翷�r��$(�{I o[c��E0�4]?KzX	�[Y�,:$&:���
ҳ��O � �Ҏ>,ܳ�C'���k${�gOz3l��v�@��Y����wŠG���@�{0ў�x���9�?kFN`G}>���mi�,h�3qA���Ge�V�@��=�_��5b�OcԢy,۱��}�sWrk��7����k���Ч����J�R_7�����U��n�b@�i1�ׯPn&�Қ0��&6$Y;R��"ϝCBbIqa�f�P�FEB�ʊ�H���Z��И8��ݽH�2#�՞��i�^L�j�����C�~�)^}����`��e�3���A��w`bK?�ΚM��a֖������BlYU=�������I� $&�����Iɢ��/��>L:�u�W��B�����Xܼ�0wv���3{g����ciGc3Lj��q1s", ��[�3�c����o�Anr6���k� ������:�7`m�FQ��IaY���d:E3+��McZh%���[8c�o���-�6H����42��Bʭ��1j|����qi�4�ǲ]��{w}B���e�x�4q�wG�Z����HN�ǲ7(�C�ٜJ�S��Q㪽g�n��	�(�Gs�.@;�rB1�����c]v1{Rr���=� n��q�%DK�v�Z.q����kf�6q��x�����Ȇ�F�L7�b�O,�����c�v6㡤D����ip���G�[�ȓ/6Ǐ�⣯G���V���T;ægR3r Eæ�9p�RQm�	hj�W�Mv
͓�x��X�A���_4��Oc�q����$u�#q�,҇,#g�\��.���=|����|���
��A��R�jk��*�1�p�g��]ĵ� 3�O'�r혾�8����d�KB��Ķ�k��i�#i���ak��2g���Dgb&��WJU{�ǌ�@�A)�/�E�8(�[ai�s��[����o ���"���ħ�|�_|�w���<�i��A�ݠ�;���>y�3:8��eSoN:�sR��%�p^u��I)�*e�3��u�����T��p�k+&�e���d�Oc-vU���+ƫ ���ItM�b��~x��a�S�W}+�CG�1|�C�3x����S/���/��Z!�~��@��5��>��ŻSh�TNDmu5�T7�RP�CZ1��@��	�􍠇(�����;/œtuv�&1Y�" .�}��j͊�c�H����.�J�������S݁�z�8�y�[�FUD������S!�Jt4)�+�ѣF�K�H��c��=�&2\ i��>\*�d1 �ģ����P�����ʏ����'v�/C&�2��N'��ы�����vc�(��F�lc����IeMX��=�1s᤹+��[-��T����V�Au�7� /@�+��;��
���F��X'�� *#�?!o����-� o�@�BQ<'Z�q�m�|��y�d�fy*��:]��o���4�{0"΃]�)������4qoF����Y)�d��U��Fy���l8��B����[}#'K=��{�ji����ֺ��NK��※�+��.x�;��ꀿ� [U� Q�����U�\��^��gn`�-UZ3�.d梔UW�^wK��:��
d��9[�j�$���[33���;Y[�f�{W�=���%1,�0?w|=�ps��Y����7�<���u �ە�ܝ�w���
ok��-��S�*�$���HR�n���:��T0��L�YQe�[��˄��"�K80,�y��M��ρ~r���46b�<�9��^ݭy�<hoD����De��|m�v]3�ǈ�R���g�l�T�5��t�N�G~�u ��*��˩�2�w�����L�����&S����>��7�&����:��$�#R.�����;�Z�zZr�Ď}�4�1=�ܤj����|jl��O���V?��{�Gww�J#uJG@Qً�fhA���e�skC4�;;��gbM�8�y!Q��{	�8�i:!/.�������Ͱ=�T�� B�~��xg�P;��m�w�!J�<�ٚd������<����`TDW�L�)�8�Q˔�dZB���i���1�'�����>:�֤\z��(�I�@``t�@�t���	�xX=�51Y��j턯�'i^�}�'*���BZb�
O'L@�O�}ߪ�L4�4�I��K��g�E�
g#q l�	uv �]݇/��.DZ	�� z�W�NsG
D�UzzR$u�Hʣʳ����a�y��>��}q���w�����~��.�r��,ZEcE᢫g�v�g�T�%0N�{�o An^X�Z�'�r�#��[��/7W�0��f$e�U�&Z���ظx3QX8a%�W�]i����.�&f���Sμ��C�<[)/�����>O��e���L��u
 �΍��8�͚Ñ�Y�|�mcÎ�lݱ�93�2m��/�������ɬ��ٜXM��/!Vx y8�K=v}c'N�+�✄�y&p���F��Q���q]���R6��p�:����<i�)v9��A\s��e��1�i/-��Uc-�u#n�;k��n��s�č�.�6`��%���/�삵4o�m��m��~sg-5�q�U��3��3gJM��5�쫔�뤜��������:5��K�X��b⬬� >"���x��|qu#,���!�����_����y�<<�7>Z�����ʵ2�&�R5a2�f�%�P����@x��J3�����~���4q�y?�>�ėL��_�`K�m	xVT3��>c�Pk�Ɔ͓x����� �����g�(DjC�^�_�̩Z�zw�4������LV�XRv�<�	�M�L�����#g�=`� � ��K/�*)���2�b����m�^L>����}0�'q10�^�u�`��@� �/��g|ȇ��|��|������ Cz�� �>y�.�sX>�)�
��-!�W�ĳ���By�͇�-<x�4����8��i)���*�0���c�a�FBcjj�.-$� ��(,S
1J/�<���<��s�ETv�+<pfV$�d�/[��r�n$��h!3�S�7��D�Ӓp���L�)��Tt���!�K����눇��䍙�֮�X������̆P�T��(1B
�b|b�bDI���.��dh�����Z��^S�空-��%A��E�Q��D��W��Z1$u��K�E�����S�!�`���J�>V�'ȶQrΉ�M%p'Ǐ�i��^6Zʲeb��ɾ�Ȭ��e�dl�J1�j`��F���l��g�ȶ^���e�"9��D�I�e��yQ����3�Ԍ���.�!��'��+�Q�Y���,�9c�A�q1�jp��<O��e�zzڵ�m�7f�k ��r��8fz�ik�
�m��P�.6��z�B x�H���/�Gy��#��׷���.�������_B�U+�{����5n*P� �����
"�ƹ)�r�6�i��jyژ�Y��  d���^bh}�	�3"�΀]���x����� ڦ�V=��@���2T$R~����I*i~\`ʳy��>&T���BP�,u	0 U�Ԃ�B�Bm-  @߿�p� A|F��^6�����$0�` 
�OG�F:�:���(�Չ@';1�6�8��9��f���5���@��@/{��3�IUY<�g�vg�P-z*�]�U/f��sg~'Ƥ��6�!i^4������pKkf��3_�U��D�}7�i]�
�6���D��֪;_Aކ^f��2��ЎM.�Z����Ŭ
�b��gMx:���!��E����8��ȵ�.�sv\�s ��2i��a�3ʴnZ[���ӷ`��J96NϘDcs��Tp�fB�G��1gz�rZΥ���9���)��:�����`�N����DRB !��C��� (���2�}���� ��H�k��q�`%����ې �\{Q]u9��ϤLRÂ�}X2�����z� .m[Ą��M�9P���r&���s�L���i�ݳ�(�	�N�Y�F���%�p�l\Ie@j��\�Cf��3�V�kK�ĩI��$���|k[���tq��Óo_|��y�����]'�ƁtGwm�����yi������Enx(�IQ�-�`@I���TD�ndA��ή��U��F���8��L��3n���?��_~��_��_���{|�k�?����`��QDع0�} G����&�<?jrr)���J%+,���0��Dx$׈����I��'!�~L>��+�����.� 5���>}�����OM-���h�`l���0��0f�`B��	��f�u�i��*� K���Ķ�|���|��'����_s��E�M���c����M�MG��&��q�f�Bs����r�543|�0��S3c����Čѓ�+��#G3y�h��Ͱ�:��S�0z���wϺ��c O���q�ȇ��<a��S�"f�"�Z굇��<0 ���¸���6��V�\��笭/�-=��8�r_�����,�8c��i;�.𯖧l=9&��ؒ��4�ua�|���l�q���n�pc��+2U��
�x�f�Ӟ�F��8�n��JD�ԟ�`��*b��"�ȣ������L[�ū�-�_&�ѣ~�\[Aj�l�&*�ͤ|�l��� }�
5��|��>��އ#WC��1�[/�[:x�Q��$�۞J|CI}����NQ�6���ͣx���^� ��\�ok �m�-C�Y����I�?���3).NP�h�ڇ߷��͔�Ű�+�Z��܁#�/n�3���f-f�k~9I��<����������ܳ�yc_�w��P����n�sa�Gȟ����yJT���#�}�
�}��.��%p^m��
� ���0<��v>\o隣7�<��r"�����>��'p�/�KљL)b�
��6�q]#�=*�f�bx)���T�UR��z݄x,������&� ۬�b<J�	�MZ����e�����x�~���	�%��H1=ě����c ��!X���ꏛ(=�ܮ�֕W�fU���� �B��h}s"M�gwYZ�``���T@��0��&:�XX�dlE�U����Gj�Հ�B�@�R�Qp�г[e�o/}���~bx������'@��d%�d�D�y`�����"Z)��tQ*��nڢ/ޒ��@��&�7͠�>*��JͤBD(�� �q����w5I�Ʃn������)�r?��מ=����s`I54`�x��D9�y*��n��}j|^O��4d���g��Ѫ�o50e�W�[Gq�s*�S�*^�y;��D�����~�©����Ǝ� o��{�o`oo���9�� f�ؒm�C���b�'�Ƶ�.P#=]�L��3�Ӓ�뙘�`�"�)��?'�����X�����hD��!�.FZ�OCZ|�����ah�#�Mf¨p#FDtK��&cbd=�g�D�bHd��``D�tE2,ʜ���2:ފQq��n��>8Ҙ��r�C��b&b��64ޖ�;�Bl���!Ć�@k�=��s1�{6#�J��ڎh[�m�	�.H"wwwl]0�����_O��{Y�αk���U�1���"j6�j�m�����I\��ƚޞKs��ӄV[���0G�D�}q�5�S�/4�O^u�*Q��U+�rTffGe�آg�j�<K�4��鐔���.\E��X����q�He��rB*��5���>�3u�&Eh�o"G�TK�)]�Պ�¤���[L�i�zQ!e�R��&�Ou3�X�{����]VE�>S�o�l\��h��9qlܢ�+P�E o��+}��޿���6�c�"oY�����8�{g��c;�r��1.l�C����TO����<�f䋓�y�^�o�q��߽��Gw�䣇�Ǐ���K�Y<��:����KYO����1<s��ܾ�����Ӽ~�2�^���O�\����<u��6�c���w�0�0w��X��0;Lld��QY6��s��o^��~|���Ͷ�c(͈��X�tq*2ũ�W��H
pcڨ�lQ��3ǖq��jΜXʃ�۹o��lc��i�'��ecM������y����Bj@ sg���7����
�c��o*n+�,������^�qM�W�鼼����i�\9~��}���/s���o�����8�g۷.c��\=��7���Ё]�_��� m&nSi9��������ٳ��{�ql�>m���G8�c7{��dق%�G����Ò9��E��;�f�$����/w�{Rqx�瀯�����?��>�ƽ��Iga!˚��R����,�'�2����&�d�
vn�;]���;�lf��M,X��1�F�VYEU���q�9�5��a�����tn��sSt�u�dnx&sG �O*w}�Ey��AI�H�{�=�9��1�0:s�5��Ρ�����!�{E�C��
37V[{k�V��;��яU�Z/�";/�}�#��\|����;Wƙ9�81A�l�D?S�\�H΢*%�h?q�<}		"*2��Xo�3��KLu"f	�X��T\Ũ��࣭���;c�$��"���5"i�L�/`Мq<|~��L?����u�"������y�!��P^~T���ZcQj}+ٝ��K����1���;���㵞�%�IhN#�u9���Lֺ���Ķ�#�����-����f�{�
��L'�k����)�Ż�^+h^X�}y�l�b��Ql:��M\��]7M��m��3�~��B���#�}�Rw�}�ғ��:I<�V^��s�p��P^,�繤"�-m�~n5�|c�d�͋^�Y�˝��Y�G˫wZב�v��I`nd:���Xޯ��S�1kF'cg�ex'��;�(.�fר8u��q�'%b�B��L���0�Ȣ�o�����b,��9�}b0���ⅱo澡�y�����[0~yR�B�|��m�J��-�b �Dч��.�2Y[jS�=���I�,Leh��Te�R`#���r�a��d��Y��X�F`��2ٿN��;%�"
���(��׳�z�bd�nț$Fs�&L�e�\8V�l��eV�L�!�2�ܚb��983_��0s�l�k"@hj�zS}vrL@t��k۟�*���m�{9��RK�}K*�\c{
d��<5���z�b�C���u6^\0�M�I1�Zj39�-�)C%qWq�T0�=
Ũ��+�=��;������7��F�b��ة����Z�V@�
m��C\�' 28ԕ���yau?��c}��i�#@���+�V3]�����X��X35�@u�����B��I.��YRjE� Tg�=�3������r����ޏ�-�o�Dk ��C���������aZ���#�4�=Z<�a�\��Y^&��9n����������8�'���!���A�����@���`�?;���T�Ɔ67���<������fJ�/#|��N]���"�^d{�錟d[S�[��J�۳���D�N���5�S���R�[�V�q�Ŏ=��7�������¨T+j��hs�a��=K�X#жX��R�8yke�M�L��D,{_O�V�L 5��D���2����-ep�\K9#O�P���õٗ��I D��Sy�ʖ�]��纁<)wRnN�V<��)�SK�����NL��5Lʌj9�,�o����j[Os-(�C�t�8�ӆ�v\2r傡'��3t*��[�е�^tǸ�>�8q����O��䙇W��/>s�7_y���}�m�i]���81u63Ř��(���0����{�2\��]�ٲm>6�b��I�_8��~�TdD2��V�����UZ�1�(�7�-�������?�EѪ�.�$��G�|�Y�v��ư��nnc��&�Z0�w^:��o_�˷.��ۗ�쵳|��%�������>���	}E'� F��s*Pd$�_�ɽ�;���<��v>|t��߻³���/��7���'y�����_C��#�N���Q��@��#e�qTi���>x�c��|�k�p��}N9��cX�`%�1I�jle�����,�]q�[V-�w_�o��G�~�~���	?��/��o�����*��3t;�l �ŏX;7������B}}=����VTR�[DQv�eU�$�C[�
���L�`���,�:���XJ��:p0��}�go=ɹ��p�&'�_��Ż�>w�S{��f�JfO���TԱ�m����(8���Lbc���ϧL�wEe-�U�)�/'/-������	%. ���Xv�^ű�Y��jq~6Ű�#����l�Kb�C(��"Y��
� ��f�w�lז���Yh�lk&�-�`��$sw�	��4vd���f���&u��܅Af����NS����؎#�����ȖFS{Z��,)34�XtM����b}k��̵I�!�ģ��xm����3<����s���k�)#f�9�G�_��c���l㳟�p���l����I�	�HD�B�;hS�+o�������&殊�a`'C��c��.}:�����aW5����nI%�_-���ȭ�fͶ>�J��"]��pD.Q�]$���2VD7w'`���S:a,E�D�N�h�l
G�'�q(>��879��QZ�Ui�o�N����v�s�3AlqO[s�Ɵ���<%��rH��ݵ��CY�(�7������!O�V���� ?��]{h��>#���mx�K^�z����Z�0>�|����A����U�d�l�[{ss�JΩ�zz��s�刅�<�Y�
�x�CR����آb�j��j�+�!.1��x�#�p��!2��x\�@���*E|R,�iqD&D%��� �$���8��c�u#I^J���6�Nv0�"�D OuQ
��Ia����33l��0����T��'j`�2~�%O��
w� �#���X
|�H��'Yψt1X�R�kŀ�
PU�1��c�[�T��ni��.�F<�AbT��u'��ˈIb��4Cd�D1F�B�k�c7�ٞ�>��Mc�x���������5��cƱ~�`���1#-����c���E�_��&E(Q�{�E�	��rpg�x�j���U�fZz�Q��{U��Z�Tw�i#N�QT��f1�gTI���Vy>�I%�/ϡ���A���9*o�(f�Fk��Z�TK�j�S]�;��5�fnOC�	��fh�7[;�3��%�,�sbV���x���d=�=��F:zZ�zu��=���A�W/���2!ю99N,-qfS�;'�r}b4�&EpJ��N��Ei��(��V$���4�ڒ�W�3�~G�&?�*���|�'�o�f�dh������2>ߒϣ5���.�GsxC6o���Y��!��6���2��P�;�
xg}�m��ui���ˣ��*�w������Z��[˒yca�/H��)��$��f���T^��̋3�36�S�}�����J7�U�1�Ї�>4���hA�@��)�� �qF�z��%�'��ʸ�<բ�x���Q��rwj&��}�aE��)}�ii�=K;VHYU��&_t����j�`n�lSR�	li-yZ����cRg�5���R@�l��i�ѝ����vޡC�YB���ar><����"���$��O92*}�.)���~�Xji�T˝�vRG��� �5D.��qQ@�WM]�Qu�O2o�]�ц��rc%�G�������OWW����z{{;}��aĈ0�\1^�!1���Mc���I����_�DFP��J}I!5����dj��$ƑFlb�1�,o̓#�ը�\ʪd��?�<'L�ҥ+���|��^}��_|����ǟλ_~���8�z#��;yi�<�j�LGo�Z�sn�~��M~���|��	�}�/>z��|��?{N,ć|���c���D���V��������ݧn���{[�L��������}>�����櫗xﹳLi�&�֝;
��W:;jc�6��g/�ķ�~��C�Y)�2�m8������ֲތj�ϊ	3hC9���5�'���K�8	��ćFRS����;r"3g�c��tΤ)Sٸk'���"9,3WV�Z���;���p�
��vq�ꀹ�&&j��8�.���S��ffg��R�L��*�b������И�ŒQcQ����>�V4�Rޗ��b���0�OCj�2e�p�/ZĠ�"��#Xޯ����|��x��V���`bk�� ���5Cs,�^وseha���c;l7S+��ƘFO��Yb�r�w%��T�{Pb�H���䋽+;Wjn��d��#�W):���e��ojM�@���el�_bdE��G��5ɢ�c���p:jxS��a��D���9�7,��
y�*�Q��� �'�:��ȻU���=��^r._+|�]�z�������6s����� �0��2(���@�O��38��8&��ǘ�+�r;��la���ߟ�;���V���w>�ˤ��j�f�d�O�������q��k?>�G��1{i4���2|rS�%q�A>?�Z/p���S^T���0'6�[�BB�`����}�
�m�D��yD��O`M'�����ƽ���Z�k�Ijk�}��M�Ɖ	ӹ]����,θFp\u�[xk�	n�.|(��E�ފ��Rp"�\����};�����ѣ��>��yƌfIj%/,��G^�ܼu��/�vF��;��W_�cw8Zџ�Α�ȯ������^�X��;sZ)[Q��㋹ ǭ3ba��K* ���G��DzG�ѐ��E9�K. >1��@<�|#&6��h��(��)N��(I��	��'6؛� _�<ܵ�F1�}D[����L��*n�<?C|���H�ƦڌX+C}mơ
i�/�⑩V!;#3m ����L����p;NQ��TQv�b���x���wC�N���A�_��"� �/��� ��_�7Eߜ)b&��T��}G:91#7��c�8�r!g�����}\<v��'T��:z����p��i�l��Ι��>��9�L�,�a��!��t١��]��zQ�}]*�21:
�T���~b��{�����;�c�q��7�[��Ǳ�Al�t�����^j�`/���䩤�S8jM�i��ch�/��fq`X1�3\�����$7m�pxUݴzr��>*F��o53�ĥ���*tcU����s^���(��˛��e���\��E`mw?,�_�*��H	�<Q�o���jU��j���p��[��C%�.�?���ί7Z��b����9��糳�Ej��|�,���� >?ן�N�������x�"�����3r���񟞪��J>>^�g�
�d_�����=��@?���c��r��ߎ�}�/������4���$���LI����5G��8X{w�.xZj�UlD�LDuӪ�P����TK�ۃA��\�Ĺ�Hf{�dN���-m5�[�'�-��TL�� Ou���R�x�UO�!9�
QrR�9#��4w���L6��S�O�"Z����2(������}��;qV��q�vJ�Q�{Ǥ����˿A�	��tJȩ�>�§�"_�i��Yy�����@�U}<+�<�<g.�q�:���mZ��YN>T) ��� FI~ �6ں�ܗ��3z&��8j��ڂc8S�ƕ�&���k1)�Uw�_0��Tdd�RRJ�8�j�ZQICA!�I	d槑��`�xv��RJWBҙ����E����OJz.	iYD&��Dj~1�%�i����~��,�(��<W�"�҇��.+���}<z]���gx�͇|��9���E>���x�<���`~G-Q�d8y�`�A� �
�R�˱��~p	�֌�����<�����sp����b��Qڶ��D�<�m�5�(=�tۓ�~�� ��������ʭfdio��4�Б�O{R6��a��꟒�Űk��*:_7/m�����.������q,�1up���O�	~&n4e�0���Hck��;U�7�	��̘��P�ER1�olj���� ���I��4R����z��2�@�
~k#�.�2 ��F�ߊX�߈4��(I"�-�D�15�1�ɝ"OoZ�����%5 �ؠ`�ll16�S��/v�@@�D�TĘz:�x�V���K{���G�<k��	�v�$ʶ$k{Rm]H�s%�΍y)ֶ��ڒjo��$Z��~r�6e6��������	��Ȼ�w���M-���/�D����۪2A�(*��8k~򛏩	�F8��T�+Ro�N���bb����R���}��^ޏ���Q�xDG���ą���7�Y��	/K�r�Ww��9���r*��Xś����y��q��I��2O���F͙ĹKc�����G>������ǋ�⥗G���Q|�m#���̷�4��p:M(1��	ci�;��˩�������>N���\X�kQNE�8���QSOhc��1g�tm<鶚����j@&ϙp�Ѝs�ژǋ��d��va��Ǜ�y\Lb�s�ߐ���?_����-y�?���	�����1�Y�\O_�'�pf�n�'�ld.�M^�C��]���U����frώ�����\pᡩ{8s�&�k���2�Vy���e�}3:��K%�p�dh`,Cc���CkZ>y	Dy�� ��CBHq~�d������MJ�7	~">>��WY;�ڑh)�q��H%V��|L��4�@%4�W������z�q����^*��&6x�˹�I�
%�?\ʙ/�?W*T�(����:䋱)����Q�&�����x���}��N]�;%9{�h1�Ɗ�-2F�N���?N������0���Vs��!�>����ٳm7G����S�;rB[Wc8��9��}8~`��b��L)Je���6�o�<��ɹG�\�rF@�(�妎��v�^����@�77y��y',5�Sc���}U���= �V`�]�N����u�.�I����M�Q�����I�Aj#��L�dNU+b�Ȕd'F�f����K5{�NMj��!
�m!�L˴f[o_����H̈%��W�׷-���� �?���ө:~<� 7½���h~yb(??3��_�oO�w&��#�Ǔ���4~}<��?�ï���S���I��dmۿޛ�'ύ��S�y�1<~v"�=;������gf���d9������O�������I|��X=;�w���Fi�?zj8�<��]�s{0���������|xk0���W���ϻ���N?_��S�|s���V���"���%�<��ę�`��vcI�3��,�	�A��������X+��^uĘ�	*=^��>G�c�<<��ա����т�b�T�5sN��zR��P*A�(n��ƀ�%�k^%�? ����w�؁!��p�*�Q�� e�^�QR���8��}'NK}��k��O�������rNU^U���=� �zZqE��@M.�ZpM`P�Z�$�U3�\s7�{p�1��	�D�r���0���cccCFF��;�ׯ���6����� E�Qm�~�7�{��x&5q#P 06$�̸Hj��נݗӧ�P[��SY(�oK1͹I6qb��/�E�!pf��1i�z:9���LnQ�u��FMam%���8
H* �}8^��S1���r3{�2�0��C�Y2��c[�s`�LV�ªI�1o8��e��:�����ב[W-po��m��>��l_ώ��Q���-��ľYY �qZ�l+���zF���-0� ��I�����|U���-�+�ajR&A��Kf@H,���C�{e�nԹ�i���At�'���35����� 6l�Τ�3��x��%,X�G�zƆD�xjbO�����2�̚3�������͢�����b�Tj|J��-)6�1����Bkّ��E��-Y�vT{��72�J��#i��T�>�Ď|[w�Llɐ�f�]�;�&΄H]Jv��b-��:`&�d#�K\R2	��#$�__�l-02��K��~��
d���1F�s��9�% �e,���Y��+v,�"�_�\+%��2�ܞw
�<�S��M���3���vK���&*������?Z�j��o�z���0��QƦ��2@�r
B�M�36�K_OVo<ttqU"u�Nt���Y�t'���9kc���"$I@�0����d�T��S|��x7c�[��84!-��Nˎ�K���V]Y��M�����܉s)�<��ɣ�9��W�����)���(~�y��r�����G������T6����#{�}�#�o�y�R��'�}.E}1I��*�N��ʾ8�Vз��!�Zz�=gr���c����=�X�t垥w�H��a�uq*o؄q�:����x#"���=x�#�uA�0����|����{+���~���wx�P�$�Ը�|-�wE���8��������Ӗ�ƶ���?��U<5x�r[9a*Dj��E�v�'s�n8��1�>�9f��7�b�6�K��~���Q�$�GiP2���쩦\;G�\�Hp�$�كDO_��=��*
H�r
����9��碠�A���V�0���V��ܪ1IzR�Y�R�ㅖs��Is&�яt��Th�"��2�
�r$�Q�,���r��j`j�w��K����I�^��>���}�0� N���<�z7\d�T�Qr��KVq��N�?æ��ث�u;��#�8���6(�ԾC��۵}�uǞ�8t��'�p��u\8ʎ�&f99��@��tO�P�����/I�^f��:T����� �'O]2�خ�;g���
M�೻�yTK�y�������%o�@���x.wL�T�t�y'j���`��f�nW�'@�B<�N��(��g�cܙX��L?��화�J{�%a&=4 QjփѹV,�u��� m���ygy6����|}��oNV�s�t���/��׫p�?����L��f������"�l|�~�
?o�J�A*�&���m";DvI}٣-�y�,eԶ����&��d%~��O>Z�-?���|�x�����_χ����K��m|��9f5=Zʣ���%"�x��<>xW���9���@�sx���e�0����ȧON��E!�2��w��N�؛O��ա>ߗϛ��59��#�9:ďm���+s�o�(o{#���C����*���'9��A�bH����%܎2G��6�L��J���E���k���w����-0yLʖ�˖N\�N�Sȓ��·�p3Z+���ak�\x��m];q t8%��Oꆂ�����k��y�	���<&�s\ʳ�Pq���{ZsUϜ+�.I9V�w���놶y6�V����.�莩;u����5�����WL,�@�M'^}�fϜΨ���ަ���)ᦦ�r�{<ω��I�N�~R?<�I�QN�/�C1Me�V�j���.��������;j3����%'/Ɖs�c�������%����8[Y�eϞd���D�'����_hn�#�O�_'�� �1�*�=�g�0�6��jdǬ���0���3������5q�X�h]u�F��X%Y�X����]X�����^(p7���+8<5�c38�������O��%��,����vr!dVAJ)�g�s)$���(��O_gW�8z0�7�>N�tx�P+pV.�].pU`,�mcK�����[� �a��t�����6�z�}�!>ػ� 6Au7'�ّe�D� ���P��Jrl4�nNĤ&���VV�2k�Z�[1�0%+9��}Hu�cdK� o����.�ۻP'���̓
7Oʜݩt� ��F�}�õ��g?�<�i�
��P���\��ZW����v��-};~<�ǎ������\�y073"T�9A�y��j��-96���y����Q)�Z�I.`�g�H�SR��/��V����2_ :Gl����Ds2�ݩ�(�U����ѢQ(�Ely����{��oU��u-ϥ�j}�F���06�Z }��+г{�(�يnQ��ͤ�z�{���ꃇ�=���89b��u�چ'b��yB>6Y%���W�Y#�M���Sԯm�gS2m1	���=e2����:sSV�c�ɩ�xv*�|6�/�_��_��������~�]sS-ߡu�j��/%r`�U�8W�c_҈CaN�}�<�uC��kogȤQ�3��������g4�XqK�Us>oX��] OZ�s�*�[V�ܴг�9�h^����~��`�[ �����経�|�_|�{��P��y��?��=?}�##��**�gF���w9�1�>Ѽ��;�ps�FΗ�ݙkya�)vMZ���P1���~��eM@�"
9���NaLX
�<����t����Q����%J�C>h��� �M�p;��V�<�~�Z똰X|}quu�A(�N�m5�զ�1��D�[�k���ЩTW&blTxS̀��H�
!a!�Z͒�oFEWc"��I%���3,]�ӱ&Y�~���P�U����\O*E����h��߻E�V�v����u����@� y��=M$�:T��{�E/&�=*�/�P�/��32��+�q��U�=���'��'�^����=Y�s��n���K�=q�3'.p��my��mn���s����뜜:���mO鼭�/փ[*��(�uV�����Ƅ���)��M��5w.����[��ʮ�g��@�'�Ԭ�cRA�$�S�,Fvl�����\�Z�b�tvȹ����bx�	 ����MXb���4���;��C[�}���e��tgڂ�+�}R-{����FΌ���x�_��k�r�xG%_��#���f��~���������|s���{0�ߞ/p�X�n�x7t?*��+ua����O�ů�����w���Gj�~�}/�� ��~������"G��-<z��D�{g�#���=Zϻ����Vk����(��IE��o���W���[·�-��{�|��O>^&`��Ǐu��˺�}k1￾��_^�g�/�������ũ����x0�_��ӽ>|{��O����4�[���y�ܘ�ű	�����p���I�@���j��B��0�8��y�z��nN��-5�V,4�d� �j)˫���<)jƬ���A��.){z��S�����8#����7�=CY����s�r`%uA�:U�_ʹ�9�{��K��Ӻ[u-������{�W��*�JTڲ3"gu�4����dm�nY�;V��)Q�g`�#k-��=c��j�;���s��/3��XZ�A�W��ju�vq��ӓ��B-S�j�qpp"44���4<R���h�Ļ�1�f���^VT�3z�{���43�Ҕ(ZJ�ܻ���j(����>5%����=5�	�_�t�^6u`��5E�jb����\
��IHJ!1-���D�|}q��#+(�b����_?���6�-��-�J�ԒA��i������m�އC39�P֧ձ�2�v�w��ՙ{Pe&�Qt׀XG�����2zE�\R��Ž91�J��3�������)���dEH<��7�kn=dU�uQ�Bim�I��ɕGq���7:���L�k U�^��HY�Y��n�@��ow<�	�����ckl�ݴ��f֖������!��ѳY<e�&�����l�R�0�2���W��Ckն�"/����|R2���:�"��,3g
m��V�bkW���l\�r���͇r9��=%U�򛇯��� ���A���	H9h]���Kh�����cq�Ф�����4{gimOVv�֍l#��kmC���/�,�r�o#p&ϤA�8�5A�^�K��1�!�܆"y�r)�j<d�������3U�,�'���,q�T�]���T��[:77-�L�����!0�Z��T�B5/_ΡZC��S-��r�bkT+_�8�QR7��.� C3��|��4Qc�Tc��<�^:8�3��Nl���!+=l����:��ₓ�,���n\{�`,��1L�44��4,��qKI&�8������)(����v�Z��ځO��E��t�����G�i#�x*c��fȜ�ԍh�xp_R��<����*)Ǻ���:+�q��M`C#Y��0l�&�a��	������"mR�� ��yq�ޝ3�Λ�rK���]����@�/�؇�@��>^p���T.
����c0�]����G/�����_�����/����?����g��y�}����� omB6/LX̧���I�����|�%�ױ��!��l���#<y�9�>���v���Q�0ޞ��+]�1y�ƬaW�X�w�-��E>�ZړQz�t騖#�D��p�<M�Dq���'�#40���Xm�NZ`,�R����r��LW��6FX�� ��Q���E�T�t�5����@�\�~DK�sp'D<<5� Z
��c�*`�&���È"����������tǾ�+��5[V��p���V���� 18Cz��A*�q���9ϸ^=�(��b䍓kŽ(;�C�s��s�8q��ǮrZ`���9}���ns��-N�>�ûO�䃧�{�>W/��ֵ{ܹ�������k�<y����S����'�>a
�\�ga�IQ�7��4ua�y��'#�<� �x~R�����j�A�Uy�R�ϊ�8 Ǟ�;)�紼��R�O����( w�ȆM�I�4�+C���`���6�ꀼO��W�wP����Z�v�Q
������>|Wc�C��\nB�kF&X��Û'f��ֆ<m+�=|���o�*���o;�� x8Zdd�<��w��۽��h~{n"����_?Y���l����/����=���nM~�q;����_~�ί����ս��v�U��	���?���R��h���b�@�>~O@��|��J�>�`������R>{w5�~���������O�ؤEZ���5|��
>�����GK�ֿ>X)��d5��؏�0|S���">yq߿>��^��o�M◗��ó]|�p �\kᓓ5|v���wW��*^][Ɠs��1Kdo�0fd�Q�aL����ne9%Ϗ���ƠHs�|�ſ��F`N��RoW�s����P�K�,�v�|cbg����rb�(�u�}�
����R'_��5�Z�V!q�D����ex��[ʦ@Y���&�EQ&��v�q�T�ǿ 龜ji�nm��,8��B�<�</���{AD뮕�D�s��A�#����o�e����Oںi��X����#z�F ������J�*(���Ok-}[	
ȳպ¦��+��*��<w��5�=�_�%/���T����)P7�����5t5U�VSN���1�{%�y��S�(
�-�wtԺ��=tuc̘q�;����QZ]M��B�����"��πD�q�8�����	����z�ϫ��j�������Z�։el���_VFyq����-#�Z3��c��96��K��;7�#�*e��c�+88#��s�
8���)�L��AZ���Z�Q�ȉ�$Z��������=�N�N^t������%P��O�� �|�jq�K�[$Dg��烹�a߁CL�5���b�jVn؀[�?�Nv�8�1�ɖ,���諱f
�r�R�!�>Z ���?�-��}�Y�~�X���H�`��q仅�n���jGO*m\�{R Z)Ǖ:�}z(�S���^���c�\Un��O3)'�d%�k]�
JÂ�4�40��/f��Qd�c$���޹;T��m����-HS��'63�D��؉L=�?G���l�)���T�Q��LqZ��Y�&N�j�ӺlͥL�=L��!B_A�)�V$[X�e�@��1�������������t���΄I��ۡ��o�3�"����I�~��>>b����O�S�J�bG�E��.130�B������+�x� ��,=�0���@l�� $@ۿ@�ob�Y$��T��Kz
։��f�PX�CY-N�������JH�@|�;�D`�����Sܛ�>�h�we�%u؋ؕT�TQ�wM�ۇ��v
���N ������F�1=J�c�Hv���ț�Ʈ�r{L���|C�3� ��A�s�A<k��3���$u���d.�j�w�)�-�Al��'/���}�Wz��֝�����`��y?�?!���aژ�'�,�����'�[,���֘��n��s�yܴM�J�,�;�/����F�:��|`/�r�D.��̮A�X�ׇ��%�
Hc�<���#���#��4�]<�*#mƏ������73�{),��r2m}D)D��D�O4��Q�D����VR��U$�4�@��|�����x��)����ʮB���x1��� ����,���\�B��rY֊��ƽe[oQԍ��{�����W����g����a=�)�#�/�/JVA���L�s��3��˃��q��]����9%�w��.������0w��16�����{ٹ�(G�^����ܽ�,7o=����9�2��_��k��u���z�W�\d]U�	v����}��m���Z��{�o�����z��J�Zo뭍O�, ~Sޕj9*���N��S-4���O���s\9.�׶�n�ǥ��X���~1���ݩqU��ڪ%�ȟa_TG���u�6҇b�|�i�tgB�����jȞN?m�ٻ�
�|O5���C|~���O����~݀'@���po����[���z?~�%wÓ���%�7�Ç�������z�����@ߧk�B��oV�w+�k�������Vÿd�������w���Y���_.��G��쵙|��>xm6�:�ߚ'P6O��×g	�-����ݧ����u����Z~�z9�}��/�>yG���â&�?^���������܏_���M�ק�����������4��p_\�ϗ�D9�������d?���ī�Kynn&7F'��:����Y�w����־�,��3̒JoG��9h�Ee,Q��KX-��V��
��G�ս�䰾��=B��'��W,\	��T���fD�I=(eꤓ��8�[�r�� ^/+m�qs���#zR������N:q@�(��zvV�tzvC������)W�-�bh�)���<ih��F��p���~�#��|�x�+��^	����rH�]CĹ3���sSBY�b)+V/g��)�r��m��߁��)bDU��;ѩ<-J�#H��ڳ������^QL��R��2�W	��2����j���g�@�e�0>����t�L�IC����Z[3e��z���ݯ�͉s�8r�I�xژRam�"k��H����y�W���L/6Ϯa�26�)cלfv
��R���E�^���,��`wr��g�G�D^c6#ڎ�c3���;/��˪8��7�W�pxI1��{q:G6���?�R��.������nQ���уZ� �:�Pc6�9�N�@Z�}h}���K���NT�8Pd�Z�<�xrv���ͅ�s��}��KeC#k�l�꽻Dd&c�d���qnd8yh��I�T&%kYTK^Im-s/e٪��i�OJjŕuX�:���â�3(�"���[W��Q�K�,�LV�Y\e�ōo_j<ܩtsr���Q�L�_��ƙbq��J��)�{�pqֺ������
Zճ�>��������65�3�Vt�H��+.��Δ�MS]�N�-�r�O����,�s��"�H@N��t=���i�AAa��+9������c�Ιoj���{H6��i�ن3{�7Z�Q��5a�>��mx�4����)[jj��*0[� �YWG�n�S�����y��OtEzc�k���J�怕���v>��z`)��?.����������=��(_lc#1�M�4>��L,�,r�1�+�8���2,��+�ǣ����l|J��ω�"-��L�
��Ӓ54�`@� FT�11����5,	�`�k�L|�i��^}wvz���M�+/��y��O뫜هyOY����m�4y�.��d�͏��	:�vG?N����3�;��@�'�?��Gj����O����y�G�`FR�'.���9*��o&�'4���m\n���T�Dp!��7���ѫ�i㘅7���8m��d���Ξ�錑J=JV���x�����g�dQ�u�h�O��Ӧ_+O���k#C!�(��|)����ĳ�/?C��o$�ʁ(�����J���A�k����"�(T`K%ێC�Z��ؠbM(�!����qw݁�{	�uǻ�IwH���Z�:��ݵ����E���r���<cD���%o�x�ctu��xjl���Fn�=��+wپ����������k��s��u�/Y��Ci��F�x�EE����2s�2:������S/r��U.������8w�6����_��C{Y����!�xo�D9�gU-*[����Jz��C��Vعs�ҍ+�}n닑�B`���R�wF���
ylJ���9\����0vԺrO�4఼yG��5�Sq��
�ü�r4��ہ&;��3%R��}�/��í�|����v���n���"�|}���N�����qu ?�m�˿�5k�Ù&~:��o���@��.~�?��jl��s����"s���"�D&���S�]���W����V@^�$�&��s����I0j����#��뙱|v{4���7G���a<�7�����7F���������r�_ޘ	oςwf������i|�`:ݟ�G���S3��i���H%��G�	,�1�O����_�ħ/N��������������x��g��B�/���=�����ˋC�`O����E�����*?و��
μ�6�������p���֞m�N��B��r�ZH)j<�
���$��(�t�d�O;��JLK�=I��੉	*Æ�a�6t�U wz8J�r₞�6fE�̩.����k� O-UK�_3eUhq���R�%<%j��U~�	��q_�Y9�-1֯Xz�8�E�^	��\P$'dy  �}!lMbg\6s}�ɗk���b�bOtb4�֮`�qT�U��ч9�g1d�@,�	����ן�!,t��K�Q�ԛCC*�i/+�_U9�k+5�j��D��-/�,7���xZ�aZ#��ҹ���|y�h+g��|�>��6Ct�'�>m&��e�n��<J�@�ʀ�fm*���O(O�g0C`�F ~bY(��-�d��
��FvNo`Ǆ"���e��6��`V��=8��y�,����'���;F�qzY!��prM=g6�rfS3'��rxU!��rxcz��FF2���QF9�b�I��-��v��U�~��v	d�@_��>@��O �N �F��
;
��D�('7����=8���)�e6m�ɢ��پ{3,�7,K+s"�eߞ�V[.�`e�7efk-i�>�D%&��82-y���e´Y8�z���q�h�,��-@�����^�.��G�E�����C�,�Uk��@����2�Z�]�1�Ҡ��ɇҐh�"��qu���Xk	4t�6o!��#ۘ�"����W�k��&�98i����A���
�Rl�&]XQ��F��Y�����Ŗ�jV���T�R�S�!E�C �&��[��?�.Ċ�Zs�6�	#��=q���	JT�n������(� ����H�f����H9_�����@O���y�=u��)���,�Ϊ
F�T�U�#=YJ=��/6�P꿑����̰s�'0̝�+bbm�r$(��m��0F�����# �;�BH8z�aF�K|m9-YdԋP�HTNQi)�%����Eej!���0�3�f�1�gI/O����p��Sĕ��{�d] �E gLU�m/�<��yց�b������ξ�����(69�j�k7x���s ���
�H��G<��1����?�������?�_���ë�<�%e}yu�y���'ܝ��q5<S2�gV�5�8.
�{ ����'�h��Wp�Ɨ'���f��A;y����l�b�[ �� .�±H c���<�g�����x��AUH5.H$V��Ԕk��=��P�M�;��u:VT��_"�~��	)	X�Rh�$���7���*F�/I0Q�.�#�J�z�P!�U*�����ez�u�.�z)d���{��(�k��;D��b��6X�U��.���z:�����^:�8<�u��@�>HG_k��ӄQ�\���Wop��y������ٽ�$���Ƶ'X0oe�5$'��JBlQ�Y�G��EYq#˖l����x���~��N�����<s�O=��W_���q,2���?��"��jл��wW%bT��X��m]8c��]n�2�xR�@���N�������?^ oW/`�GG�S�,J��|#5v��w�܂e&�L��5�"���G�����9M��L�2�h��D�xW�6����u|����w��hk�m.��-�|������kc��[Ƿ{��jW%_�(�y|��H[��@�O���p��h�g�����T����ף��� �8<����#���î>|�U`r[o~�-���"}�~�{�?��χ:�a;�88�w64���J�yim����u�y{}���z�^'ϴ���t�۩��H��;_��'���ǲ�C�y|T ��P>??�����׆�����P����gw��݁||�����������A|w���/��K�xt��o���+���X_�.���m\��qq�-���[�w�)3���D�@��(�k��_�]�U��6��jB�J�f���(JNI=8&��yQN/����S�8���F��d�ee�x�7��x�=�[��)��cW���qC��U}+.�p'�3e��X��uʹm7D��%j8���-�� ��~�О�v�֓k
�]�{�̕��R���Z�8�9����i'��֓;b�y��1L*~���%v�N��SQ]*y CG�s`;��[IIO���_w'�m�gN=���)��c�CyJ��b7�w�,�5��,�כ��
-��
�R���^�ݡ_刅	�F��
��ީ1yj����f�p�
j���. �GZ\)>�Z�x�]��f�&�z%GTpvE#G�4qlV3'��sX:{�g��_˃)u6�hEQ{��@%�6��cL&�VWrnC-�wtry�`�nm���j��,����B�v��Jn:�S����pCZ��ks��ŋ)WU��4�:���J� r����`F{3B�j��}�\���m1ԇ�P K�]��% ��=36!%�����R⓱����ږd��Lsg��HX�5w ]��1-���8\����'@��G'o

*�*(��̴ٓ�M�����T�� hoSՊV/��`��w���/�"}T=Z���uq��ށ*G'
�Y��-ɷsG6����Ӳ	�}�d�oP0CF�b����5���O��ZXKKk\,,�ws%��L��^��݂Xi�ݪ�Z���'Jͬ)�z6 2��e��*eTm3�N`�q�n@�81*<N����&�nez��j��o��9�&�d
���ifɈ��n�21]�m��$;7��9��U�}+N�{�e�� �/T�y*���<'�*�_�g'6U��������X=c��&�g���Rb&��D��Wy�Unn+C]�-M�ԃ��*�
�A��ߠ<}���M��/�0��4$,���H*�i(���0�ּd:�3��F?�:��h�0� &X2�"��Fެ��d���M�8�Y ~�����m1u�Z��5	�y07ͼ�1yOY��p�6��l��v!�a�^���I�H6:�r�3��>�lG�ы���݇��������!�{~���}��uNL�̩!�xo�~8�"/�����C���L��p��7���\�����i�)����{�ؓ�����'/s���J{�-70т��e�P��^�2��@W���b+����{��i1v�4�$Cʌͩ��ݢgD��&�Z)tUr�R��y����TK��L)0�b����W5��K/9F�N�+�BS.K%���h��*E��xJj�*�Eo]����{��1Һ�{��W׈y�A��
t�)�!ʴS��S��U
`Q*�<��ȇ�*FE��.)�������9q�-;s��9Μ�őC���{�A-��x�i�ڀ���<2�K�Ϯ�$�����r�X<%�=�w�]���+�:]���m�|�^�w������Ō6'Qf欥��oJv���5�A� �j��Λ�s��17z�sU�U�ȩ�׿�k��mJ�N�l����$��R�*ǜ��xJ޻��f,56�у(�Gxh���hJ��!��]��7����Ѯb�<Z�G��x{Ko��0��e9��4������,^Y�ë�syky1/����i�ܝ�ȹ�p�����8.���ָxn�����(.�����.�6���R�l�J���4.L���4���r�)���!i�xk��g�H�l��ܠt.�1�R950���S��Ú�VW��̟��bCe0�k���)[kB�����x���ќ��̀$�I���N�����l�O.���"n�,���"�^V�sk�xe[���5�7��ޑzk�b�}��m��}y�l;�/���N���d_Ⱦ��yo�FD2�Pi��]��MK������䐅���	{rH��:�/���Yʅ�����W�Dq�$���K���Λ�cOM��)e���?��D�'��\�-e䚡86��ⶡWu-��nU]�ݓ)̹�o��n�-��[���%�um���B��������Ӓ;��+��{ň���r�HJ�l�ֳ�����rW� ��&Z/������n����N|R<A�A$�%������'b\\���ٚ�ꌷ���(�����8��kcTk_F��0��Q[*��[ZB}ny��%�hAۓT��T-(�����!��ĐWP�u�VgWw-�hQY�@I�>A�y�s����RwՐ�X&TD�kl>{��qhv	;�+)cˈL6�e}{��'3�!�tWS2��(sK!�:� }CzGزgJ	75qfS#���ܶ!�����-�Y�[��ӛ�9:)�c9I\�*a��M�.�d�{ C��d17?����LH�CW`�8xI̎Ig���IA͸�M�=&�!9ET&�bgcMtR���e؈Q��;S���#N�rr�����qbt�*k<����6n���� �(NN�����j���JeUy����[�{,dь�T����K��S(�\ ��38�����/�c��Ѵ�JF��0&%��Q�Z�j�k�8���Y@�#E�!/�1�4d��)`���HFn.�W��r��N][?s�P�t���Ɔ(g*�"�	�gq��I�cWo�k<Tw�=e����S,�X�ZZ�{�����۲�]���m�FΕCg�
(�ٷl���Q��ήe�r�G6�(&��p�N�ϵ�سb#;Wl`Ϻ��݌����*o�jT���	��j�S���k]z	�(�s��K�<��V��o"u�B�uO#m���՝�2 )Q-~RO�d����j�J���D+��H8�w�'�6�X�`�l|��.�3�<�V��F��3�n�4�X��hO� y3)�.��qa��+�t��m��
S/֛��V����Ft�
q$�K=S��C�w�8���9���Y�{q���{FnZN��-�x�܏W�xS����/<#�$J�IP��~x���7����G������_��k����k��8�uq� b�9��̩����ͰB��n��V^����|�r��(b�y?���y�܇��)����;z���������,�}������5�zZ���X L�`�H�b \���k3�T��}�J�d�@_CcjB�t�-
�^��F����bX��")(J
{���A�j)RaN�K��LΡҮȺ
j�D�_&�
)D*�E��%����y�`�%�Qxa���pCĀd�i��|���R�*�J�}U�832����C��{0j0�;���~�:��αU*����9|�$ǎ��̉s�8z���ZLTIQ�	�Ѥ�$N�)q�5���s$9i�t4��3���3<}�w�R?�x�����S��ڭ�̨lfO�`�^���{N3o�T"�}�@���G��]_�lQ�lܵ�a��]_�/FX�����p��F5>�l;-���|���Zw�ݡs�1l!˼S��. pQD�������D�.�Ճ�PW"})t2�0e��$^^Y�g�+��X_><���;�y~m<O/J�ɹ�ܟ����ܞōI\�ņ;������2+�C(>"΅�7�z�7҉��T�P`Ey��~�T��S�c��	,��!�[��V3t*�m��Yr��f��f%��F�B/;
���v7%�Ӟtk�̉�7%��D[&;���`)�R���u%N6��Yr�</k�]m(sw��ˁ2o����p�>ܕ>�n��azn(�ʢ�n�M�b�噏����D�N�������++
��Ώ�T��`i䫣|ud l��-|z���7Vh1��{3-ۅ�p{Z"�i�u�I�{��g�ݥ,Xjݥg�T�a{�@��f�,����/�㙮oC�|[��L�4RC02���e�\`"�9�'w��4��(�[g�V�׳���9�U˫=M���jy_@PmBφ�rJ�X�P O��r�Rǆ���h䤭+yN���☞u�K�O�2�o�u����m�'b��8�Mb�}��qB^Vvb���f��y,^�����hc�6n����s���"��IsTk��2z4I�	�+��nGkI��*�kfp}oM�5Ч����,�R����!7"Z�3�ڇ�g�6"����&0��ၻ��&LbѢ%�Y���[�3k�Bv��O������Ζ1����	��Saaʐo�NfӸ�O�c��N(f�t��c~G(ۢ�n�<&5�eݸ�T�Eg(���!�rtU={�Tpj� �l�]\��ŉ�m��!����y#2���w�c�t
�}h������Q��\��w�����Y,*-gVV6Ó����\��"!�z/&��y�Dq#(�K����Ik�1j�w������p�CgN���-~��^�6$ۺ1�o'k���&+d�!nIͤ<-g{;r�:Z���g �;���>�
�6)��Y��?���M�ۼK�)��e��ļ2��aYK?�͒���W���2�E&R! �,���M�S\Ș�޴W�k�_��������h%�6$:Oo_��\��=�X��8^��ֹ��>P�ğz�Z�C�q�5*j&m��M������L*��}�%���&ϣozE�q�4�������Y2O��+�1k�tr<b�
�bT�`ɮ�{�;e�\dR�$(O.`���������Ԓ$m�^����y�Ro��<xu�j"��M�
���ޫؙJTH'�mk)�E��o�I���b�X�1
=囨� *�L��!���d��)-1��H�R��Rq+���m����'L�C�Sì����%�f��c�,�,l�D�=�c�Tq<�TA�߬��$�r��{��9pN�ʨsU�sE�}]�;z�<����޼n�ǻ���o��f!|f�Ϟq�[���4v��=��jq�6ȣ�_����;��y������Pk|�ۏ|�ϯx��eΌ�)4�uY+
�C���M /��SO�s_<��\��!�m1�O�p�*�sB�'��9m��q�P���wa�(���,бe��=��(�S��"ޫ�מz�E�[hA3�-���+РZʚuu�5֡�T_kU�𨒏�䕉"VR*Rܫ'�=�7"���:�5��K�Y&�G���G��"�M��@>b��+!�x���ꘄ�c<��	8���� ��G��N�] ���D�R�3ir|�>Պ��U�����1p�s��HoQ���]���W�q�)QP�9v��N]�&R,]��v�7�0��;��")%��P���7#U���Zb#�II�b�ҵ����<��<q�O^�˥�7x���y����0q6S���7}O��Ū�[��Ѻ���A�,04b���M��,��<��z���祠���~F����׫"�����s�>b�@^��{1�z�9#�謱ˌ�[�D�C�h��ԩ'��yn}_�q��O�W���><���[�x~U�f�sgj�T+ݘ��gK[+���aM�p��l(q6$�J�k#b�	5Cn(ޣ�>�����sZK����D��/�Ay�j,�Jkg(
D�?�7�2d.�H[��}�D騥�My��%Q��T:%z�f*Ϯ�w����lS���c8��{V����WyWV���Z�T�jo#}Q���Y�agJ��1�n���`X�=������,O�Vr�3����e���2>���G�{���:^[_�k�kx{[�l.㥅�\��U��ǚz/GQ���.��Ϊ�&Z:��fܓ�R��tO46���.��U-x���z:���4G���ˀd�5w��h�l�S
Pu���*|�&���H��!׼&��/y(0���5O��~R�����<-p��(�g��b��+�N��cǛ�l���]1b+��D�[�hn��U�e͌>D�;�0$A@p�NFv�IA�-���kS�,h�]C�F�w�ᄇҷ������M���ڊIcFr��1JR���oc@c^�Kh).��8���2�T�R��BzD	�~�F��"eօ��f���-�KO�t;���h��KKKaɢlٴ�M�6�k�^������Ft���6��R�i�M��S#d��kf5�������x�����^�zz3��_�˷Vqa��fS���=�y��CZ�����
����.����g������sG������y���y^{vo���u+�Q��;/��գǈ��gxVg�/b}�1�J�ad~#��ٚ>T-]������_	��z����������_T�e��
%��'K�eegP][OYm-��'�c�,���H�����v�ㅓ�ٱ*Hq��]�8���6DE�w	պM���p�p�/���:����g��k��7��˙��D��jc����'!�b�H
�bHt����y�����倬<F��Ӗ�Ċ��l�5�э����Huz
�n���Z��Dg{�;�;:`)�ZkU`dwї�޼���_��R/G�@�|�㩆V�������EKS�f����V����̓/ʷ( s!HꝊTq��-Μ�Ĭi8��4y1���0t�(��K'o��os��5���CZX
�R'��9���Փ���+�E_��΅Dkg-3���7P���"L�ɳ[h0�g���9�SXe�P1T��/��t��1�6vx:��f�IV!U̅,��03q���C3',,\�7���2�O��g���%�c���j���e�F��|�-
�G��\�1���]F�.�3�`��]fJ<*�j��3�乔�6wb��xG&�}�6we����,������؃}r�c�>\�
䢥/�D,|�"�x�"�6a<g�k�����;�q|�˿��!��b39��1���E�m�`-���l�����)��C%�������~��=�ɉ������v#KvY:s����=���-��-}x�#��RJ����A�6�G�q\ �bX*�<ψ�?��N��I\���r{/-��j�@�Xz2A��FSGR僩3��
����< \��ٍ>vN��r�ZאZ)�u��T���R@�R��
=cʤpT��?�T
P���&�R�*�d!p�,�Z%Ǩ�_��h]�"�"1b�s�u�9��X`g���wz^U���1}�Jz��k���C��E�&i箅cQТb��q���FZ����}��B��#Ļ���e����]�t�iN\}����f��S�=t��w�f��U�Gd�ӈ_fN)��4�V\CAI%eM��������(�M_��g^��^���'�t�2�o?������[���ae��>���K�/^��W�OQjn�Q�{>" ����x����%����
�.i�s�Z�e��<�91�{BSxf�"n�Z�A�KWn��*��E�+r��RIvH���c��z�jFs�S
|9<��wu���>�����6���\^\��3�ӹ?5��C"��'L˵:8ɝ�@{��M��5�ǸfD�Z�og�����<��I[G�鯼�=�{���.j{Oy�I�:�/Q��-J�}��]z�yu�MԹt����5��[YA��j}��ʐ0Z'�=��sfP�c��YX�́~�ܘ��k+������Ē$�Y����yqY*w��qm|*���h���R�I�Vl���bƝ��|�k�jf��&U<�K�^p3�^+��1Ժq��ޕ7=�ځ'���/����yE�K��>�i�-���&��5��(e�Q����Z��zWD�
L^�i�u�>�X��=�k#pi�S�Dz�<�<�a�C]K^��y�ԕ����Ə�#�Yj�LCOs��]��Y����#y�Yʛ�<�U������/0|����g���4;�Û��N#35����Ji�͢�9���B����1g�N���MIl.�x9��ʍcd�jf���yټf>[7.gk:S���"���T2�´�k�N�غmDz��"NV������Đ�KNf<~�΄����DXH �����B��"?$D3�#;��"�q����U��[��׷��&�6��������������ə�K��f˒��|��ҵ�y�\;�Q��W��˧r�w|��y��K����r������bU����#��iq;�.Y�u�M��ɏo}�-�m�T'�ӧ/�z�1�����j�ԷR�[AC^%��ٴ��~��'�Eeh]u̜7��#���BS����n���T�C#���(/�%-ԗ0'[����뷞���^!Ll�[#�yi��%��GEu�}K��VFSK9�鴴��r�7��n>��+w122��%�������Jrs�L�!, ���T���)I)�*���ͭt6�ѯ���K��Ԋ�VƤg��?6�X�뙲t�b��a��8���3�L��Z���s� *�ĭW�<u>Q��{Pg�E�ؘ� J����E�����k�m����䩛�0c�
2�*HJ�c��Y<}�)�\Jrp���<"�	��S���m��u�$S/�ą��=Gm� �$6�����ǯА_�3�t$��U��5��k��"{Y&�Y���P��#��3ɶ�}��m۶m't:�4�L;m۶m۶mk<�c[�zWU:}f�<�y~�矙o��v����Z[A��y`��{P.��3��y���1X;�Clj.�iE�D�����[4�Y���bX�i`,C�����nx���ݳ�:��x䊲���!�;�P��ܳH�L#�3��b\�H�s�|�I��S��Cn`)MBʩ*��=�*�xZ:G��1�n�	�pK���|\b��0�xF�&0�/�1�LvKe�{*��RX��:�"6��-����y�(�hlGBs��X���|���q9*�W�|�Д{�	q��k4��Y_ۅ/�����z�6����S�������_~�����߳k�<X/���܎^����WN>���P^䣾��n�n>Y���������<������sc�,��ObO���4��u}Yݺ��-z��Ig&��2(����h�[CMQK���������(��>�	}2K�%��3���������cL*�Sh�DۈDj���e�٧(,�6!	oT/�a�,�RL��_�:�F3� ���I��W{8e�Q�D��/}ӨK�')�k�&h<�D�h\K�8�zs4�躕`핇�$ZD@*���j���h�`�}�M�TOe�{0�K�2(U,M�-��-�.�˰���v��瞰j�Yf���(��!���z�Y�o?BہS�j9���s��OnGbj�mZGNig*[$+��^)dH��]��3�p����8Ͼ�G9r�"��
������ �2����S�4m�:n������CK'EF���ᶩ��!O
�r�qy�'T�3Ta��;':"p�)"�ۃgpn�Lf�&���#R�+��x�.;�sת�Ċ]�Ěwa|yۆs{u7�j����Ʊ>Q\���Il�gz��"�)����2��^C�{m],R��l�����cC}uvme*;]]4�ʔv
��/R����z#e������������ߤ��"y�2��<S��OO VY}IC��`K�]��v���Ì�p;';��e{zGs}z67f�qaRצ%rmr
�Ƨqut:[;�00=��n6��6g��%'�k��#R��]��zd����$&Y��,i�+q読���t<A,��a<s⾁R}��#SO��rGǞs���߄e7u�� ��$�wE@O�e6EJ�uW�7���Y�P ���#EV<ֶ�CwiY��H �SKo^ɳ>���1F��96��f�F�X�c��yM�C������t�7���݇X4j]��if��Ծ��8���~|�O>}ȫ�����������g���>o����!}p��~��9�aE!᪇<+ԇճ����9��������>?~�!?���ߊ���=n�8��ɣ���pd�:���F���:5c�N���'�}�4Gmg�Y,�?K����у=qH�͡"!���p���I�ꎸkooæc������|��#���_|����~%������dFD2s�L��C���:.�Å�����W_��?��O���/�|~W���O>����Glٰ�vU�o�n��=|h�Մ���r����N ��������������wx��s�<��1��خ+������u|��$�Zv�oT
��{���~��3��{~�����+��Vֿ�����O?�D��y~
ݻ7����c;R���}ؼa;6����}\�r������'��ÇRx�����4��c�����jS�mU��4~
�f�����{�-[�y�~Vm�ʢkզ7+��f��a��rul�:�N�λs7r�� �'gsp�~��K~�ׯ|���|�����[|��+�����_���*�^5��Iy���������Z�:�pʭ�թ6k�l���Ak'��0֧��#GN��O9��������g��r�,�#�ɗr)F~s=�K�1{w�G�͑25�n5�x���Rf�D���26frۮ��u�A�eȷ��Ė�b@5�2��P�3��B�B�j��3�8Go"��ȋJ$)&;�hl²�����=��|������|�}�q��' �)I�D5�x�zV�����h�E/b8���1���Y�h\���6��FV<���)D5�Dt�8b���1������B2��3���ᢑ��!<{�9#I�Lb|w�c;�݁����t�,ZQG*��S�ԙ�)]h�ѕY��e��k�@���;0���W�18g"#
�0��\f��ς�Y�}.G,��Ը<���/���f}x��q.�%�J�rc�.|r��@^#��W��Q�)�|t�{w��b�
yy>���ϧ�޼4��rX��.���'<?}��Goqr�e��9˦EX1o?c�n�װ����ÖѢ�L��M�H %�p ���H(�'��A���j҃&M{QUݛҲ�4 ,.�������%;�yY5�W��֔̔r��Ϭy�Be�&�D�zin-%���mŒ��_eڤ7#=,�����  ��IDAT���mݛ�����kAeF3j��P�ݞ��6XxW�q)G�\��s���h9����#�&غ��!�OH?Rh>?��v��)�iJ�P���1��a�f��WJ�-�i��As#*|3�o=���61e�>&�����5q!��l��ɳ,۴����H�)��މ���Hdawɜ]��FtN=�Ø4�0ǯ~��38q���?���;�?s�C�s��Ox�i?�<C9c��.��2s;	��*�)�jJ/B������i��3/�<s�!�� O�(=gO��y)Џ���-2��C�pa�lf$s����'O�cZ&��Oi\���Z�A�&�s0�e�+cJ�Y׫�ӓ;rtD�:Ų����,�
cB�/�!���t$��_=]uh��jT���L[��������9a-:e�}]Lt<zF�җ�Qʤ�Z�^{��'���O/\�����۵*��� �u��`m�r�z?9O��ă�����&�F̵��֡��)��X�ڟ��#96<��c�<&����8?4��c[BgwkFI��Ҋ��֪�N��c��
�ݶp�o��]Tϵ��_G_���8�Ȗ��)|"��D�R{�Ȟ�R�3�S�X��pQې���H�'�{b<<��+�/�T� @�P��ƌ'Z���1�m)D>0��=+>�o��{�k��Tc�G��|f��g:�|m��7��<	M�N�`�m�@[3{NF&�<=�%.~��c˚�L>\���S�64��b�=:s���Y���?����6|P��C�Q���)p��/^$��Um�ul�6�G��mLAD����4ܾ~�ӧ�q��N9ȥ�'y|�On^�����5�t� &t���]��ut�M~[K�N�o���ߔ�����;�%��_���j�>�|�Z�.`����t�[�V���P��o	�~�!����珮���u�yr�Wo?�ٓ�<��E�Ƒ����x|�m��I6�$�Ã��k�.b�ҵ,���%��3w�8f��~۳7�:Ҽ����R��̒IS�	Vn-F�����C�D�O���R}�'��+���G���Β�޺�k3����}��̴��]?|�69j�ǿ�HSڙ�)Ѣ��Ґ,L�_�Hs`�@聳T�Q��ǟ�m�*�كܹ|�����m.�<*�q�G��0~���ҩM��ɓ���n�J�w`�ȉ|�޻�"i����?�?�����/����>��c�N2m�TF���N�0p��^���C����p@����:q��O�g�1uԝ[�n�6���Ī�h�[IJ@{�f���4q���[�Y��^��l��ⳤR�q#(�S��l�N����|t�{'��ֈ)���(/��a^Q;����V\K[sn�,�����[��۸jnKٶ%�-_n8ƃ�S����X.yE��kO�����V��z{m���.)7;���7�-u8(�ءY�[h�^Ffb)V>��K�Z*�kS|Z����v�:��J0t/���	�^Ͱh��{s4�-�xwA�M�P�b&��8G�N�\,�V`���A�n[���uؗ�Q�-2�c������.�4{�*Ì���0mF)�1M��y�\�2�`�>K�U�,lrb��X]Z�.ľh	��+pi���584_�C�f�Zmƹ����ülvM����8�]����6�}��?��v�`��[�;|���ss�at��B�yr�3�u�	��V�{�o�'������Me��W7/q�ow��x�ͯ7w⸓?��/�ݹU �2No�Ė��X��4��]b̒��y��3�Q>�IC�>� ��v��f���B,��c�;ۂ)��N�2m�q}0��]Bo|�x�������&t�&�3)=T)���q��cL[��`��ĺ7rO��%���mT)�nq��,���s����Ӈ����Ĵ'�x0Q9�K�DDb��[�T��O�X�vMѲ)D�.�|t��%ҳ/��>k��-"q���;���J��	v	��ș��sh#�*�hmN�8��I1��6��glc���Lț9w5s�R�]�~'S�m�U�1dv"N`1$����4�<��V#i�f�d��{�����c��3�ʗ.��Щ��9}��O��ʚ��ㄭ?{;O`��*�)�<�|� O��)�w����<�@�����ŽasUț��z����F�;(�]��u����4
�yXS�L��0&7MeA�,�(�x$�1�؟	�����݌,Ksu�&���~M��Td, d����gkS<,q47���GcCuV[�7��(�F)���]�75V�*���V����?��ku�ߥ \#�(�y TU=B#yWygn�up1�U���,�ih��,{��`W�H��K�P�vtbMm ���m�{K���qY
��Z��0�咾%wl�o�#FC�:��2T�Ҡ:X�@��B��矠�{��Q�ΜK��j~����Ӷ�\wU���� �綾|`ᮮ+լo���R�\-<x�ʓ�mD��|h���n|h����>�p�3w��W�0~r��[�P>3��_	Gp�}�i)y6SϚ�1]-y�1sj%�C܃�9�������=�=�C^1̷�a��y�>w�M;ws��9N>��C�p�:���3��0	1.>�Pϓc��Z$�1v�d��GBD��&م�.��eqSڔTQ�[H��L2����bńiزC
��Ԍ�c����wyt�)���y��/?��g���y��'|���|�֧�)mA�[(����_mO��w�heCilc{�bl�ތ�YO��m�Y�F���iמA]�ҫM[rB#H ڻ|Řo�@��y�^�S��LeN�Zp�D'S��NuJ6]�R��CVpQ�Tg����}VN�A���:J��fj<}��G|��7Rp}�;�|�G���׿��W�|�?|��={Ҽ5�GM�u��ڪ�%�NL�­Gؿe�������?q��.r��5u��#��/�aX�j�����pM��6"�2??���i]]AmE%-���!09�[o��jOMIS�S�)ɑ�hVCbP������W�7�9����}���E`[)C�P�R`��_Uؒ�:��\��,�:��U-9Ҷ'�4�jڙYɹ�iBef9�	���f��T@Zr��9$Dg����w(ޞ�x�8S����W�3q�
y���S��+�w8:�Wɥ�S̯��|�ǗqYܗ4�l�^�;��ڎ\�*��ֽ�:q�k�� �:�ם�x�v������!����Zs��p��x5u9�br�6��ǁ������s/�]y�+���!ܴ�Tۛ����PP
����G�6S�!�?�v��)J���+C�J�hsl�J۵����]3t][���L���X��z{�����M o ��Qh��B;y!�i��$.A�h�XQ�k%-oP��ǯ�c�V���s�e=u�[$��ʺr�|9O�"Ǔ��R�\�*J_ӠQ���hr֡)؄�h3�|YnA�DT�M��/���hZ^AS�M��h���q�K���>G�����_��/q��hE�rA�e\Y�Ȧ�����}�����yb�I�l��FO��>�X���F{��ys�)�w܂y%�3sO��qe�|no�̚a+Y<a+w=b��g�:����n�2����b��6�/a�tE;�/َq����Ģp�y��M_.�������(o	���J��J[H���O��a�L����e���<i:Vr�e�,��&c=���`�4��)X$�G/v��O���^�1K�QpO�l�$cI�h��m):VZ`*օ�&������S�1�F�(}�(4�����d@��?�v����Й���4�r��I8}��	��.�)%�n۟���Q^ڕ��z:���_��L���b	͛����&2m�,.X��}�9�Lyv�w�����\>|�#K�^ڟ>�=8���ڳv��3�~���<��Q[?�t����������k_�4��Y+յ��0;�m�B�s'.Nj�ɺ�f���gl�&�Mތ7��#R�5B�2��69���ԞLJu���)���ώ�Gr���dG}�=���q��Ռke�=�:�BK OK�i�P�#�Q:8(0ckn���1�fF8Y��im������Y�]�������@��Y��a�������PGO}n#t�
X��r%��=ޔ�߼��3֕��"���ĩ"e[]W:��b���z����0��H��$����%�������
���Ŭ�6v�bS�@6t�gn�;�S\��HW{u����CC+�.j����ޏ[!)ղ$J��m��I�b`���t~t��#{�57$��X8p�ʅ[Y�5���v���w,�y��;q���s�8�����'���Q��[A����;a��HQ�~H&o��~1&>��������s�,��K�o���q\�fY,u�R�2Mی@	g7s{^�'p��U򢆁��*��p���{�p�l.�f2U�N�5;��"I�Ϡ0����4���+�ʣ"��ܨ*R���f�o$O�\�sbW9�>�ɽ�=H	��8*�R)��'�S�SI�*Z��&3�֙٤���p�.��xy�×�o�]^k�4����L�>��×1��D����W�~�2�!��Q�I�$)��ݧ�z"�7�f��0��O E1�Te(õ������V�[L��b�F��!�K�����=z�b� 2��T�NUv,ٱA���g�УE5�[��Kq	�*[��S]Cu��E�y��s�Wh��%U�!mY��s���U�诿��W?��P��xDE���gnݽΨ��92a=ˑ�Zfeg3���:�"������)˫�������(ȩ�IAK�C����:>������{t�M�Y@ �Ԙh��H	�UakX���hӍ��\�R�ԩ4�Cc�H/bV�0~8|�/'�`wI;6�ͻo=�0�*a���������F�})z��7�X�����8�k?����ul�ԆY�ړ��@Xl<��^����{)#'DG����#��~Ĺ��!�\m[�x�<�����F�	�@�Ǥ�eF3~������o��V�@<����f���sl�ЕO��x/2�/W��ƶ�,�ޓk+�����\�x�-��Y�U���*�N���)+94~1O�cGρ�q�`~�$>������&\2S;��樑'�ͽ�Q6�Equ�D��ǀ�2ں�2$�%-S�qt�Rk�][a��^����]Z5ȵ��
m�����@�i;֠���:4��򆣗4��q�J�/H�mE��k�Q�
��Y�}�U8T��1f˹SE3Ѥ�C;C�1M�/M�/]�S���_�@^�ke�e�- ��+9 �wM��h���N�m"�<d���Xz�m�x�擟rq�Y�6ǋ��\��s,k|�94`���/>h����נ�@�O�OP��k��׻�@��ZU�Q��#N��%���x*	w?���#�pu�Q���f�������G�b�����cB�\E��%45�E��.=�v�qy٣薜���F�'�͕��܎&w�k	�fn��ΐ�_�.��(M�;e:I����DſH?y%)�%�W���H"��$x�L�D��$ɾdQ�I�Y�If�6-��h:�5Gת#�r����s�X���E�����U:�D4�qh̒�览�2
��<�$����s��X�`�`�,����h�2�l2�XI��n��3��CV�k�*FM�����X�b'۷���K\�t�k�op���;���u�d��[l_���9=I0��*$��;����ϸ��	g�=�آU��C�
y�g5T��i�����4x�޵
��2�@�o��.�,u�(�_!���Yo ﬀ�yGtM�+�',m�bbI_YW OiT^�G��P�|])s��[������LS7+u� e~C��!�����ӕ�F��JK�kKS���-Mp��v����)�<l��&�\��UT�O�:Y��r�4P4���T�2���P�I� *˿�@��7��|S=e
?�KCC,���1���$<��f�e"�7Q�uT:�(KU���*a7�{��bi�z2���1�p+��ĕ���Z�m/��1�W�X��n�k��/��b� ��B��9��˒Z;��ګ�koXqM߂Kr�}-^���*��X����~�Xx#l\x�;��x�H@�Іkb,(��ַᙉ+���y�!�۞��#r��3��a`�t#;f�80�ԑy��̵pV5O��16����Zl��R1D��H�m+�=Yg+筰d�m ����,��"����10'A�c���� �O�d�@�xmK[x�+�����Ҩ�ܭ�Ȗ�\"��pru �3��p��0
��i.��MQx*����n�L��tR���u�
=S��$�4�u-��u�ez�Y�u�tʮ�KV���]^��=X7sv���N}y~�2��l�B�G���M�b|�,�����.��'��Mn��%1�[��
xy��k{�k̀�2���B��&t.mƐ6u��nEϊ*:	(�P�o�+�6���*ټp�]zD�2m��;��Oa���tiUFmi.-�rۧ;sGQ�q��T����h�DZ	��{�![��&�Ά��@N�Zăk�y��>�~�.���!�1?� t�g�7L�}��G,3��c�����m׉���Y;�/�YUeU�d�p�R%Pҩe;:�zw�EmY[�����6]�:�f�w��;�!�%�^��Y��Ѷ����Lj�Z������Ѯ�MR��ZӁ��0o�X�>~�G�泡i�N�̝�x��[|��s�U��W�r�;����է���[8u%}�j��e4/�`���N�o�\�ϜB�ԧ]�;�n�v�ȋO�(-�����~�RF�v�"2�Kǯ�x�"*%t��Q��z�R̗bT}bć־�k�ͻ<t��NH�;��_o=�L��b�$p�:�������xy��N]���=뷄�ⳕ�y�n?����~��Z��i�x�v+�[t����\��Ui-9��U�({s@~���9d��1;�9�p�~�����K:}���ՒVyN�
�5��@��K���t�O��[s՛���\�-ǖz�Eǫ#��h�GHy?G O)��DzR��U:wz�+�M[����N��ר��N��&U�.U�.u���tt3g��5�la�T�,�S�|��"�����r�Zt2׫��ڀq�fL36c��	��M�����hf%G1ir�ꛘ�{�Y�;$�}ĺ�_��������{?��3�)ϳ�j.Xq�-�>q�(���G���W�����
{�<�����I�x�޵s��݅�>~�5sd��7��x)��b<1��^d/ƭ�Ҍ},�����X���>e��g�����.�izF�U��
:����:�V�1��aP|���tB����� �&������d�`������A�䖿�n�
�e�^�Jtb�5�
Ľ�yѳ��XΕ�
5q�� a!:���q��]���гj&���Vh�4E�4-��7Ҷ�F�&=�<u�e&�'�gn��K&~nex;��f���}&�9���ܛ�QN�W3�;RX���3�2b�mz�=���g���6�w�b��S,Zs�ek��y��o�����Y�xK�a�����I����X����;|t��P�o|��7ܓ���9�8����X;e#IQ8J��+
xpy;�|�#��y��y�ܷ��ޏ�
�)��;!��C�ǭ�L����~K�5�ۓ�P�MIv4�.֛>	�T9SbcB���Z��T���j��h����zR_ �P3!;;;�l�\�mqw����7gk����&?w;+]�LQ����5����?�m���Nv�X����R��7��|sc0���q��Tâ���Q­�^�����
�z)�jg������;s\�%����x��l��v���-]�<݆�2��2�t6p7`W�4�X��6̉9��qdp�-=���� �����l�q漾97����<�2�g���WψH�O��I�@�@k{��򾅷
t�nh��@ߚK޷��s��x-ߚ3�M�r��+	-�$��G�R�V�݋%��d_�r\��d�ْ)ʗ�jc{��[R`l���_edKS-+�	@�ZSlh�z��L-Ԟ����#��6��w�y;:��U]���e�ǘ�|6�af����Ђ���tmRL��l:ee3����C�n�Dn���}Ϭ^��^��6즓���6���fR�zz6��}n5I�H�`pm{�N�ę�x��S���O웷�%�Fsr��ͬT�9�j9�G��SA�$��-#�~��t�ˢMN��3ѯ;���fv�nt����փt)o�6qX�_<z��EK���:���5�7)�}N&S��3~p��[ȽK'߷/�������Ԙ����>���~������Le��!��Z�����h�\��ͧ�É�{h�Y�'�g�u �N�	�% ���y��Z�ʑ3X9x:kF�ub�*P����|��w|��mƉ�ca�.n	�-q���:���FӾeK�
��ݩ=#%������}�6t_��%��^��[Ql�Ƽ����\�̔���ޢ����ש���;��W��4�Cwүc���k��{$�C��ٮ��kX�ۧ��ə�<����N�p������cX8f�z�د`i��:�>�Yt����=<=�	�1�m;�nCˬ"�U�Uÿe�*ɗ?`Nǡ�eq��fL\L�{$ͼ8U���MyO���n��^��Yw�ň�n�����ɇ�������\���RR9_�]���wp��n&�q­�s�m�e�F���{U#����p�E�n���Պz�V��"�C�>0qb��%����m��{@c�	ӱ1�X;v.u�9t��fPN�m\�v����z��^Wٺ�C�)K�Vh<Z��S�ie��oG����	�&r<i�U���S���	|)2�m��c��^�ä��'�G7y=�)
OHٯx��]��\�|�K�`\������Ehg-C;SX"kU��N��m���henm�����)��S q7�٢�=���&�g1jr���{�~�'č{��3_���;L;��d�3�wK��8��s.�\r�f�̇�}��X���߫�-�~��7��_!�����z��)v�wb��/�M�Yc��A� �	��g��Cc/������\���ee��:x7���˒c�������.=�*.�] �zy��N��>�n�QY
�o�['�t)��+Њ_�Q�D�,��t�N}�����i%����k�~� c�wKЍ�{��^��x���*jEJ&���������a0��mmѵh�Ƹm�XK�3�G�8]�L�L���w������c�[�SXk\º�2
��Ixe��5�/�)�J�]\?\�&�^���xWoĵ�\��[����E�V�&�r�-f�[;����d�����$�+���ӝ�����&4�Iѭ�.�se'�]��*���?���sq�;�#R8�����H�P=;�pj�H��|}���7h�@^�@�g��a�Cs�e���;�#�U��20"�ˍl7����U��
y�ڤ��.�`/�H�4t=�����.�&��[bcc���3����;�ce��;��g'�<7g|�"O'�\�Ȳ5�2���_G+�m�&_�Go�T(����ܬ�����|��v
�)��l��˿����ZNjG� ��t���	W���۫�(�v����Gs��Sz�X����c��ħ�ġ�@f��55�V�Nq��#=�����"^ ���+k�ԉ�o��	��Tۂ�=B�`��O���
l+յ=L�����5p䡁�u�x�g�~��%p�'��Fv�P}e�p]B�� �A���6~��t�d�G��W���7R���1�&�Мlck��ݨ�	��'�b_u���`*���U�>t���̜W���Ɖaƶ�Q:�$r%2��-������H�`U�	l�4�Q]���D��t..�<:���&l�6�-�fqr�F�Μ�Vu��ڗO
zd�+�ٷ��5��2w�0z״�s�
��e1�]7��X��K��㋯���_������έ�����땑��nXǆ���!Y�8�ő =��|ݵS�uej�.|u�6�<~��>�wѱ���	�w���;�G�cb��j*�hE��4�̟��������/8�n=GWm���cTY{Si���^C9��k�`��V���(��f`��\�t���~���+֑�̻W�y�l��SW���^+j׋.��i�RF]J9C��J�F2�L�o�͉M;Y�o$���;ę���)���[Ϲv�KW-c����֕ư`�8z�lNY|2Jj�7tC���$(��[ry�1���l�Č��o8uU�1l2��d��	L��9l���٩7C��%���nm����Y:l"E�w��4eb��tJ.gTuwvL]��~uCƱh�X��t�cF%��M�^چv�%��:��K�S�C��/}��0��Pڗ�P��J����rU0Z�K��0���E��:
ܓ�Uҕg�_1{�R2�é�����)Θ;���u������"nŔq:��[f[�q�j5��E8]ı�&��nρ�.�o������m��f슯�hj/�&t�g*oǗr�7�����m���2��Us�3�-v�l�w9��~�u~��^Qp
�PB!��/b˴�����ݯ���h��+)+5n5q�:��^+��U���V����l������nh��D,et���W����4�V�޺K��[�^�z�Ft7��;�'tS�����E�g��8gNesq.��}�t��cU0�����/ǨP�"O�._�y�)ڍv�~�Atr	�$m��&�C p�z\+�:��)��N�{�y�N��D�~̢����s&|ɚ�/�7�*��0��<�8��6��Q�����SJ�?���o�V�U�����׿�� x��v�V��F�{��I�w�c�����]k��~;_�9E�U�X���.��)TO�����뽋m�>b���l=���_���*Q�m�Kn�� �8��G��8�n�	4i�D{"#��4��ꄼ36��Q -n�D��W�0y�$���$�&C"Y���-��!�I��M���4!l�����%��K�IX�^�j�U��mu_�P�Hq��'��~��r&��]��h+<K=�
4f�h�U	d����FcS�ER/,;c�
�����0��qpN��G�b�J��T��iďG/qFYK�+Z�q����FS��Ry%#)u��k1,ٌq�,���Z�猱8���9�N����ԫ	zN�d� 2��鴪����w��%S�����'6�e�W ���Z7����'�����Z:c��R(���Ɨ{�^o ﲾ20�g�t�iΔ��h�U�S�_�{3�d}H2��N�d�Y��K㈹�
yʼ�{��ث��N�v�Ȇ��w��ĀG2=���g��,Q`�O���R���m��uu�*R��H���33�s8S�F,VV��\Y��:��E����R�{������s��\?)<]�>Nv�r��ߤz����vqRL�Ee]����79�6x�O�� �?�+R�k�ع9��Y��/R����	��.rU���*� E�^R�W©��W���T�*m�����0`7PS��A몃,�Z�)ڎމ�t	w��Ê{Jl,�mn�5���.�Ѷ�ƚ��B���P��pI_��
�}M�y/:�O�x�җ��N�Ҷ�S#g>�O��_4����26%��eN�<e��|��2#KJ��Q�V�bPF�/�cJ��s�LgXadJ+K[j-��u����]J��I�;����ґv��<����P�{P��I�䏦�-���7������t�O�����ѭYFw"3T���F0i�HY�$�e̲5��l�\f��D�Ҷ��5��/�ݫ�}�������l����;�q���l;�q��Ճ7xp�_]��n�Ϳ�@��g>��>��cĠ�*p,=���ǰb�B	�0���F��6��[�r���C|�� �����Sxx�6_}�='_b`�����/@3�9ç3o�L6/^��Y��2l4[����ʍ��&��zη����'��o|-a�1c)C[wg��)���>j*�&�gƈ),���5sV0��No9��w���;잱�%3���{_��ɇlX��c;N�|�6�Yš��پa��l����޽ON����K<�y�'������֏|��"G�g���%�����Ü�v�m7�w�^V._��5[X�t��-dբ5�<p����w�dݜ�l��������U�w�['�s��5�;/:���9 q�i�
��ϴ�s8��$�-�o>cՊmL:M�Ge�-�Vpf�&�H����s�7��ZVL�ˢ��9~:+�,�ⱋܿ�D�a;�&Lg�9�^�����|�|�._ɖE��<=�g�b���,������ܯ����|��OL�7��h��9q,(�wó�f�ˣ�R>[����_,��'3��b�Jޚ���W���7}+�^��Ƀqk�?~�F��ѫ�n�ޑ}7�����U�?q3��_͇�����<��G#�b�r9�����DSx9t6�M�����9�U���L��|��a3��[���Ɣ��I�@�[����`�K�#�T��{�:UZ^]D���鉖�@��Ǣ;Ì��C(�����M]�n�F���_jS/���Mj�0��M��<g�)1냩'��Z��V����皋�W��M0i�U� fc[��&��-؋V��fR�{T�i���=�?z����*��B�����'1�8�^�%4�70���v������^���]Փ�j�S.�����!\Jh�kO�xƲ�#�c���Hy�t#ohb�Xm����w�S�k�������KV�������V����s4�D��y /bJxk�Z��9Ȳʙl|�ek�0y�6y���/���J�]|=�$"���a�~T�ﴀ�����
ܤ�@G MKh[��M\%@���mhenF?oFy;1��%��⭘��Te(���͕k��.�
Ib�n�{I�*��\�� �"�X�8��Nl =UI���hMG�c�N�w�G۪m�Y��a^�F�<�2)8����G����a�g��P@�6�����$��)}nys��^�~��p��XT6M��g�@S�	�����
�:�q˓�WE���J[F�09��Q3�b?˘����-S������X���;�'�i�rM���w�>�L���/>��+N�]�7ov;����t���Ļ�����t�0ң@�w��q����o�S����O��9�!φ�rL��v�v�\��4h���^&�R����r�$�͖L'3r�)�ԣ�\�,@e:%_Oe��F�ӈ�ޮ��.���9[
���#@���&��*��"e��U��z������+����"��(���7�C���S���U}�����T�����j�������$����L���,�'������C������]����@�����O�@���hk��#TO��W�*յ�TAʜ���J��i�L�8څ:Q�f%�Ö+&Y�rN�膅3���jW9�n��2Jc���+�@����|����|h��=��t��-"������3Sa�_�z�p����*݄ؗRX��n���R���s8��}�L)dMx<{��8Z\���"6E'�9*�=	��.f�o K�������cgB;Rsٖ_���j֧���ܕ���������+fs~�7/R��+������Ïy��޽�����g|��}�����7y[�}��#>��	�}t�������xy�9���{gnsi��@��u�#�pu�1.m��M�;.sc�i�]q�����a��_s�O��;W^�΃��ѧ|s�=>���/��7?���_���3�{�Ƿ^���w`�58�H�Ht�<���n}���Y~z�}^]z[ �)�$̟�{���ˏo�W�����vg��	���}��=~:y�O.?���᫇���ŧ������|p�-޹�/����d���u'���}^����}9-�vq�,�����<:p�3;���	�X��K��sy�AN��¥kx<s5�����ö+���"m�$�^�����}���o���M�8ýs7x���_|"�x�g��7_����\=p�G�����nH:]�y�G$]�_��G�U�����|*��`�V�� ��qv�)��;(Pz���.qt�.�8��}���y?�����|�J5�����Y+�;}!�W��@��gv����ؼ�#[�K����=�]����g�r�.���[U]���+w�s��ɽ.���A��ڌr�8�Yx��%�w#3y�����[\^��ӣ�qv�t.���1��{�:����8�s�Ύ��ȉ~��{�z�x�1j��]���HU;��gkmo��髮��<�������N�]ۓ�ͻ2��%�z������͢�r�M]&�0�:��W0�j �IR^�*á��k��[��x��e۫C�)^>�΢�*�iy�Dǻ�@�P��&�� C)u�_7�JY#���T���M�(� ����b:k�%a�:A��.ew�44Ʊh�G��H�����Q����h�%-��wC?~:&���8�q�Q�4���.8�~ɑ7��-��)8�n�	�ʤLoz�*�<a#�O�h{���O�x�S6�����o�z�n������Hn*���I�P6��sb� �R����������]�z��a�~�A>b��R׆�!l2vf��{m�x��+�H޶�y\)�'���£,��Ŧ!���&c�_g��9�6*������	ܽ�<�,�d����h%�� m�$�n�I����fnk��e
	��Ű�&{�.]�}�e�O�<{�*�	X�Lšd.���m�ݜe��+"�ꓶ��Y���5@����z:	R��J?��;�Y�4x�J0V=yyuX�O�2w<i�q��{jܒ�2����C0P2qo4A��z�;D2�d�yhJ���r+z��c�f��wcX���X4�#s��aD"���Yxo���?��~�d��҃��>��wB�7�&mGr��3^��=�>��[����� 6�;���K������z�	�=ttq7�U�x�i��]��򌸤o�V��7�;af�_!o�@�^�2e����	:�j�L7-"�,Is�S�uͰ5 �B�\S]�L�T�k��)=M�kX�N ���O�W�}������V�%��zy
���נ�z�T/������*���P
T��x�j�F�j��)����u�?��psx�<���������a��ٍ�T����F>��l	����C����fjO[#��Y2 ���V��)K#m=�W�2_����� +j#�i����lA��>�L�8���3nj,�,x�&������C>	��{+O�����9Ep=,�j9����|���z�zK^�����-�:���+�=��Ĩ�%��_���>���Jx����e�PU��|���)y|�Y�/9M�&!U�K�'�̟"S!��_Қ�s�rM����CLl���I��o��P�ws��}��r��&�*�Vݛ�R`�oQ���CX�s4[�f�Q3�b^��Lo;�i����~8+ۏe^��jG��j:D�& ��������k8���j䶁1t�e�_6ۣ*x����������ד+i�(���0��(������^(��;1��+Ë�1��0��e@Bkv���U�iP����˦��s�Z^������l6�񥽘ؤc��2��'�;�`Q�x˻l�4��B���u:�6�Ǖ�,oZ���SY�s*��۲��Y�΂�qLk9���G�^�ao�0�gB�X�3���03�)�C�08��Q��LNh���L̪ah\1�#��PȰ���0�;��7�fw��N��م難�^��Yݙ�י�9��؆����^͔�:��bbZ[����$�`|J��>(����/etj5c��0!��(>�ڞ�{@���ڴ/K;1�?�Q��M��w\9}J��E����5gBn[�d��c
XQ�y��WZd����z�F3�'��Qٌ�e@\�"2�����<F�4aDb!�����B�n
M��g\�<��L`��A�$�9G��1�
�<�h�N���:�at6�R��Y/��>�])�ٔڜm�mY�єy5��iƪ�R6�5e��V���1��%����bIz*K�2������xf�f173�����L�d~vs���S���4&�%0.%���N�aZN�33���	��+�F�4��󓗪���S"�2��HJS:`�R��[;���|��S�#�ޝ^��
x��r^��zރ���V�T)��ohǟ* �*e��ف^�Nt��!҅%�bR�ۼ��ס�)e�E���h4.h��4n����1	��3��r^�5�9�_W��$�s3�`[��ֻ�+�g�r\�&�0:�GD��+j�h�Wz����W\D���Q�5��?Ų�C
'�d���X{���>gي{����ø�T�1�`N���=�cC�W+��˨�����O?���ȓ���W�)�����w�8�-Z��?��fnl�]�������>����x�P��)���������Vf���x��Й�zy���UrG�����1�3���~�C�<�V�>4���$�Rd��Cc�ڐ�8_ �|?֕�p�ȹ��$��K��<CId�"�t�"�T>���X�(U�S�a����]�����6�R/V2E�F4�zqkЉ_+��A�̡�*�yV_���ÓW��y4���
h�I��&�M��3'��:��>����)�W�K�Y������uB;�=z�=�O�$y� �4�(���}4e�e}�h9%k��؈u�j�R�(��0�/�ݰJ�C�<�F��= ������낁XL�m'2s�e�zȣ�_��+M�n)�j�.���]g�|�b��Qں5@�>�z��h��*�[�>y�0*��h�5��e�Bީא��W� %@ڿ��?@�~�;u�XmjIo����l]�6$9ۑbgF��!Y�d�h��B�z:8	�)^'Փ��������j)��@`�'a�|����*�5z��@�_�x��*��F)`����( ���M����T���}��5� ����:��=�6J� �{�5��E��JX<���R��㎗�O�BWl��L������� �2��kHV�r�e�M_C��e�V4���H�3�ј3m��s�х˦�ܐt�#z�Z�{�5�әit�6v#���g+/��拐Nz��Sc���kiE�Jm��;_�g�;�y�?ߙ�_���z�q�#=W����K�@�r�'9��O��$�7�>��#��������������Ǐ���g��+�,ݨѷ��̖Z'9���̇J'J�](�w��ԃ<c���)6s���%�r��YU��E&.�{P��Bs#/J��RWʍ<�4�����Rǁrm+�Z�%�^�kH��5bH�5��L���	w�}�h'�gّ!��б�B���5��lm�E��t��;�RXu�`�[?&��g�<��(N��;CXTJ�fy:� �L|�Z
��5t��c0�$�&ۅ�� ���۔��K���-�v���:'��=��N�4����&�2I�
y�*y��Rv�#p�{VK~Kn�����k�(�0�X���#�����Na�_2C|��0�h��'��5�ђw��G�Ct�b��[j;�z�1�(���T��P��Cg�@ZIu��3��З��^���ƕ��������2�z������}$��B�a�y�t�,��%P�qR%K�(�b�F)�Zڅ��5���j;��Nr�K��}�Z��N�ELK�.�R~��U`�LgKzzEP�L7;�Xy�[
�^�A^tC��uò��'=m��n�M��'������|�`�CksI7��պ���7�������󪸎�b \̭�˙k��E^���������p����_GN����q�(�_÷v�멃p�������U<ݸ��v�䭭[y�i#��/�Ԍ�<ٺ����pw�R.-�����U]_=��K�3����O�����Jn�Z��S$��0T�zf��v�©9�����������p���
xO�z���O o�@�(�������h+ ����� e�zt�wc�uH�wS�ļj7�R�Z��A�s��,�g���=f�;�6���:G�(�%��JX,b�7�D�8-=���5Dc,כ�Jy^�u��oĠl'Z��W�pu����D��� �y��.�[qU �:���{�u�GOx��'?d���r���q��j��������s�`�O,���O�ZS��OYSzW(��7�S������~WG�Sjx�{zj�k��݃�b�$0��^�x/�R�6�'�~܎���U\Zt�UY�o���b���:~�I���&��{�2��4�//./�#D�yRC /s��1�9�N�DL��^�$F�v�
v���<��;q.��Q�$�C��B�Z
Q{4P��WI�ZG��D��#���V#�;a3E��5�ԥX��E7k�d�T�{�C�N�Ri ��	��u��u�׍n�,�|����e��? Oc���a^��
�y���|fy���`�<ۈn���i��B���:b"VDPUz!�1��N�0tR����M�@^�Y�d�h���0� o�)c�z����|�0��g�h���W2���17�^P55��2� K7���ɧ����b6�[pH
���g�t�fb����������ڶZr��O`�R�����: r��)����q�I9�l��딹kׄ$q��t���?�;��f�����;�'��7d��_)�(1�#�Ԅ8G�M*tI3�"�R�s}⌴����� K9_���z��(��0�%8���`?bb		T!O��[���#�y��~�+�)Ra����������}��
P5���񑥧l{�M>>�u��0(��7)�z(��+`*R&LW��)�)j��"_��F��y��W�Uyo;k��L134P=y�x�/��_�<e e�m�2S��(�BC��1���y��jF���@#}v�9q��]�2L��w��y�j˱Ff��r���l��Kak�V�F���oJ���}���<,�O��xWہ�����8���F
�͂��"�_M���&�CA
LE�5�;���/���ȯ�|��η��,����r�On!��s�槀h�I-�\T6�\���M��?���lheiMkGg��ZP*amc�Hss�M�i�o@[sڛY��Ȕj1��K~nah,2���1U:����:F43�}Ɩ��	 �x�Q�kB���@�>�F&y�����C8�
X�+8���ɴ56 �ڀ\+�%Ζ8��vn0���|N���'ǔ�h7�2`��+�G$@H
�'�iR	?����tJ���)�0W�{43�����ڮ���?s�>��� ���bn�o���U���x
�E2:8��R��x�*���܍��N�.��X�����"S ��?����cZV24ؓ~1��K��Wl}""�Ɛ�`F��00*���1��	doX?�V�kt�(���p1,]���5-�hg�@'O::9�U~#l�b�L7yE�z?/?����[Wn�W8}=����T�@�$@Z��d���qz�B�J����Q�FO�O��$���E=����z�Hh*y2���bXv�_����+@�L� zK�{��T������0��x�,���;�����w��V��t�𡛏?��;���A���X����u�颶�.j�g��I�����,"���~���>������o���'/�����\�~��O���r����f���:t��op��c.�|��{9v��n^����ܾ{�;�o��ʾ�G�1c�x�vΖ���+�Ό���;�.�)LN���n�h�U��k+��:���U��������k�;U=j�|��z���x��O�����[�����?u�Y�Qz�j2��Sr�0)^���<G7Nx�#ko�%O���Ь��5�iZӓ6��Qֲ;��-�.�70�,��"ѶS�c�F_`�(\�)�i�q�ތe�蕝FStB�RTx
��Kx��*��JS)l�������E^�|�u�n{ȼ9W��nϓzq5��c�*�)Y
���ǒ���`רF���!O�*���O�<�����������.c�{0����b�/?��1*�=�O���k��� ��&�����Ŵ���p�.S�<&h�4-�=�{�V�%t�Ϡ�sV=����e)c���{�*Y��]ؕ��4a�Uz^w��0f�[��&�FNj5M��QӬ'��"6�3�@bR+5i	�����.�q�b���Y����jM�(yZI|�z)z	
�Wו8�s1���� t��'�櫐g��#�)��������8{4�Y�1���Z%�Z��k5��0�`��E��
��:�"{�3��ْA�
�C��z�k���j49����1[2�d��&`�4Ө��\�a���!��HJ��DV�U;~�L�ǂ��]}�mϱx�Ƥ%�C���O���6���L��O��l� y��yǥ Q��k7@�Y��AVI��A����@�&CC:˶2�U�@G��>�&D�ۓhkI��ɦ�dX誐o�E������:�jx��)s�ZY���bGP�7!��G����k��w�U�����O��+��O�'乹	x�������R�M�3��g�T�y��ӠF����s�s��+�)��U�+�@���T��D�B��C�<e�vE�����m�<?����j��`;b�525⠋�@�m�x�h�T�l�@��T�%����J')�Cd��C6V�H.e�@�	)�>���}#'�Ѷ�+k~�N���<~�B�/�Cr�A@�Ǡl�/�QB�f�Kd��d�Kt:?��2!��s�6!�D�$��S\�'��Gb>�G��?J����[�ɨL�;J�i�H��7=�}�uv���k'7w�е13����$_v27���.mt�� F����k�uh-�HK}mZ��e[QS��j��-��h�g��Z4737$K�Qf��-F��aY
`�Y����V�#�TC���:��I�~�/���x~
M��&��b�� �/�ϓtn'���3F�����Ф9��Ȃ�(������21��ʖ��vt���LSW���@̄�R���C[�gF';8x0�ه~�nt7�����\'�kNc:�7�������q�j?����-9U���PO�zK���#$�A{�����>,����u�d�@�o9�[������g�|S�ۚ���F ܊��t�������m�hcI';k�z�3�׋�n����ް� F
p���_8��y�r=I��/�q{E��.c��=
�D�=0��~�r]8#�"e=�^�Q���;�=��NRx$�����Q q��=B��@^�������K/1*����;P��
�����Ƀv�>w���x(Ko�*�$_V�ﻳ�'�#�$��:��#���H�����y��G���G^|�'��a��㌘����WP?q>���I�~4�;�����܃��è�7���i�UU�^��:�Ү�(��N�a�:c.�g�g삥�۴��GO���eƍ�̼��X\Ϭ�rnN��N)�1���aN��v�ة�.�xJY�&e��,�2��T�l <)���!o���y+1�ځ^�Nu���([�"M֋�c��8f���RVG�ɷ30����6�9s��z�v-�̜�[X��(�w�gɚM̜���O�]ҋ;b㛎�D�N�P]cY��1�W;^��+���A��x��AG OS� y��h��Z��{���Kv�����l��l������j��� �>��:F��3��C������o��ǿ�y�`ȿ��/�dE������NQ�m�c�@$������^r�%��Y�k=K�^g��;l?���������Cy��hJ����K�E'�ڙ���;,�Q�J��)؋Q�>,�
�N���2��������D��;t����<x*&,`����ڸ�^�&��_Im����w��r��Y�l8J���l>���7ٍn��0)]��^���Wq�ʺn�f�#�yJ�<�v�XI��*�+�+DG��@�n���8�.��r�X#0�(V�d*�h��E/�#&���K"���VrM��:���L�=��k��yM��G��h�<�~���I�H�W�]�5q�Њ�z��b�K2X-:�m�O�OH��d[����������,�p��kN�P>��S�hl�G�t�΢���	���ii���4@��S&�?��i���T)���S %+���@������3Rح70��l'�j�4�#NO_�n�@��=IR�&��b�C�E�Eȹ�zZ���T/��j[2cS,͔^���U�
�)ՖJ{�FO�?�Q��
m�
o�����y�R�5z��o�k��5�ٿ壪��}Uyx��j�nT����������k����W���ꊫ�����Ӷ)ղ�8���f�W�����z�d9&q�`�xP�j�[�4~y7�]�!�vK��ɻ��-���@�Jl_'n�Vp*:����N/J׌X#S2��=E��~��';/>c�s}g��N��_ǂ��'�+ ���!l�e�k0;|"���(�����;�M8[������H��$�3$]�If�o�c8ǅ��GCh���C
 �WrG�r�aC�mg7ںx�����Rx�q�@Mɗ
H�YY�Rאm}ڋQ�������k%�K3��j==Z����;��R-�^�oA������В��洰�$O~-$~�iكs����'��.��I\��PjeLk9o�\��X�X�yp�kR�`�-��� c'Z�[S�ѣ����!�?���@<�ݛ�R�݌ӵ�����ԌfF&�7�������	S��Kd�@�(��>	t��y������r���q;��w������:hY��3����w��=�b��=�P ����vb�����8F�%3 D�)0�.>���
b� ��P�x����!�5g�%�,ikaN��mLm�%y����,�����:��ŋAn�����'��.�E�}��
�]�c!Y�V��Sry/����?�7x���"�Ő���I~H�g�<�m}X������$F
ޱ|��J'z�۪��������@��~�ܾrE
0��l��)���\%v������*������J�"'']NI��c�Rt!�������X ��O��_�r��E���E��#��FJA[2�IL�&R������$5��p13K�.�$�����\�Ǧ�)���@dB���$�\LaY[z�����8|k��f_��̍��̄e��=���iL.�ɔ�Ȋk��m3�=�L�Ӹt@�KYOw��z��o�!�G�U�=�(��'J;G%�${��{�-v5��O�r]��k~ �R���=t𬼈�ʣ��h&����ݕ�װt�r��-Y����ټo/;���ą�\�s���.�z�.�w�OD	�蚅ca��^�pJ�:֟U�Rl[C�X�F��S*�iU\���U]C���mo�1����cɞ���r����pJx�Nj='�K�&F�i�vy�pd�@��&�_��;���+������G^�=��:7T��x��1�w�Bxb�c�L��Ľ��Y�c=K��`ށ����;��)�<�)�+����ZyhN��;��~�y��˾�=���îh��|3�� �;4��x�кm�O�Ǵ�+'�7t�8ƌ�ƴK��h=�'Ρe�~����5{��v�:�o�����0v>N��1��m�*���2v�&K S��J'��Ͳo;:���
����X
�}Ѳ���,�
|����kT���S O���n)VͧbQ:Mt'�9���]�L�N�d� �P�:��Kݯ ��x���4[�^��N~���{h��Do�5t����S:�(=�?�h	Wx_�&a�0=���Y91�v�%��&|��c���it�}J@�;�ț̘�D6��ޗ͝��`�z���א���Ҵ�l�B�q����@�:��x*䙨:�������;V?�Y�)0�T�)m��J�x�Ȝ�Ff��v���`�$��
\�li����T��
�)��fa�7�K�0&D_�������ks��	��>::R��Uڣ)R�Y�������o��@�Z5����]�����񬽆8��
}���kT#�y����+�)�� O��>%L�b�[I�(ӱ)�g�#qg ���D ���!O�Ǜ�ii@��Q�j:2�g���͜�&�M�KK?nx�1J��%��R*�g�_�@��Z}�cD���Z���W�[���~�r�3�,=ժ�Oӛ��5��RP�50���F���s�����lbI�䳎���X��ʆ�6�Ԛ[�BW JǚJ��"yV��B�A�f�{G����O�i���m�# �O_�E`���-�J5�,��{��۟.���68�k��mgaC�n+���T �B�C����Pc`$@gD[3{�͟w͍�)ӱ���[S�ZX���B¶�)�Rh�rD��9��#N��G���9%z�#i�����~I�O�x~r�K.���
6	��Ҙ�A߁�fΔi��!�^���k��kߥ��"�53�Ы30��H
��J��
�v2t`�ƆO�ZBn?��@s[C+j�]�l�N+':�;PkdE��I3�=7�tP�U�j���7T[+m�I���*���r��o�mq��S"3��OG�`����Gཱི���1�7�b��+�*����@~7~��ɑ�t�
�(i���F�݆�F&ۘ���Z �?�!G]�*MO��{���Y��7�(�B����4W?n���{j~N��R>�-g��}o{��a�z�|���*��#4B���#�^ώU�>�S R#��/�E�s����������X��`���s�W�l�l����K7� 	Oݜ���Nr}7�`:��j/aj��M��UfV�w��R�%5��~�yԺ?[�u��8~�"�;��,�5y���&,,W����ĕ��Є<�s�ɥd'�%�ZHvr.٩yd�>�޸�$U�!����&�Thp"^�l� Ua����PU܆�]�p��Փwa���L�cK�1��XR"[58M<�JY+��\��G7�t����t��j��i|��"���=L o�~��<#e���������]UG�l=�H��0Mx��l�N�Đ��:y!�Lcܨ	̘:���V�r�F�o����ٴg������#�}x�[����I��EDF[m�04�� ]M�B����� :%���*�y$��S.��TT,Ts�vW�+���.�w�c���̘u�#ӹ�ܕө�l#��s�=�8>t�@^C�����Z]�H�<����^VV����U o��;�m�x���A<��Il	�^�͹{XZ0�5]��l�]�~�֓O���9a���J�N����h��+0w	M���Ƭ��B�ͯ���*�K�Xf�����Ӹ�ːә1s	#O�O� ���N9s�T�]ÒU��:`em�1f�,6����uX�n#��s�A$fW�c6���
i��ۊn��]�Z�����؎Q�J]g��8�hYw@ǲ��h�6Gc �g\���E.��#��릳�^b���@/�f��L�I|������z������~�0|���Л�Z��B3�1��c�O⫩y7�S&G�s�jb��0���U,@��[�ݹC��b1����G�����[�`�����n��i��7�&�����&�SGO�0�Q~�,7�p�̷�ݝ�)g�`:$�2WmC������	���{y}gp��,�x��G
�rl�h��2��4��ʶRu�c,  ��oD��ў��{��bM��H��i�qf�x+�X�bj���6�zy�:8[Y�j낿W �!�*X)ß���^�.��X�!O�,O��=m8R�J�vp��n8�)=U�I)��]�x	�g) �x���~���
ܩ� ��k˿��S�n�5B�x{s��ָO�V���wj��,�S�������O�����+��Ԟ�"�}�r�J��xi�G��.)����Z�la�hSs�	�]6����S�5�!�@�p�i͔�
�)�$�04�k��b��e`߹G𵃧�C��l�3:�G�E�r���%%VvT;����_��R�WJ�����k�8��ތ�b4�s��@^S{�%��]��(���	ImRI��"�Ƥ��?��I9��o�2���I-oWv�]8�ׄ���/���;�z��I��Շ^n^��u������*cSZ	T��5���nO~W���Uu�����=�$
�pl-�2����V����Ěf��i/���ٙ�}��j�fط�_�n���k�_ە��
��驰:�߇������%|�l9߯��׫7�񊵼���y�Y�(:]c��ؓ/i�74�KÇ�ٚu|�z#W'LepJ
m%�)��*��R�8��������`�Z�^�������S����O;�Vb������{�%�P)���H��L�|�Q��u42�N�a�7���Ӫm�q�,�?Äڶ��/`BuK�����/���v��TW���My�q3/����b	��}��8���I��o���M��[��v���_F&�Z��[F6Ë*�S���ftr��
S۾���d`�@�P��v���դJ~M�˄�j�ȭ��^ ��W8|��˘�$��J��FK�\jL��e|j�!���O�MX��Cos���;0R�3�>.A*p����$ AwY���<#��1�>�!�񈠝[ �r��!t���F��V�~�{y�T�D��qr	����s�d����@uwNJ:8��J7sg�<��q���?��yn�����|�=������FQ����l{X�wU����)�X����a+����1��"+�������������o:���\���5�&S� �o1�������:7��s��GW�d��������4������O�"`*ZA�1HZ�~�.�s����4�:,��)l���$}�0E1�Dc��\?��v��a��U̞������h�*�\Ú�9v��n?���k?u�3�Or���=�ϱ��h�s��|3u�z�&S�lM�9�%�gLǢ����ESv��s*�
��C+�$����U�ǩ�)*&�`��{,�}Y��ISr�|2��;p( ��O�;��3^�6��JX��7��H�S��? O��B=���O��_�ё]o����{��@�y O��y{�2�����܉��e[�3��c��~�������:��;hʟ���n���
Z�B���+�-<* ( ���s��o+�����D�'�魨�=��c�0P�|�8F�Š��L�?���f�y�n�-�L׾c�<w9�v�f��l����;��`)��z�WT��M��`�����q��w�,�$l��&�c�i;0��wS o8��=��бh��itLZH�)F�(�u��4B�ε�0ʛ$0V�A|L�`�S���E�F7R�.�:a��
�q�PL�'`�lZ#�c��;��f�Kt�H����N7����b��F>^�=
��hGB;n(��S�n2���\K0J�I\�U/D?�/�-0`�Yf�:ĦMX5g3K��`d�.[6v���q���u�H��f��/7,|�L�9�o"���o�Ӗu�#����yg��b�W:�L�T��)�kd�'�i�j�[;�,I���G���uq5�"7ʏ���ۚ+ �b�G��vAzZ��>O}�:􊳡�ֶxغ�'�qDX�����q��
yJoY��S���_!OYW�i���)P���"�\�_{�z�6m���S��"`���U�����?�o5�W���&a������,���k ¿C���6Vj/d�z[���R�Q�v^�h�Ke&�אf�K��6��:�G=�ʁ)&V���㊾7�����
���B%��	�����'�Q�r�K� ��)��=�����\��%2��q�̑������y��7�NaѴ����7%���9��+\<h��E��9r�$s2llI��!�ĔTG'���ܾ��>�sOqt�-�̭�;yg��Z�����������:�G=s0.��fVT��A�/��Li#���ꪴ�2�Q���R��m�eH����Y��:;� 	�R[ed�z�Z���ĞF��0���:U:o����btA>��w����c-�?~����JUpsC6��!�OŪ��W����u~�XZA�~��ÃF��*�]v�tg@Q����ӷ�Σ;|��>_=³s'�ҶM-,�*�j}��Y٣o;�O��[��w�<_<|Ωu���\¬�O�ƀΞ~�Y<����sb�6/���u˹� �[��Hi��o@����ߒ��H��W_p��&ƚ��yz�k��Qe��0�H�m���ʺ���{�>;�ob���l�?��:1*-�J�����cƔ5����xyU
�n]�oڜ]�����(��N.�xQ

�������Q̯	J�p�5U!o�O�Z�:"$�����v���J_����a��u����=C�6"�_�C��/���KY� �F�w]�Q�^�������G�h�U`�A���ջ�9!����Q���K�>|#i��'�T!����4�;&��Cns��]�0�j9�}]8�`	��d��ӷ}͋�hQ\H��M���\��iS^)���4'���l
RTUf��,����ʲs�JH$9*���`RbBI����p�\\�� .$+[�="Vӟ��Xތk�ְv�$j���*���f�I���@^'t]_C�{wt<{��g��}ϑ��Թ������3�����M� hFC����O�Ձ�u��;�v����,ph���WUm�1��4�v�ǈ��1k��,`�����w�����l��K?������gܼ��+w�q��c]:�ʽ���1ǈ�b˰�.�ʪS�&h�JJ�bR"L��ZM�	НD7�0�9��=�&W���F�/���U��x�CV�ň-��6�0��&�0�=�������a��{D��z|���<ū�H:9�ߕs�TAO��?~��������'n��o�� E�l�B.L��҂)�ﱇ��2��S��}��;�ã�U��۪'O��Ky��h�^E��Z��.8%�rM�I���B�S
�H4Z�t��C2���̚�VdC���͐>��ޮ+��`��l�r�1���DN_�ŵ[�ٶm��56Ҧ{?�K�)��wh�P4U8TmǴ�y��{�Mۋ&]2K�N����%P�<m���X�@�J2�y�O�Ze�����S�M� �+���>MLO,2	��%�Y O�>�E�}z�[W�M�ptk6��Fg��h��f�}4��°��ae���h��C;|Q���vT?tSG`�7��Ab�T��ĭ`�ͦaݝ�V��7�8Ӗ�f��}�]��U��36�_!OB�IO���7X�p��W��=�m(K#����)���A����n�|/�o��������-G��J���b��3����+�����liJ��!��ll��@A��=�b�� �F�4���jb��(P⯫��� ��	>v��ۻ�#娨���U ��W<lJ�lCU�F
�)�+m�\���e�r^�
D)S�5��Mկ����
�)��w�z�>��_���XC5n#�)P�o��;�5���|��0�]��6*�n:F�|�#q�Lcf"�7�'Km;œg)�J��"�4��k�����ځyb������o�7Ȼ�'����S&������ `��k�^�h��_����8���� 8��Tےo�B�W ����)�%M�xP��F�j)�6�y���!��.�?�.���K�	�z��jhEZL
�{�g���t�6���zӺYW��ǝsw�����������'���u����,�ʮ|XT��@�K�Pz��������=T{ߚ�SadL���
T-%ߗ��+ �x,+�Zۻ��N�T
�R+ju�6c.�(P��^��(�&��)"�-�ܱ-�&�f�y?z�/^�����I���Ȭ�b�Ia�w�
u����X�b˗����(C%�]������e�[��d�V7�ke%cf��Ӣy�9�o73�{�0��'������ar�:�H��5�I�'ѧS�M�ÆYK蔞����ʙ&}�#��)cٰpkW�Q7w��6g��,�Շ&6�;(l*q�xf'Vײq���ň�ChY^C��*���3������#�[{�P:�����0VI8��M��tʭ�eZ	�R���Mw�h����;��������.]Ȩ�i�_@mAS���O_1&�HY����'���ߏ�n^̱��Nx6���Axd�񪠒��Ju��~��O u�>�U{�*��띂h)��F�{��Fd�K���SR%k��kfC{k{Z)=~<���I{w���1H�}X@�
�
�ֹ��m�N]\���H'oZ�q�\����]�Z��5 �*y�6�m=�����I)��#yZ;��e��}'����|��K>xr�sGwp��!n�?ʕSxt���������9��]<����r� �O��q��>�����]رy5{�������޺��G�i�N�ɠ}pp�a@��m2�U�\��������'�1�]T֋�rt*�̪�S� y�^���튖s=:�Rƹ�G׽'F^�1����0�GK=M�׹(�'��Wǥ����9�y�e�6��l�@bf;��� �c�ձVmd���L�8���vq��]Ν<+�?����}�Ϟ���ӷ���7�����i?rF̧݀	�7�5GO�p�I������ ��ƶ����ǰ�����#Щ]p���Uq��Wp�;E��,�q����3|�M�L>ș��;��v'_����)���?|��Bt*�)���
y�ʮ_���;�7������7sS��=�C���&~</�鄅\���Mf���V�x̂��Uț��C���AS�M��4e7�h/�04�ѕu����7=�A�246�wn��clFAeG&�\is?n*sg�g���6��#ƨ	�e�Vv�9��q3X�t��z�'O��k����3H(� ��%=���}�A���KB�h���|/&�1��F� ��y�{�v��h��\����/��K�x�%�(�l�q�$��h�
ю�u��.ɀ��0M�#�#Z�0��Alo�t�z�>��ay}�čǦ�!�&?�l�/x��1�v�ag��tŖ�DM@7Z�6J�����U�~u`�9�&�1����X�ytB+�bWG|���9���;Y�e��dfe�KA�y��n ��a�����Y_W����;�b��(c�pJ˰�4&z]e�P]�'���aS[��p^ �d}��B���@�Q{���S�w�}J��T';
\���Q'����Q�I���tɌ�]�yv�-��g�M�@h�����,aU�x�qw�� ::�P�+ dg���x��H� /o�3���=�?�����k؇O�����] @ �`!	�ݥ����Ipwwww
��-Ji�o�Is?��>�����3g�dΞ�{����{���⪉���&j��U��+��j[&e�?gg�I�Я+X�����rQ�U.�˨�S��QE�����̫��9z�ܪ
�T��7��7���T���ͣ�r�)�SC�j��r�S)TT䭽Ws�"-	��R�V{�ڻ��ܚ�z+.��rA��=Qp/��9��@��R��Ŋ��<x�Ff�%K�����^| ����m �U�&�8��֝z.��󍤩�aS_�:z���W�\�����0�KW�"�Hq�&�ڙTQ���a6x���&m��V�T���G/]������L�_@��5�����~�J�L���E�x�6��z�����Rc�kǡ�l:�=77��o��Q���i]�����ռ3x��.�30�<b�ݽ(01����S�Ԛ\C+�:���S�א"sG�;z021�^��TЛQ����^=�% 6y�Z�kK�Z��$�a�#"�ōZ0�C7�D�f����3ܻ���c�Фq+N8��ISi��*�ʴ���+`bfI�ܺ�[���vұ]{
��iW�}�2��訆S3��D�X&ϖ;9b<��Q),�viU��K3y�U�g��8֬B��y�ڻ�ƭ�Q�V��%SA#;Z{�=�"*T%U�w�C���d+�ס;q���Z��Ui�@;�D�
���c\�!^}�S�Ѣj!�:+j��2�b]�V����Z���Gc)_avU�����M[�;n:Y��Tw�[T�#i��K_:��ӗ�N�\L@�T�s��\����1��O����eA��|��q�CK�\�3c[ZH=��r��\pI�����Z�
�PzX�A^9O����#-<=h��F{Oo-ʶw@�C�LKw9WozH���S@O`���VvZ����j�B����{����MR-ΧT�1�9Q�-��w�;wE/��������k��>���tn7����#<��ׯni�'w�����|��������cr�q�9ǃ�g�s�$�����gy��lO��t�N��b�"�<�ߞ�u{�<�>�',fU�Ѵ���Z��[�+��u� ϯ�y��yw��=�-��z��錙w+�n���7�ַ��B>�!�1��Z�8k�@�@�����w`�wӌ�\�S�]Gӧ�(��Æ�ضy;�'Oe֬9�8q�s�.p��Y�\����g/s��E�7�g������®ch�k
�����W�{����?�J��c�Yfch���.f4�5K�.<,�{/5�bXS�W� F~�aUt��i2�*sJ�������3~�N�ݍoɾ�4mM��_�v	��[_�z��� W��ߐ��j�V������G9���\ٱV����3o�X�jy��D���cK��z<����s�2��d�w���uי�����A^���5��A�6\��9y9�4��m�K84����M`)c��F��צc�Qt�۟�=�2e��-]����;q�o'Mcێ}�-�Μ�K9q�,�?��ͫ\8s�'O0t�*��Xԣ?��a�����)��M�t�2ǂR��t.[�Uݍy!���g�����PL��a���Sg�[�E�Zda��"�*��:3��:]l�a�����X�tC�$��	]TG�^y��a�5�z�q��~�p~ב� @�|��q�w�'���K��.m��h��I� mΝqJOl���`��e/�\�Lk����Tl1���1e�v�7�eٲu��o�j�2�[�f"s��$% g��/�d�j(u�M �lB8c"֢�%'DQ3����i����٪�*'��Z��B-�.�w���H{��!o��=%.t�}9f!���@��*;�!�blL���'����B�T?����S˝UЗ��� ���#Z:noQ<�R�������<7�0*� H
䔗O}��qrr���;�����<�倥�FI9h���y�|���s9��k�SR�[�o8��9��<>�����[;k�x9��7�))�<%��:^���gU^uj��UC�j����E��Y��d_���'O�ʣjjL��%A�F�X��`�`{W�Y8p�Ċ��社��}�˹�z���V�02%Q@+�Є$c�71�R�(��n����1<�9��;�Wb�/6v���r���o�Sh�BS{OZ8���7��y9vHU�ں%�|>z�,�	��r�I~�V�T��~�(�HQ���R'�A"!���F�K UܥM'��#���zp��u~���'�C�(�|^��Rmgw�8�����a�1Z
��.^�OgPd2M�lm�P%����l�`��d�@NoQ�-l�{�obI;5Gρ!r_c���$���G{F=�4��oy��n^�An�jڰژ��ȗ{h��K��dꈁ�l���Y�Ԝ���b����W���>��۱'��2[����0�#Y�����|��7�z�'s'L'�ٛ�>�t	Oц{�&�>!�(##Z	()���O�x��szujG��9-"c���>~ᴴv�!C��}z������G.]�N��
Tt��� V���IY�J]��ڰ}�*������wv��#J	T�5!�.RG���O���!�ص]sF���/�#��J�/�ۘE50:�=�3���׫N�^~�y5��g��n�-��o�H��:	0��򡱻�)��zJ;ِ��ۤ첄ٙ��91��b��r��{(}�����u��m)ZGO�{�"�WZ{i�C���˿
?'��3�.&6Z�>���<h,mEy6U��^4�w����@��P�"x�Ǥ��+�6�tv����*-��M\}�'���7�T[14�9�ɷ�S�9�1j�;�du�"����Cس�����px�zΟ���[8}f���-��?�K��ws��6.����[9qp#�d��>���G6j�9���r���;8}z/+��cl(Yπ!Cqc�c���+����BN���/F�$�jv䋼^���5��!/p ���1�i��6I�)����D&�`"��̫��������C�>��l�`S[>�MD�Q��Z�:|�����1޷����2s�r68��78x�<;������������<u#݇-��q��3z#f,���k\}�?|��??�������C�w� �Pc�j���lݱ����[E�Ғ$�ދq�>�y����|;��ٴk�-��A��U�8Z ��h��u�hLe�=�)u	f���������yo���+�� O�W.*�V���~Q)T>���˻ֱ��� ���G /�'�1|%�S�2�{2]�}�.�`M��,\�Y���cfnyAh�k��<yy����'�4��7�l|���I�Pt���0�M�q�1,Z���w�pf-X�ԙ�=q�-c⬙�\���h�'וl� ����ܽq�'nkI�IGPت#���a¸�̚:���G��"m���s�X4��Q���e�$��1L܀.h>^�л��ܡ��E��5�خ�U��be=%������4]|G��6ym�:
�u�<z��v��qR��{`�3�:�0˙�N%8�Q��N�$w���Lkɶ�|)�,���C�.��,�2��A��A����a8����a��t�����{j�;�fȂ�,�x��]�X�n+3[v`�(Ey�[O�_!��ؐ4�\b�5�P�9��p�H�|a�a��? �\���'�-��ĉ^�9�i�x� �\o�ߐ��֛n��!ǬLL�1#/:���aZ�l�W��<"-ꂝ�\%�����
�����\��LS�y�6D����懷8ѱ�DGGk��O�*���7��Þ��ӛ�ߞ���<�UR��66n���uN����쬬,��4����?����!e�����*Sy����ʇv������$&*B�ީ��jN�ZW��3���kC�*�`9�i+^�y�f�D؛��hH���"������t�Գ���R�7�|��٠z
�D�
�EѦ�h޼8c¥�j�w���y��CW���r+@ IgAuCKj{I�KG��,[�i^�V�~ڐU3� *Y�!���ڜXQ�>֎���9�ყ��6�0:(��@��9����㍻��b�CH�w���@��`l`����m���~{�%���]j����H���y�^�#Uryӵ?���i���<u)�aInN� K��s�B~�1V�n�t�ʹ3*f���+��d^����8V�+2��_�ٻ�!�ߩ����7�Һq#*D�Ҽb:�^���h(���;:�a�\m���OV��Z�գm���Ո��qt�׆'U L�����S���,�2�D� 2�Ԑg���8
}���ՠ�??�$
�~~��F#�Ғ�N�O���a������z�r�,�|���;�P�z]HA����k��
�3m\	����x�x��'��!#H~�XG� _z�D�7.���ěR5:�#�����_�����jьd++�Z;�'8J���N�� s�ޒ�����e.?Ϟ�{����y�g����~!k�4a]�,jӋ���pa�D��<��ᗪ�R]�$eR*л�B�*屮jvW+bnS�5o��sf�p�$v7hϞ-9��͇�
|���l~J��J1$�pmK;G��;i��+��ߔ��ړ��#8�p	[&Mca�^�M�J+�/e�4s�gdNm�g��;�r������il:��f1�� z%eq ����8U�&?Ǘm�11�"�)t�ܖ�7���G<�/����>8˭g�q�Wo���\�}\��w�r��I�^<ĕ�v�(.����r��_9�����s��I��<��u�8P�u���H� sϢ.���`IZ�LZĂ~ch�C��N���]��z��<���+}:�����3�qp�|E_:��3r��֝��ը^�6AQ	�;F�w�ǣza���ڻ�U&t���.<(\�]@?���Ѧ� F��6}�6n�Ͷ݇�/��z�N��ڣe��p����d�&�wbκ�L[q�q�7������_�y'm�ы�\�u��O����Mn<��9%�D�.�X����*��W/������z'0nzώ�h>���ޑr\eD�E&��ʙZ�x�ҎC1�{��5�^Q��A�o?��%?V��/�S����zϕ(�� ��_����/\޳���55��j��:K_vڕA��.e��T���Vr~�7�Eq�],�t�����#�ozNp�+e�W�l��0����j	�5��i��XU�)�WE�+?�Bk3|�������c�2g��72d�L���F�m������-�]���J8-�ۃ{��y���]���[L�:����L�:W�Λ4��'3e�2�[�oF`�S�]���5=�A-�j*�v+�����n��{z����E\K�LM�0Ч�Ie��լ*	�WG��J�0M��%�� /��4�6�)��E�^����8���ӝ�V�IoЇ�-GR�h�M�`�. �2D�����	@�0i�\�6Dl��O<��3�ϛ����T�o6�����y>��a��,^��ً�1�YGV	tmu�<ysG���p�oc=tF�ڄs�*��Μ5v����j�)QC��g.�g*�����LN��ȁ���[A υ}r��C�a1��^r���W��Tw���0ě
6�����'��
pFٚ��J�J����O�DG����:ȒK2,	�x��U,���D��㵠c
�4��R�� 
 gW\~�g7Q���+Q�J��r�R����C�n�&g8�7{Mll찲�����_��)���� �\ܕ����&����K�"�!T�S�GOݫ����6>6���P-�V��⩄Ȗ�ڪ��{wy:C��D�!/Pk��1.�my�(ֺxsJ�\�ߐwZ ��? Oy��!/^ O�ז�Z���%�g:~�L�z`&c�i�w��;T &HK �<,�\}i)���8{���I� I��4�����3��v�;�lE��17ӆ�C����*7��gice���TQ�I��D9��*���7��A�mZ�՛w���W�>���*yp"�g�GB5��,�Ϭ���J>�m�~�����c���0�~ɣ��?p'�O��L�U�i�0r1n<����p�6Vm�eg�¼"�^�b*0^oOQ`˦/d��=�/-�y�|R���������0�������L��ׯKWΜ9�y��ΚG�\�%V�Ux�6i��[ ��3�l��g1�eG�����-;�Զ=i�!Tq����X7���Q�ɑ[W�f��N?��C�)
<C�%��]޻pm�McK����d`�n��Zǁ��Y8o!�D�W ͓v��Տ��4w������ߵ�Ā_8{	���#�+@�͆�f��
���P��E��)U|<ٹ3�Ob��ԯQ�Di�U��ɳ����@�O0�|Hp�f|���͊��(��qt�}�]�_Z��锩R7��k^o9�o���p��� ��k����)��u��ZƳv���Ih����~'��8�_�ϝ�8�[ m;,��Tּ�*𢇅=��5�]/�hvͻ�/���+Ο8ͭ�xu�/��c���ԊN��W�G����sL�ݛz���
�O����w��e.l?����Vz��s9�:�*׆ɋx�| ;k��@��5k�>n<�ϝ���=�nX������G��U�۰�����t)+�,d�ֵlް�k�Q�v���~�2�nY��c{ٽ;{���?yJ�@ݴy;��M�.t�ԓ�L�(hCiv;��hõKz��IHU�TiG�Ꝉ�]y~m1�넹oL����"�?�
�ԊV8����R�\1��qw��������.���^�AW� V��a��A�/U�I�&3q�|J��a���E%[��`Sf/c���,^��}�.r��5y)޸��w�������	�d���~��������[��v��1Ν?%����WP�I?̜���W�{j�}���\���6���Z�<�(٨�@^�i��ƻ�qZϿ��}Oٸ���_cܐM��1�;1����ry�彙����x-����K~y�+?��A^��NǇb��|y�Q�|~'����|��O�reo	��ՠ�7�M�5\��K���� o�2mŋ%�3X�k���fơ{�zĔҧ�uQ	��k�g��	����.`T�T�9t�`VxHh�� W�(�X�,��lˈ��Y�~;�LgĤY����!��{��Εƶ���c��5l?x��/�q��uܽ���?�����'P�h5�N_�x�Jf���iSY�x�4ġ�������0k!�&0�#��]���6��v�[���`L����bj苩�F:7)�7:��$��ur�_��~�t�0��� O�YR'c�`����z]��u��uJzO]��{O9u��X{9p�K6�bc��.�$��(~��H-��Z%ü� \�O���2��Ʃ� ��`�\	��Bj������6g'#��a��)d��������9�V����|�dd�{��9c�A�QQ��
Z�d>+�<k�N
�����ɮc9�n<3�3�y[����6~���kõfF8�T(���lF��HZ%��bk*���+\eeoA� �;�=ٍ!��W�O���Fy�l'J�	wQV
򒒒		� O����(���悳��~*j���7�2ϙ�������U5�-L�����'O������昙Yh�O�S� P������&��
��5�^��a���B��D����ۧ�����Q��U����XQ�꾣#õ`5<��F��ks�,�B���zcm�m�V��B�v�U�`!���Wsɦ:&P8oa+u�㴡�S� O]��Z��SC�Iz=y��vSg�8�jA߹�p%0�����8i�"�z��|�w�����}j.W}Wj)��P2��Lp6ӓĨ���ڮ���Ox`p6v�Z��[j�*@ F��L��#�Ǐt'W��9��4�]���7���\�؃�	EQ'�Wp2�����1\�Q|��Wp��(��G/��>���]�J���]8?%k�������Ù�|=b.D�q�� ���ؗw�����]� �ؑg�J�*5h]Ԃ���O��u�k�8S��N����H�<�
q������7�eN>��蜐I}'o
l\�(� �"'8��h��֡a~=c���6Q�?���
�����.��D��r+U�o�^4�אj	iT�	"[�N��7M�TʓzR�D�1q4�+�[��TϪJ������]��4�����6�T� /�
��
���E��¥��Hk8�QH�S��@�vw�~��:b�ծP��u�#�Ζ,gw��4���"� �Ʌpy/r+U�Rv61ᚁ0�Α��q�*(G�6 �c��-����bN�����eğ�〙|:.I�}����Ws&��F�@H���mL6_��o>��=��I�W,X�C@*?��f���Φ*�ևV������j�=z�7��E�>d�FSP�*k�,���/�o$C��[�x��7��ЅJ:G���r��!^~��	�{�ܷ"%����G�1��K՚q:)��:�Y�"�g����L�ڋ���Փg]�2�Ab�����NTl(A�>%�&��GHx))	��E�s%V�srb��'j�sYU+MbR*���ZԨ]�z�M�*IRL2���Q�M	������1�Y�c�@{E��ѵr�}j��h(��=��]1��>�7�!}1	��>��ZA�[wR"�ȪP���b������,�1N5c��]�	��X69�e�5y=�m0���`U)��1t�,���L�a�5~6;����ï���5o���~�齶���W�9w�$[wlf��5�ػ�#��^�ҭ�9s�s�n��9��������3��IH\k�Ħ�L�v�V�P˫)��<y�/bTt��n'��9�}Ŏ�Ϙ��6m�x���6`�o]=Y��,�͓�����x��7�_��ߩ!Xa�O�����G���VN�Y�����G�������F�����ʇ6��t�@�+�0؆p/�6���¤���dS�}Z���o���cF�x@P���bUC�w��:_6'���ć@�
y��,Д��I*涙��tc����ۼ�I��3p�$�����9���D��"�\b�|_�� �_<�ї��}�2o�{!,��3ϳ���cg.r��)vl�̒���=i<��,g��Y��W���.e2�EG1���j�1�9�i�-D[g����F���M�040Ӕ������B��d��j��.D��}FW�ڢ��<yI�L�E�l�����3�������L^��_~� ��Y��˜�|��^P��h��c.�4I��a�8��*��-m���P���f%����^K�{�anS���Tl4�F��v�Jz^��n#���RS-^q;���kI�K�2#@����)�WYg�*S7.��pZ�͉��l��9 :�2��(���Z���<�����b��j;��A9"J[E֪<y�Ml4��w$Z>�9y*ߒ��V����-'�6ô%�T^<7m�Ԃ\QxE1~�Ȝ�j�캾�
�������Hhd�tJ	ڼ<��& ��i�p����	�����7�o?<|���\z����{��ꈙ���������@�VU�7_
��V/�<t&���Ͱ�����J��KA[�mq ����мs*Q���s3�܃W{k�\�q�7���J��s#L�,&���<w�7̓��OA�Z�6..F�o��,���9##=��fx�w�K��� O��A����S¥�*(FAvS[3�:�r�яk������n
�o�9y^q�M� O���+����
R�)��Z���"��|c��}����	�Ka���F�-�����E�-j���7Ew]���yh+qD8�Ѻ~�!�����$u9�ozw�,�܃���}���N��X;��!�.6&���D�BH����_EA�4�+6��U
�*�ߩ�$�R�Ǐ��������4�s�O�.5��oA�1��:��R�nAl�ܟ���rh�x����z��;QT��$s�S�kF~sI�Cc��Q��Z���6�E5�ɐ����J��TuGW��U�q���\|��ߩ�zt�MA!�#��B��x��yQ�Z^DH�$88Q;)�F5kP�VU�WH�����-��H[oj�xQ�ُHk�#VX��Z4�e�|m�8��\[�&G �Szڦ��"P�7!C�o۬m�7�aAmR#��(��ި�7U�]�c��6T���Q�\�k�P�r&��qb<�v���O�M�;��F��T�@�:թU#��ٙD�xmnA��q5;g��y�$��O#�M���ԮW��:9��^��r��;��m5�r������_	M�#��[�h�3��S�qr����0a9���{@�d�o��7��G�~���9��Ƿ���!B
ߧ�d��?]�i/��B���V��
�Ȧ�ܼp��Fu����[���O�f�����n���;xt�}���z	eD��� ]>u���8�Ԉku��a����X����=V⻐�<����9*�i�~bx�K��jdB3dЕ��Oq����GceP�۫���.Y[I+�bk炅�#z�le���^t�7��Ǝ�L��>���ٜ�����GP7�"M#k�,�I^���u*K���c�ޘ���з:��x���P��z��Y�J�YT��"JmG�0,"Z�Pk1u��'��Q,�ƪ�"�#��Q��z�`ԤeL��B�Ә4s&��Щsܸ�59�0һ�>k����m����J)ټQ���Mk8y�0������y�U;ϰ|�9V�N��[��쀱�5��SR|
bSP�����aPwOY9�]Ǵ�M"z��ߚ/�r�-[N>c�������s3���	,p�f�k8K��Y۵�yϟ?���ۈU ?���H�u��3Q�4�7��UL�Aj*�j�����>q��NJڵa�@�z�C�K�0�مpG �Ɉ�\����ufP�{��f�B�/��)��o�k.�W��'��ҧ�Ũ�e,��c��VF<F\�v���ѝ������y��?�y�zO��7kk��غ�@��^��5���w�z�����!ۍ�w�r})��d���۾��g1w�D�X�`������&���U��r6h��9bd	|*�q�(Vi�vf���i^#C��KL����l14M��Q O��B��,���c{�����C�>Z��j���YTG"��{�K�g�~,�2���[޿Ǘ_>����|�΃�c�T��1H��M&5M�7��.�7�V+qk��:#��~]�j��G��C��g�������s�exJ,����ڎ��;r-�~���U^<y����bXe��YsO�{r��U�PQ�j[���oh�>#;�Zs@��p@�ʈ
��=�=�F2C���#{�)O�N����Xd�B� ��tfz���hAOQ:Q�t��GV8����8��i�a`@��O��9�bMX]ư?�ܬ��W���՜<��
� OI��5-���]��%/V����������-���OY�<�ٳw��A��I ���
;ͳ��FK(O[�|:'LLL���6���5�+��YhP���\o�����L�-�R:R=ks�k��}I�#1:�̌*d������S��,�_u�J���+�SwL|�fm+������U�%0wOo�0�4��w�U �R�dSz[��3�Z�$�<�v���䖱=���w�\�@�m��x'p>L I�_���6gdH��u��y*8F�v�7�P^X�O��+0�Ȟ|s����& \����/�_Z���\@��ށ|/w�|2�5�I�N��bl�Qą�a*��J��]\l�q���}V�n�I���#i�@������/	9|�����~JI�sd>���l�U2�cx����	3����6�?{N���c��IWN����a�a�5�Ʒi��U@�ua��ȉkyX�)���� �U4g���؂a[�Z�/�̚xs;�T:!�M,	�����ٓ(^0�����(3�dW
}�ɵ������b`J��%Mrk0�/��Ψݩ���K�w�%�Ɲ4q?y��}|ԭ�Fb���b ��B�����<�b(D�Yi���O �_���ڗ9S�нEcTg2��eJW0���D�@X���U*2vp�����h(��R�s�IP�g
p(C��̘v��=�/S&g��QT�	�g`B���
�yx)��DOvi˸�Ø1y$��b��OO�S �6O�6�9��u�QN���j���R���@��ܖ\�>�}��m�R^��ό�L����:P��o/��ɩ;|�p'���K8
�I�]��w����P��+�Ti+:�Er}��_|��4��~p$���ݗ���X 7��q��]��@�E #r[qI�p��el�h��jxV���Ѽ6�n��ɵ��ăWV��
�̉�j�6����G`B������^ڰ���ǿD󐶦�U���7W_m�"����v�n�K0�qpӶ:�t/S+�[��X��c�$(��b�L�3�z�YEץ(���0s�?!��O$Ht�[!:�=[��4�jN��|jT�#�{V^�X�uǮv1z�ZpZ�F;�ȚKT�dj7�e�h�v #�-�̅��{x��OTj�G<~�R����Cǎ�a�VN����g=i.�f�cei	7?�s�v��F[tE��K<o}g�B�	��W#{��eL�����`��vbX�]��^�}��B��]������e���p��v}â!��Vu�
���by/w����-�������}�xȳ�')ͩ�y�sw�+� %b�k"V:v�ia~��Y~��o���.��Sw��X͓���O~�oO�{���S��t�2���Ú��������7�*����+&�|�_�w�� O��9̪n8R��00L�̦"q�ݘ��;g]�&L�ͨ��<v:}��g؄i�\��O���4�{��)���?R�:΂�+Y�e;v�e�Ɲ?p��k��|��K�:b�LQR�tQñj|H�N�RQ@��lj(���A�X3���{h
�@ Hm�������t�C^m=�/�<Ô�e�<�:�u�/�k�QX't
����h�����������;����~���q�n��M1H��.v&����sl��K�;
���b]E�P�����E�1������t
尅7��b)�<��cW�"��LK��r����&J�X����cF�z��۰Og�n#Kvٲ�XD��Ʀ�10�<�]��/��ȑ/&���HF���G:����v����FzJ���g�F��T�0ojeF����d�YQ'̒.\�_ŝ�imM]c�Y��6���ZG7s��%��k�Y:�h5l���y�T��J��A�_ٲc
���yj*g^�~�~�x��+����O�%�3TC�*U�汳����yI�Mp�����c㈍�=�XY豷5׆^��쭱�q�q��\��.�@�������P�,0)�q�$40�D����T-�i��U����іnӼ�>.�F*o�����@�ܻ��*��(��bik���=��A�xzI�6� �_����Kcc͛� ��-ǃL��T)Vt��3�fe�F7W.[;sI�Qi��EA��^��EK�P��3�-%�~��1��:j�w{����ɇ/Š� �8*��:+-(C���HSc+:�i���b�,J���5-�m�_9���ӹM+�c����$�VUl,��6dmdN��a|L�64���FzzBB��j�R�]8��$A��@�J{���M3Gg�C������t^���uR�V�JD&��+q �
�������������o�_�8�r[@�zذ���u�,]��3�x45�+�e[��\���'W_�a�j�W�2��I���ER�[�-��ط�e�&�቏<�Di7��	��Z���NM�p��^�?<��+G�ؤ.ّa4��O�N�v!Q�����MoƘ��t�8W.��գ�+��<�*p)[O_1<��PwW֮X̽ۗyt�
�L�#��i	��X��[�h�y��`�x��	�?��1��2ǈ�i�@u��
��I;Sy8tiυ�Gyp�n]fH�NDXY$�AE�d��D;Gm���V�&��ҙ�<�}�緮ҺFu��&P�+�@[gR\\��!���s9�8��\�r�u�����hvGVdO�"^��ī3����Of����=<;p����r��Pv�4dS�!�p�W���h��\�R�Y9\1�g�N�u�F^�xȓ�ۘ����Y�e�i�ț��-ɧVhi��-��. �M������_{���p��m�;��)+iW�1�E��hܑ{�1��1T2w�eD*G�����_r��tN�ʡC�x����fe��G$�7o�C�&��#��!}�Z��2�'�:��=x��]..� =���9J���]�m�9J ��zb�,�����5���3ȳ����)�{�>8�S�0k�$���:�P ��T��y��i+]	��}���Z�m��1rUs��h��F�zm��m@V�|}�
a�:�:�1.8)�!���Z;H�|�a��0h�*
�����ql�q�{�r����8�ν9w�6w۞}sX�q3�.^c硋�w=�Ӭ�GMg��L_�����۪?�`��U���惖����m&��U0R��-��5�����Zj�� �VN��W�ux�e��$������u�g�z��m/X5|/��EX>�Dw.u���-�`m�~<}����<�;W����/1���L�@���X�8ڈ��rz�^	~���?~�yAK:t�X:�2����}�Vy�j�@,�K����`6[���B����A����W�����{��$k#:�fK"��%�vgf�aV�ncƬٌ?��Sf3n�|�Ϝτ�B�p��m~��;�|�e鄾�M��ݏ�X���k�s��-���M۵$�%���x��-*a���89G�SgL������V�/��Al�v��i���_^/⣃13�kQ�j������Q�<5\kl_G �˸���u�(�ߐg��I�UC�ֱJ:c�}L7�����d�����|��^<�͑C�y�ݷ,X���v��1NS�7}҄���-��h1�y�1	�+�DAѵ(����o2p�f�<Ƽ��̰p紭?}�Y�c*�'�������9KG�ed�j;/N�yp���cb�)��Ҡ�����o1x3f��N��am�ҸL����0-{�^�$����MX-�l��$��T7m�Q9fbn�������E�8ɝ�l^ݎ�=X�4�������b@�-mmtt��1�߂~�^J]�K��� �9$b�+�S^���-���:�g�����&������+��(U�<�5����]γ�;��N��� '�6u�ԧJ��$U$�?G[7��Ā�03֒ks�䳽�wn�"��"�w"�;���H�T�L�F�(lЄȘt\��<�@�<��4HIMJ���O~7=5��
)dU�@�v-i׮���$&&BbB*	�����k�<5\�����H1�\�.��O�������t5��g�עj�,����z�t���u�(�3r������U��|�^��n*r��`��!�LԐ�\��T@Ò��f�		�g ��|����ʌ���V�h�J/mav�ٿ�{���tu�c���ʌx����o_��vJ�ܽ�!�j���p���8�(uMXh��<�0��Wiu��RHI�'��GKّ�Kn�UŐ���Ę�x�H]����Xޏ��֬�t�{묳�����ڙZ2,)��ort�.�Y��N��	�!<�/�}�Z����Epx�<��~��縶�$N<��ӏ,��^�t��В>G�ܺ-��3�>���'��۩y)#]]	�6&m/�̔Xwg"|��:a����#O^�C���mI��͈��5���Bڮԉ�(�];���_� /�� �r�U��]���Ovr!Lڌ�@���kW.����D~���d���.L�1�vZ�i���]�T����|.�[4i"1�΄�%�y	�Z��"m-D�Sݟ>��w�����]:�# !�@��q��$z�=XX��Ή��废��x��!5SS��qr�xU��::F�j	���s��j*��SKS����-����A���%[x��{v�:ˁu;���{�yB�:��b��@�ر?=|Ź%%�����}s�6|��-CL��jS��yă='����|����sh?��`�[��޲�{�X ���BK$}D��'�P2w+�go�˯�SZ���1ը�@C1p�����+��s��.Y����@��$�-�ŝ����|�'k���b=��T�s�㕃_E�q08F�$�ɽۄI��M3)�&�&\�A\9��� Oy�๹���n�<Z	`�;�`fk+:����b�-��g���vXE�N\Ĝ�Sh.��>I /2_ �&fjŋ6�o�k�ךxw� ��o0����h��s5�"ꑕۙČF'4�&�=����+������ �@�i�s\����#3V�u�nl�w�ǯ^�i�V��d�&��϶]�y��N\�������/|ώCWi�z�[����q��7�VR߭Mg��-����1��1l��N�2(�CU�t����`�����������Qt�Nb��2����a��.��/3��{��z�������9kG�IV?^��e�"�D���%eѵ
�N�x�/�p/>�E��\�����az
7���%���q��W�}˯�r��6voK��ެ��e�@�
��F�]kSy�&.����ll���_�c��L�s���2a�sz�D�֮-Ы#�W�v�U?�I�˘d����%bn�ADfk��l�u�5kK��n�e��b��)a��U��R��g�x��1��J���)�|~���g��|;��ɳ�9}�[wS�f-3�N`��9�)���A3�s
`Ű�L<;]�X*BWU@��N��l� B���g��*:��:��DD�L10��ؼ�v���4�<�5����<x6��4�N�El{�b�c��}h;�zb�1�̞�^�S�������y��6'���7�2e�&<STdnoL*Jc�� }�)�&��K�u���4Y�s�x��Yh}L�R��KN�9������3��(��RYcl�.k/{�1��F�YNXP�@�XaF:-��U���-Yn��a#'��8b�A�^��*�V�>٪��=���ܩ��mґ������l�>�>qlEsX a����rN�Q�+�؊R66��X���P�tB�h[#�q-��<��&��_�FT���l�̠��;s3tLO3bP��6��[
�y�iJ=*:���m�X7w'�]�a���pm����_���,��j����
Ӓ�::�����X��*����"���܊*b͏Sk�B�J��C)�b�{1�)�;�U0-02��s�,߸�$��T%/�:�נyQ.�ge����5��M����_>��t�DGk�8_�@�նU;�ʰ~��7m.v�t���A�&m�H�H�8y��pXER����+mluz"�|���5��]g����VZ��J��V�=�ʙ��*/��;%*��ޚ�nǥ�o���=����d�V��I��]�9sGNa���\X��[�s?&���!\���t���-c�ҕ��^��m{١�@�#=9���x~��H��VNL�O��3V^�Y���)��($i�V���Yӫ!��H���}%��Qe�u<D�	P�XY��M��D��m�J�Ѽ-�Ϝ-����O��ӛL��
r�\i��d���'v�����ʨJ%�?��H+���q��ٻ���C鼕�v��}'�n�Zn�A��=I�t���z��.�c��I�����~�U��`��-5�U�E��1�!�*%��ƍ� F��}�5�fS�rU�J�T�.EYG�a�fc���'�v��*�ƻp���鸙�i��q^�$���͑MOM�νۼ������E�;���@t�?Q~��!��H�
�w�ڙ~���o�>j)5���r @쿒2{�D��X�NZ:�E��J)T�?x�͗4o�{�	Q^r�ў�Z����5~�۾���������][����҂Pww����6�������7/]���R�wL�7��1�b �;������۸r�9��PQ�����xx�%mr�S �]}�#m����K�.�@��k�JJ���ؼ� KW�r��5m��%;�(X�����P*ԣ�!��6t����O���jU�Ɵ]yH�*ͨ�ρE������+M��B��Z��ʙ��k܆���\�،�]�q��P>��ě��97p?8śU�9X�5�ê��s/�y�������Y�"�F%�W�y
ܔ3C�2P�(����s��O���Q��A���Z�i�W,F��(鳧/c֠ɴ�ؐ�U[�.�1���0�T)TZ��z���@�A�1	�Ex�bE��t�(�Vɓ��J�f�Š�A�Ө�`���j�X����5𔖸x����ml���[=u��{v���Q��\��S�v�	��������Oq��7,�|���73a�j�Kߪ�z(�ߑcg���K�]�����Yw��z-�%�!�n5Й�����(c&y�>�K�aXx�1ir�֏ѵ�����qG��|�-��3��+��U�޼����t�z�G1�%���{���n��o\aw�J����Vr��b���O�G~�A���~�Y�x��wy��г��B�(Tyϼ�E��:�����1}9��cm�9l鵛�k.1e�m6y��/�O�ߐW]*B Ϩ�@^��J��$�7O�3�.��f��s̖����̚������Vi�w��e��z�Y����O�M��o~���J�$��N����c�ض���k!���c����ţ��54u��>�̙�4;�Iͽy;�e���V)iC�9W��%\=����TD@D<Cw��02��ȶ@�<��6e��TtmLL��k^<���X�w�<������N�CZ`���A�vd�4�_��_>���������_����[��	]��*N�,s:&��L��i�hmY3�zӰn��?��k��sE\��R1o���R�zwZT`���Œ�e�JOi8ûN����D��d`��2�gb���M,Xb��ag�
�hs��ܺ��08$��AS[���c�LMY'
e�g8��u��x6��j��؄�]#�N`c�މ��^�4��~���?Q��iT-��]+s~U��o��u���_�m��%Mx:�.7�&syd*��f�,�'w�P��"���$<"������cHII�c�xx��OJF��$$GS�R��7�f^3R3��[�Ԩ
�yG����(*��H��5d�0�V-;ҤikMT�Y���
����`mXTd��jS�^��b���̜>���'P�fg��m�\z�iD�U�NN�փ���LVj,��d6$��S�èv-صh>�ӧ�y�.��Ʃ�k(�:��zӭn�+�� >��H?�E��H�`��H���l�I��i��̩5�c���"���N�Zzq�܅�6G��9-�s�ЂFfZND]��!�7䥋BUôݪ���K\>x��rr�8p�Cǰ+2�G�G����u?�gͣX ���ܽx���)����L���_�mX'�l�Fߌz|�Ә�inĩ�2�eɜ�)O��Јp�B���.6V����\�lD(@P�9#.����-V�������_3jv�T5�����m��50���%��u��rd�v��dl@]kJe���ω��Y2s	>A��.��K����X�Hyw2<���Y���9�a��Ў����W3sc1���qs���
0�9��jۙ}Or��e�/[C�(z#S�]ܵa� 14������}��Б�kشm��N'>2Q[
0�# OQ�>���xyɱ�P1 G�e�1BVQԪ1&z���
0�i*z=08H�R�R��g�`��u�^��JUs����)WhP����e�g�0q�d�-]Ƞ��H����kШ�Dݯ��y�x������ciڲ���q����Ko�`����&X�ZѼy��m�S� �\5-��ٗ��(vl���s�H%J�Ÿ6�x��{N�>ƈ�ͩf�O���ܺ���3WRY�����u�ͺ�s)]��#Ns��#v?�ɵ�`�V���BpUH�g�C0}���yhK�5�w�KHw���Ԏô��NC/f��Ǐ��qq��Tʡ��7�u�VbPio6�T�}��x3��Ij����t'���x��9|���'��.e�w& �����x`)F��@ζ�zʋ��!��w�<u�蔔�C�
����׆h�X�;abi-�� #=�Do,�[m�Mit��X��a��٘~YmiӐ
>y��ڠ�ꀡG'�=�b� ϫ7>0
�q�0#��6]�D���N\���:j�Ǹ�)�Sf(b�Jt�i�f���l;����Vq��1�}�5��(�б�+7�жw�|͓7?k��K�cŦ#o;��g9|��]����ܺq�{��pV�#箱v�u*�I�,�0��D�OD瞏U�9nE�[�W�s^��5��a�'�:�o�wW ��m�mV/>
�P}`P[=�X������*������{�B���tod��@� D���?TJ�~�����E�㯿q��͓��/����ȫ˭��]��ey�)�M��3��e��4��{]� ^C��|x�O^��՚�݊i�
���(c�X,<�i�i�T�y�/,�W��L���5��0w�Z���%�뷮r��Im���?���,\������	���Y���Es2a�8ƏŒ�˘�p����oZ��K�2{!V�Ojf� �)�Y�d�y���Rq�wv�zt��wnZZ���硳*�<��6ЩaZ�ض��~�P�id�DԐ�apS��:hį��L��s8v���ܐ�������F,�փ��������T��S0J�e���+��7�{K�%��j�'R%�;���t�a�]�n����%�׮�d��.&�7Q��7ȓ���T�%]`��37͓�Gˋ�� O��M�X7ܭ��c��-3L͙`b�l�p��4go��,v�c��(>9�Tg�*����j#sV��j�B[�[��U�seY5#����Ѧ"��r|Qsol����rC3�)i�����bUm���,�L�
���p�{T��ID����3�^T�Q�&�
5تR-��5��o�@&������8{�Xl+��[�ş>s#�Obp���mM�Ju���K���t��4�欢t�n�/�@��#hѼiIY�=�]6ӯ[7zu���у�6~���g��)Ϛɮ%+D1l�J����U+1,�"����+=�a9Q���O�������k���>x�p8�����\�ޕ�Zq||S���Ϧ��oɺV��)
�da�;��83!S��j���bΘ,{�Ř��SGsW3�[PhoC[s+�8��O ���J~l�9#mœ�x
��-�]��W���3��⩵e��.���K��QH�ΒQ!�0z:oW���UWn���۽���T7i7aR�+�O�Յ{�i؉/#ӵH�ߒ
8*���ΎUjs��E��l�i�l��Nmq72���/7-���)	ӠO�MT���N.f4iR��S�P�ru+Dkk�޽{�J���t�����g�BukW�lɓ{/0ѓ/�I��U�}ؿp?=����ѨJE��뇏�6l4�sj����}�
�1}�d^^{�H�d?�͉��"��;3'L�9���FhX��m(F�
�Q�y���F ���3=�����a��B8R�G�<L�����5V��l�<05��T�)7/_L�}s4��U��Q�LM͌0�4���N�
׋����q1 �hpm
��^6�L%�3���F����9�`.������z�-�My�ռU��@���M�?։�_@�r���곹�K%W�E*�M�G}gjn�M�Q��|iq��a`m������	pk�j��ɳ3�����7�#�A�l[X��#��SВ+z��=p�7��g����o'���^��%K6��Y�f^��������t�>�ɕ�l�u����<�ؤ�S"�Gf��X�6��ͩn��PoΨ�xx�6�v�o�NT��<�
���ۯ�c��]b��e����x��=��q�~7n�iǽ������O\��ASx�l+�L^���l��D���/]B5��*$��	�����Ft�WjMY/_-�BE�Z�8h���*r�ΪLĕ��վT����U����K3�2��wȳ��m$�gFk��@^�<ףy�FϦG�"�WiKQX�^�:	�u�ģ'�"j�Z�O�Fb8]`?t�}e;
���;ga� ��k0����ʢV�bZp�Z���͂�x���Μ`���Zƍ��O�n���ZL�1S��tG/�bױڪP�������Ҥ\�s�=G����I
��>t�(�O_b�ܭxE7��*C@/]$��v�5ل��tN
]���%�_���-t�i��/2G�b�������[��Zw~	�ƾ�����E o�w[{|�O�����|�~����a}��{��?��'��|�O��z�ul��;G���[{�J�<�y�}�5�{dʍ�Z�_ f����Υ,Z��h�7n�����B�E�n���4�h�gi��}4��ڱx�af�4p"[6�g��D�g.bǑC�||�/�T�����훬߽��{�K\b��=,Y����+X:os�Mc��٬\���SW��/b�U`]\7a��"FU�����֥�v�Wb6��>����2����cf��޼�H-L�4�3�m����ERW��Θ%v�2�����N_D��4��&j_��H���UFaә����6l6��ϡU��4�5��=�W��ѥŠ�4L*NƼ�$��eõ)���3���p,��{��Ʀ��JjL�DF6"�4��)��M�N�^�R��p�u����8�X|t�e�'J�C:�tS�[:r�x{m�im�&G���sg[z
���ٯAoъ��YQ;��U��D�d�9�1�҆%�F����h���Ȃ��vL4���(�"kG-q���1ՒbhZ7��Ѵ.�dV�*lW���j�/7��-�x��*/J��zcW-I�����)VK���$[Q�j�)>.�N�[2rh�v�HC��۴��捥\�v��5se)W/��ճg<z�ӇOq`�Vv-.fސQ�j҂��kѬN�g����?u�Gg/�m�R�vhG��ήĀFuX;�kF�a��N,ܚ�S��o��ނ=�X٧#�G�c���m�ώ���؈ݲ81�*�K�="�kòx=�����Y�yQk�Y܎g���|aK��*�����X�ϣ�9�X��˹Y|5�
/gT����M���D�����D��ߊfS�rcV�?���fCO���n,8�f��SG�	�(�W+�P8)�Z^��;��\h�@�iٲfy*¶]Ś�<w�S�j����b{o��6�Ŗ��L�ϙ�K��i41���h"]��-X�7r�vK��Xҫq.�
�ͼȒ�Loݍo�~�Q���4 �Ԛ(SOC,�ڐ|\L,�JA�Z�@%�q�(��L���ټx|��M�޴6�_�㟟y��;�}�-�^�����h�هlCk�	���}523���QZGfұZò	�o��֭[|���ݻGzH��m���Wܸ�������[��,��]B���G�(S'�����@����{�R7���*Gc�|`#�3�$�_�� ��h004���)�^�5�@' Z��^`�sKML*5�1���{� JE}[ژc�h��@��F��^@O����c�+h���sv�r�V����;Q��9Cc3MtҗhPg"�)b,uo�����P�{#�K3K9�@h34��I9�`Tpi*�f"���Y������ʭ�70�R)@5U *���:�P��P�X'��S@�������T�����	_[O��o�̓g����\�y��uZ��+�1���͇��~�ێ]��ه�|��'�~����,�4��y	�O�ù��x}ﭖk���9� �Ti�o�:�(2��Q�e]��p1ϭ���{�����<y�I���O�=�q��wo�Qp�������߾�[/`�i�vɡ�S���E~��g�{��c4Ǣ�����2��+�o<���)�W��������s�`\\�q�c@�\�zn�jA���D=c�y�'�H��Y�DJ�)�Scf6���|�V���`����}���S�V�|��f�a`��4* ٭.fn��|�a�'�ģ���S��gʛg�?�/0P|0
��a�m�Zyeѫ"ub�w���q�{�kp��o���L�ٴh߃Uv�z�A���ɤ+��pK�nf�����lcӮ�;|�}G��m��<��K��� �5�_���S7h�~���Ty�ʼxn5p�4����5?�A㋘4����u��^Ǡ���'�:�²�#*	����-�c����-}�A��]y��z��6.lp�`�o��p�o��ţ�y��'ỿ����e������m�	����X��)mߚ����7sg���^����i+^ܷ
�f�X"3�pl�:�����k���3�?�/Ƭ~T6'O�6P˚����?��+��֗p��T��,y�01p��*ۀ��_��5�XU�V[�v������G���s޼���3����w�r�6�_�ˎ=X(�W�����[�?e<�Le��b�^K���2��1c���'0�T�\�e�DWU$s������o6~_`��	����7�N�.��e��dS���6�<w���
虥��:�;���qK؋j�Ud�QE���з��XE��,���\\j�]�	����wfsmi2�Ď$� c*�����fiS0I�I� �k�ƥ�<��,ǻh��l��=O�0ܓ�`�G�.9~�T���;����C�1L���h�Hܤ��_���֮�#�IK;.�زO:�%�>,ɮ̜�BV������yt�W���IQ̻�r��A������Լ1_�F3!ؗ)6f,��|���6o�t�3D1�x� ~��[��ajI�g i�~$�zQ!օ��~�eC�,�N��Ԭj\[]�G�+�bSW5��ߐ�hAHH�6�-<$7Gg�b�3p���1�� w�ͬ!c9���s[��z�$F����.X?n&�-b��)�5�=S��@�-dR�l�ul���=�2wwWL����Ձ���ս*��Wbo��l�ƎΙ�"��CkqfDu΍`W�#3�0�*�f��xA�����_ې��ߖ�o�d��	��j��m�c_k��_��"��.�����~���}����5��|�ՐO;��a[c~�Ԁ�J��q}=Mެ�ɋEY<�_���ҹ:*�S���X�Һ��J��K�-��i�`�0��W�z�S����9�-L9&J󄡉6'ﶉoBӹ�N_Q�)�fTZ�hc[����u{�O�&��L����ʉ����t�Wl�D�VL6$J����9sxu����W�
�)#�s!���vS�މ���q��%���Iz6Qz[��yFX���=RSS�@���""��9�q�	ڱ@� �s�����CZ	�ѥ�~���?����Ox|�On_��{L��Sڤ5��v[P[�k}3{6��o�^�g�!��?�۷��׿�/ �y�.6,ݤ�<S��^?�^8���w�\���cp|�v�H��?�Զj�\5�E�`I)XM��q�|���5���Ū@��L�J��D��� Nj[.
�T�nR*����g(�(o��)1 255��ՀK�M*���`h ����D S���f�V��8jDS���Y�@ډ*�ڪ�j啿-��c�\u=D�\3�����W��74�-�}٪�Us_�g�7��P=u�
���}H����X8k�o���ͯ��ۿxp�>�g�b玃�|���^�໏<�����v���S{O�v�r�����[/����^|���o���^��Ώ���~�:ެ-���\�}���α��g��֕��t�%�.<��'����w<���Op��Yi����s����ۯ��/凟�����q�_N����g8ܴw��y��C�p�	�����s(_:i�w@-�f劯�+f�~�Ь�UY���H�5�[��t�Ս���iRԲ9�Z4�Aӆ�oҀFEM�m��<��fki���Oyg]��ݵ*fvb\��%u�S�W�y�Y��F�4�^��nS�Չ�ɭh�_��Tt�g�Vy��أ��V���H௕z:�nz+�^��b0Ӱ�����X�Q�}�S+^Š��U��U�)":��Tj>��m���Na��匞��Is�0m����U�ݰ��t���e��:t�CGNh+�(ٹs'����;��-�F��-�	:�i��z	���Q����ڲe�M/`��
�MD��ĨH��՗�:��{Fֈ�L��-[O}Ǻ]YR���}K��҆'���yE@�f{GR,:���k|��?�1ʟ@J��:��������,G�|��	�{��G'�e��?���A �=T����"y`ʝ�:<�tv�:�󇱩�Z��d��gl>�'Ϸ����<���o��=�c�eܚ�2WA!b-�a`(��Gt��ŷ?r��Yz|1���q��}���[!؏���g=Ϭ�Śk��Gl�z����D��E�7|(�kVh�5�����_~�U��v��H�k�oTi;���y�1�v��5����k4f>C�;��ġF��1�n��E-�����ljJ�l�Ibg��Ժ���:b��Ȧ�D6�<��!����@Eߦ�=ka�U�G�\�*� �VH&�r^T!�҈L"ŪI�.}���&a�1��I������h�f�a�t&��s1J�α2����J�chc<}�����X޶�:�L����;w�Șq����A,�'����E���weW@��B[��NIZˋp����lX]��#�9|�<�o�c��Cl8��������#n߽ȃ���6�a@/�UHa���D!����Ē��?Y:��|C����Ȕ��]-C+��"��Hp2#�̈́��6t��dT�K;��yX4g��rwY]�MΣW�@�-���&=<�Jсd��R)ȓ��+2��N�=�����og���®�}�1�;+;7eA�|�;�bC���֊�c�qtBSN�o�թ�9?��kc�xF{�h�ӹ��ra'�\ԎW[�fQ~YV��ō�rfML����:�XА���rI}�ZQ�����jm?��ǃ���pS>jG��ɖpV���vp�'\�������}�|��HW>]�̟�z���r\ι��w��J��Z�#�$�lϟ��j�1�^>:К;��|^������i����!����e�=u<Mi�hK_gW����ׅc���e�چӢ`/�Ly��ɰDz�bVs�����r`n���(�C�Wr���6+G�U��Q�:n���Θ�,p�`R��ؼ�'.rR��YV~�����
�w�$G@���+��|i���!SؠY.���Ri<-̵`���D-e�<�Z��)����t*�^��nކ�#FQ19��;���k-1����-��W����׬�<�Za�M64����E�A,nۗ�β[`s���oߟ�{3�� ���˞�r�KY8j#�bh���ܟ]2��h��^��iK��Z�K5��JA���V����@�B[9��ۥ��zvP�\��)|�)S��EA��-�l���?������5�˗�+_�E�}�uԾ���
��//��/_�<�����&��We���r��jTp����;��D;�m�С�W���YE��Z,/�ڪ�UeW��D?�G�{��ү� �O+f͜��x��[Nqf�y�m?��՛ظfkVne��,�̶�[9��8�䫯~���{��qF �+�a���S���m�ٰ��Jw�x+��m�ⶃ[w�-�w��%�]���k�ѧ�`�v̚IX6y	�[��gAS�4l���S9�n�vۑ\�6�}����P��~g3�3y��϶�<q�O�������)X��=�!Z2fo{g,}��)*�F-g8v�X�>��;��p��.���v���Z�¶�;���j�;}�A�SUݛYi+Q(�SC����^�+l=�b��V�L�\�����ۓ~�:��?�$�:e���\K�f��c�=c���4}X��W<;	�����@*z0B��+���Q�AWO��α2O^�U�|��Gpn��J��JkG��������sW0v�|&����u%�]�V��ݴ}��fׁ��>{�˗/s��I��8Ωs�9t��'m�3���]�a1"�4ƶ�\�;���1��� ϰ�%�^A��&y�_�� /g�=fl��G߰v�=��<di�U�N�"��Ht&��Y��T�p��Qɐ���W_i��;�q���������<=}��];�N����7�W.<���^J=NY��)�7B,���/�Ť�Y�6\��MrS�;xQ�� �<O���I,��������,rt>�{�%��:���.LZ�����o�8�=��o^���Oڜ����3t�4���͖'پ�ū6�bI1��-a���,\���/2bZ	ޡ�b�bh�E\W��7a�PG�C��ڊ�UًYui4�����s�X}1qꎑ}l�jó吧7ȳ�,�8�#&=1M�&�&�6��~�X���7���X�E�S��Bt��"Y�y�%��<Q��E[��4�#�1b�D�C�4@� ^�VZ&��+.�(}��S1J�"ߏC�3��I��5�*�^�wRk��qJ���M[��V,q{c�]�h�{�&l$08U~��v���=�=�����8��3�E&�ɔ	3�.�x�*�l��p���6�e��m_ö=9r� �vn�:��W/q��N�8�Ӭ5�b��b��BCs�H�0�И~ DF�0J�N)gS�\O:�Z����%�eoO��+]�����<o�5�`Y�$�U��i�;�����Z�L�aN�(6w���a��݀�jp}\!7F�����_�g�j�rv]��/�}����y����4���B>�y]CXל?�7�����uKC~�ք�;����%���מ����)_oj΋�mx���vu��=y��/w��Ѷ|s������'���p�'���h�j�_N�Ws���E��z1���/2���L�������T����L�z
<��o}!p�.t�s��D�<%���ձ3]D��#�����C�/�Ε)��Җ�Lɋ�� u=O7��o+�7%5���X���N+ΘZ��ĞGn�����ԙxab�-c6�G/�<F��4��l�Z���6�T����Zj�-��h�
���d�|�6��-��1UĘ�b��9��ŊmK�gM��s���O9��q�&Zڍ�2^,���;j˻�{��)�S[�b��ļl�a�3�aÆZ^���_i���'}���¢a#�+ ��Ȗ&f6t���W0�6��5F�B��V�F椛�Q�ʚ����
��g �\�r�"Y (R�{���zg��hT�I�qڻ�#��,*awPH(!a��i�*B�i�WR��QS���FCl��[x,�!e`�OQ��D�������OQ��)*���.���ʡ��(Q��e��CI�����Ͻ\ʯW^��Cy�j��?P�Y��$(8���0<��������j&*��
�P[�<T�~[�F��Zڮ��d�J�<����*��:GP�5�&A��_��vch�f|�U��՛ҿr�'Ԣ}P%�;��9���orj�9�4���qh�M��ZLNo��f��i�L~�8��=��ȁ�^���E�Z���1�6��e��d�R�֗�֞d�z�%��2<�Ս�r�m?n�nǍ��\�m��E�ӄ��.����v��FSy��S����A���}��7�I��������6AZ�sCSͳ�v�&�\�Oמhش��ǔ�-hDN�zT��դJ��4kݞ��/�t�z1<�11����W{mΞ��
f4�G!5\��ڗ�/[��8>z��ddAw�t���.��uл5B�Z�7�@��yz�<�v�����OE�@�m�/8�Qóeɐ5���?'�!���f��aWc1v����j"K���e�a�o`��Eڼ���V�p�r/[���ز�GO\���+�|�#W�r��������	LlY6L��8��D�P�3��x�F'���	x49����C^����v��Zc�3w�O���%�[o�b�]�_ȭ�"��U�H\%քĳZt�4�0�������7ڴ͋��tT�_ �S����Qv��JI`�@�+������ڵe��(�>w�-���5��3���J���c��a��G�p�_O��ٽ�c�V�Q����#X7=�}�-H�5"6Թbm�*�Ey�"H�ӕ��q������\���?���\�O�q����M;N�z�.J�x���ٶ��_f�eFU�
q���s�tB��þ�s	��²�.t�6���#�'ǣWa�/�S ˵+F�1�k+�)��2CK5\[y��y���gtC&�}�a杅�_5̽+cT���y�p��s�"���*����a�9ӌ��ƪ�`t�]�E�$�["�k=���J9W`�����s��S'
�M�"SMLm�ξ*>��G5�޳
����댰e�RMx;�Һ�L�F�t@N:�){Z�س,��վ>W�eC�QL����ӗ0T��9��:�|��'��j�&���qôI�%+�i�
��,Z���&2x�X�/Z̊�R�,+f��q���c�@�X#3=}�<_�*�7�Č��F�����!�:�fT�[i��s��h�nM�`+�'�1,Þ)5��Y/�M��#��O"gGepwz.����|nm^ͯ��K���1li�_��������H!(�]�x�>�_J���������D��xK8�V�e{F�]��0�p��G���p�;��u����>՗o������`��1��oKl(�?�?�}�ǟ����O������}����D���U����7˻Z*�׊���%|~��?~�n�����Gc�|s �/����%�ŞerI��r���W	������P+~�R��չ4��'��S2s��>)�*�N�x:�#5�uE-9ޮ��Yca�=kފ��_��t�DQ"�坳�8�� ;Wm`Z��l4�ǳWro�l^.Z���7f*�_������9�Ɵ���>�gWZ6E���{��?��䲍���,ܨ��K�)bĘ��mb(�[���� �����r�PC�*���(z#QF*�0A����F��
tn߃�[���O�N��g�0�Y;���7���&�li�L;W*J�L�w*Mg�Ь�7jB��YtRˇ	�4���[#���Ӵ)۴fR�N4N����R[3:=*Y�ۦ"ˡIM5HJI#19E�W���+5%]���V�H��*IJJ#-��+��R�������J������R+�KT��J��Ř��S疉�m���}�_��*[B|�v}�F�B�����:O�:G���\�?CKET�r6)i��K"6>Y����"b��D�����Gk���ˣ�����%L@R^x�J��R�H���%�ݛp#k�"R�	#j��KJM��W�("����i�A���Ui���-�X������~LKd\�#�"��$�ghR#���>�%��s"�g��q10s����3��r�.a	���a��9�k�&Q�-�	�����p����)�y�kϧ-�J�A\j����E���~�[̙���x'���X��_!�K8o����D{1L|�\��U��t�򸖔nce�F,m\D7�E�Z��T�ktF�,:i�:��l.[�-_- �C#+�t��)O�?!��Ȓ�6�,2���,�-�9����%#f1�A'�綣n@m"��`���� �6\�O�SiU��t^=������b4��27bZx�_�g�w�|5%�X�m����z�5�����ٴi/�cc�V�Z��k��*+�n�t�!N��˙;�9|�&���]���)�Hi!`�&�$VX 
3�ژV�m��*��=�A����Z�_��E��n`��@�Sm�־�s�{��}?�|�CVn�ΪշX�r67�h�w *�%ޡ�'o�g$�z���{����|�����;����Sõ
�'�4 Z*ȕR{?���/�o��xb)�א�3�s|r	KkgS�M,(�˄4�����	y�.k�\�<���I�)m	1]�>��&o�Ttid�X�`f�#ƛ��zl9pU+�K�)-Yŭ[7���w�.�����Y�a��&O�߼�5��~�Q�l?C�!�	K���DY/�`�Sq�=��0�+�_e/F��4O�a���ư�A���!y��УF�1�o��mC���L�E�b��� �Χ1��]�W�ez����k*����V�η2�A9؇�b�+�VayX'��*��)}�ŋ$E�9��	��|��X�h��ey��%R��WZ�>c.I31O�*`X�a��Ӡ�X;����A�p�����S'�Ll�0��3��!�f]��g�z�\bDQ�k�xv%0�ѝ�+3��f.*a𨥴�6�!SW���Y.\�����Y>{>_��HQ��4�R��[�`�h�Ξ��ƕKҫ'9����s:����0�MZ��Y o�^O?C���d�`���]e�C��mbdJss:Y��Ò>Q����bV^ �[���K$���svL:W'W���j|��:?���˦z|��P ��9Ј���N��Ӊ��u�#����'����+_��� >��/��������F��/'���p>��_�L��W"o��N���|<�=��[�4y}{_����y�x,/�N�������%�ƭ��[��+���j�`�� ��VM��k#��?>���z�&���W���ݻ���rx;��O�����|�НO���Lw�:�Kட�� ����X�8!Pz��<9�P;~�֘'�s�2;����?4������ ^�����Q)�#sfq~�x�G�q�̎�}��@'��4�#[m^��#3����g?j�azOd㬵|��4o�.bK���ZR��'o�/FD�J�雚Ĺ���/3�z}ۺ��ӗ���T����/��u�\��NZգ#�ss ��W3c���=��HIIѠNA�y����w)^@/�+�1d�E'Q5,����dx�* ��P�5��rk�9N��AϜr-](�p���m�z�k�:z*Z�,:���sd�6�4iG����P'���2�CG&��ˢ	��?��
�7p4�>$��$�Fckn�������+�q��W�-S����J���?EASR� X|� a��m�?$U��:V.��n���z�-���Sy��1z
�T��)
��5Vݏ _9�)Q���w+�S�������su�Ҽz�|%Q��ЅG�j�+$,�?�?�S�W.ʋ�%����͍H?o�~ї�;�P�`=[��QNm�7h@˼z����S�>]���d���'�/V��{i)�}藖�^��5�Q+!���L�4�H��ft�ތV�H�����q�;0�]
���2}
�.%�֍�Y�~���9>w�	���g�8�G��=iЬ�Z��Qc�{�8gvf��<[��c5Z��lCx��S�8m^�3���}��N� ��|�  ��IDAT�H����uP�yfVZ^Í�7h+@=�&E�i֪�۵�G�^4oۊ��D��kޔ:M�4��ͫ�lߎ���9+g�=�ul��T�t�ެ�	d�@�Δڜ�����g0�yzVkA5��;��Dy��ۢ�h�A�Oyޢo�y��sO��>y�� OתU�j,:�<�B�(O�z��|��
d�?�y�S8l�0| :�"+��{�Y�ٲ�0[w���}�;y�]�q��-_�ǎs��x�v\�y��8���	�EO$�=kQi"��Ob����3��ø����HC�<�fW5�3lyG �1��o�����S����gV|̊-WX���L�nr_Ge�#0��^!�z�1�5�ub���?j��y��d���2��'��ڝy�6���A �@�+i�o��yf�㔆|9kggn�8o��o�>fھg��RK����L���G�Ǯ�Qt6��w�XZ	���������.7q��m�o���'�y��-S�aڲM�9w��{�2�n��$/�Z��A�ꭱ���0��&�8F`�>���4���ƨ�!L��A�n���>�j	|
�ĔA��W�{`��E O��X�ȳJ�ޯ*��)X{�`瓎�G*6~����<����eT}�3�`��}�aV�e�$k����T��FcRq� �t٫1���%�.�(c�)���U�P�A�&��*�7z�",\�rhErT�-B� '@ؿ5s�^o���-^V8����N��s1��|�,z���&�C��LN����s������X�-ɶl˶����̎�03333333sҤ)7m���4M���}{��4������뭷�����hxF�|����=v�o܅�K�`�����c�L\����`�}8�s7O��3fb���(��FmJ2VM���SFbͼ�x����gV��!cM�/
�1F�%7z�T(��c%Bg��$y2t���V"Ek�ݍ�e�S��X��m]�qh(�vF'���T�>+7f�Βt�>�^��~?��$�nEPC��\��|8�3���?oO �O�� �] |3��3�1?6	?|:�}��a~�r��v�/���.��_�ų�f��ɸwg
ݜ�'L������x��ߝ�Ǐ���O�᧟	��XO��Mϧ[��'k;~�c�0����� �O�+���R�@`��:���״�%���t�I������.��Bg\;�n�^�݅���t�O�:㫃v����]����j�Z����d���4�M�=��] F${�� ���Y:=���0�kgܺq׷�Ņ�8ܠ��d��Ơ'1C^�8$GV��+{.a٤�ػ��zW�Î�:�>o���7��ۧ/���xv� ��8�%-h�8����v�(p�cB�NX6q2���6���P_=T�����9E�����Bư�?�оܼ�c
@������9"M냪�T�O+Aǔ|���#�*�2�m�\�x��h�C�D�bk9R��($�У�6vE^d:5z*P���Ҥ4Te墹�-���߹+捝��;!R�d�(��m����jd�#��,V��y��Ý�X|/�e�cY��e?���1�	�}����D�Ȗ;��#�GF�1��2��xD��9��������?!�]�����V�`�WPX$C	�B��C���?&� A�e��E&o_��Q�K�m�tl�
}ztǰC�Rߌ��b�mjA�vСuT��#��#ǎ���c���C[��[�	��ah����pr�n�X�k�l��cgp��Y�������c�H�U������Y(O���9�pp�2��j1��_�.�r=G�Cu��H�j�D:��mUY��H���^�V5�j�,|��4^)�߰w
~v�{�2�
����x� ���#�sur���G�����9Ϭ��������[B�7�o�}�n��Iu��w�"W���۸�֛8��e���1e���V����n�%ON�cE�5zFk=���������c3�a��٘��}��#۳~�հqiO��Y�<+W�5O�<#/7�� ϭ� y"S?���B�7�o�'�ɫ�i�e��/BVuF�
Q�+hq�8�v�¾x��S!r��6���z���(5s��Ʀ]{���a��}�mC��s��0�t�Lb� �b
e:ľ�`�� ��B������uH*.ú���5:6qOI���6�B����]n�� o��߱����u�_�Қix7��Ұ�8l)5>���c�c0�����=!�c��?�PǢ�����yO<̐���y�����G��z=�u{�a���~������<�ܳP�i�%HJ.
#Q4�!����n�؍ O�MRr:c��x��G�������r�Y�������m����]g ��/b�[���g'�I�johrG����-�.�8�U�aH2i>n/A�I�K��:���7� o(A^_���/�ɫ�;䱻����+��;��1vbakJ�ƿ J�bh�T�m O�y�(H��A�7j�j��C]2� x,��c ͤ�2s	D�k!J�;a�0�V9�!�`D0�AH��)Ӭ=� s��\j�V�����bq�i�X���rxy���1q�G`�c �;c�c����5�1�)��{?v�:�<��/�Ĺ+�e�N,]��gN��#{��{�a����׶sF��	�1y@Ol�u�,^(D��\�R**�@]s;�f ŠG�����Џ�� �~V*t���uBo/'��aN������^�8;6�f���\���7�f����ZV����p]��h�7�;�׳=+ݟ�Z/�y�~����c�g�h:���	��#�����<���L���t��c^΀�����|��}�� k)~�|.�|4	O���ۣp��Dܻ=nN��n3�MÃ�s��5���m�������Mmw�Д]��l��?��s���Zp����bZN��MXA�&���@���:�G�������[�\[��fl:�(��M��@��S�Ow���b!���e��`^ޛ��W���������b1��#r�9:E..�w�#]g'���J{��q�qn?�1�<�p= 3D���6B�8n�=�0��+V��=�����xc�b\�>���Q~q��L��	���ux:u)~�9gbJ�Mc@+�ʝ���wAC~6*���� ww�ge�� >NNP�1��
a�$C�#c��y�X��9[�	
�ء�� �*�Z�`�]��7��- �.>(ttG��yZ�i4h�2�������;�*�F�^�l/�u�$�"F� AV���6#9Æ^d�O_xIm��H:��*GN��?�>��%���|�X���$�]D�#�R�R_ҿC���u8{KB<�xӄ���2�1�q_:���;>Ǘ!���{��CZX]_b� v��``��%�ݵyl��m�������78�@���^�\_��Op�M���Ƀ���T��zG�*�Y�(I*D]vM���goĸ ������=�r�"zWQ�����8�{7գ��ON�F�-g^��g�y>�g�����2��zw$ѳ=�l=�^�X�z�c��u�+k�@�$�g"3$)qH��GV`�]C���]b@��K*�૭'q��5>����P���=#�!�o��F��A������O����~x�m:�������=�;�u��h��]Pe��j��]����-���*�A��8à7�Q�*�Sa���8�"9&:��B��m8:})�_�I��Gr{dz��ǥ
�Nm� ��!Op��+��z&=��f��wȓ�\���j�AZs���=i�%(�B�x�%k!�N�6[���U��&��wDznD$��GH��8;?b�4Q��!
l�u�Hh�7BO,���q�y��B��&D�t<���7�\�l�5�I��6D�އ��=�w���w���wXq�&l:��s�aE��QE���=��X� X��xD���|-0����e��Wȳ�l��4������/ܵ�dN�f�SNA�Œwo�&\�{�j�`��X��6f��O=Ĵ���Ջ^�G7���!��/�c�[TYv�B�l�\x�Vgah�"�v���J�� ��������[���Ap|%��� wJ&�ʁ�GM� RG@d�k�ȅ�D�E��_��P�1�
N�9ܥrȔ�z�`M��u�X��1C��pHy�!�n���e�1�!� �&�7A^g!$��gA^�W<n	P��@ZUX=����+$i���!�	Y�`ؤ �I�0�<V�c!�[H �����O�,�/4!��h�jh��	k�e��PkS-���/���b�<�J	U2z��ӛ ��ЙX0f9��c���F�-���Ek1b�^�[�ӗ����k0p�\��#g-���+1c��X4�wo��'�ѣph�zL�c�tØ^�Ѯ���iT�D"�
�PzicB���,$��0"��R)z��"��`��N";tҸ���	�+Ᵽw&Ύ��[�S��\����
�ʢ,��8� /o/���K����
|����������������A��A���a�捡��!A�G�������3��	�~b�ZD05?=��_>�|E EЇOx�����\��l~�l1~�d�}4���'��[����$�N#��G7��[S���$<�=�}����~������{ҷ��O�����׻��+��������������q���$���ӛS���a��� �pa ~:���o�7������٦r<^[�Gk�_L�-�,��_���3#bpt`(��Á>Q��%
KZ�cL�/z�y�>ȀJr.�p�#���,;{����>/'×��T�8��E
!�Y(�]�Ċ H�T+k���Ȗ�P�uƔ�|��c?��=|:f>��g��GUT�.�/ĕ���قk������;�#���.6�0-aTi9�$B�������A�,����8�[u�>yl��B��	�
Lt�ٶ��@�������e�J�V�t>m�Ftt1�^�G*�[ �A�F�;�	�x@P���M:D9�	��9+�R�P�����$�''�,%���(MKA��<�6��D��& ��m��8	��\|���k�m���e �7E 0�Y �a����ۇG!"��M@�����^���b�c����~q�2���Ű�S���3aC[�,ֻ��r�y�A���-��K���|ʰ��(@��
��V<~�R��_4<]=�s�o�ع"+"={`d���o���-��l&�:��Ж���0��<�C;��Kl)�]��Bpp�:|������G������w��_��;p�ѧ8r�2�4wA��[�|i�a���:/�ӵ��)q�Ȉ�FaD:�֡[i���CJ!��2�>1��%
�P=�Ɇ�8��
L�����nA�����ḧ��gZ?|�=n�hQ��इ�ݜ��D`f�("��H�#���$v�ʵ0���	�\Cp��D���n�l�>y"�L�� ΖG�:z���$�2q�F_j�Lr0`'}�CQ�85k5��bB�`�#�Ju����V�<+���<�'-c7-���͐�@h@�7� o1��[��w��y��;����[Q�)��NBD����A��t�N��f'l�B9R�nik蚩>�J�{�H�;M�`�R�z!5�G�,x��
}�!طf�$�+1O\u��sF|̮Z�k��ZIk��`�Hjy�67 �� ��>@�7�l�ǘ��L]y�g�º�i�U�ǡY8�uTO����\Wj �L/�s����c��y���#�?��O������������M6f�;��OL��D����^����y���z6݋e���⓷q��cL[w>�_���y��B�Q�=3�ٔ_���
d%� %��*.���� T1c`��H�K/��`���ht�p3����A�Bl��B���	bkgZ���]iʖ@z��ٰK��C�U҃.>
Q��'`�{Zp�
�'�-?i�>H�V<���y�!�v�؞^]+U1D�z	2�<��Y1L�P���"�l����+*v�c^@�6�����K�'��$�/���x�Ix�#��ۼ�P��2g�9# �Q�Hz�'�*�`0f �����WC�G[p#tupj"�lk�Z:�r�wB`t)t�@�R���w���z����4�w�9X;j-6�d`U�"31��H�Y��o���+�{�D7}�LA�q�0t�r����oƤ��z�!\y�]��G����q�0�ww���FnZ⣩p�zMp��]m��3}����N�<�\��6D"�P�]�vp6aHzv���upce�[V���������J\���+��qyV
��M�;3��qs]nnh��m�x��#�>�?��_��¯���38M>w�~5׬of�o	�>��߾��?���?���?����F�'#�秓���	���p|�� <{w(i8�^������O��oO���F��C��� |��h��V�����cHC�w>��l�{�'p�p��8���_w���:ໝ����v�bs3������Ex{6�t\��s#qrX<NI��>	��-
ۻFbc�`l��MB��M���bqc5bYs���0.�CR��-���Zdy���U�(��W�/�\�Q��)�Z���8�c�۾K2*�(R"��+�yg-F��
I�)���EV�����l��g�q�-��^*�`>U6�.�,:�'��W�j\�H�N�ր*OwD8�!ШER0�Bu���:�г]36�^wT6!2[m,�J�.�#�6"�H�#��C�^ѵ7��+z��c����G���/�:�a�9����≩�q�N&��92-24:k�7�޼�߹�w/���.�����x��Y��:}��*��o� >z���(��ē O
g�� -�!aB?�0j101LY��Y��"�����I������U1t[lE�A�n��������"l�@K îg���?5�3����z�� ����c����I�5�9�z���sb�>{���`�ҏ�G��	�pN�fP�b��Ax��5�;r���z��7�{���;Op��������g٩+\�m�{�n\;s	ݢЖ ����v�|��.~�?�NmD�l�z����y�.]�đ���L��Z�	��A����ӱk�b̘3s����K����Gxr��]�2������Wq�ֻ�ttF���Ěz�5o�`�{dJ���X<��-� ���;>��f�:%܌ΐ�ʜ��e:����+�Ð�NB����yJe�9x�5��J���%5��>qк�� %��V
5�c=>�ç�ݱ����ѹ�0}������;�R܊	6�`cl�A����w$��an��r�k#�{�<	��e�=� oՉ� .;H�pVp�
�/�g��y��_�@@v������B�h+7��p)l2�C�0��	Х̀k�"�V��_��pow�����*�uW ��
I�UXWqȖ�t|�<Ag!��$��ŭ/�]���u�?�{7[H�?�#1R뉯a��0y뻘��
V�=���q#�����7+=���*�M�8=q&��K���,�W��d�����oq��1���#�Qn ��zy�:��:7���h��>w?UOǆ���f��Xv�<��7ރ�7!j|V�BR�!�*߆U�f�+�H@u��3�ʣ^@7>�(��h���c�8U��(�>f d^U��	����f�D �V:;X[ka#������~\��PzQ�a��s�-�M5�v�yX���`.���c���q��\�w�l3�MӨe1�y� vh"ȫ$�+4C�<� �h�.�����/_pת]�`k���9�Jh�C���侰N���P�Ā�.M�h���:{l��@�1��M�:o#�8� 󮅃O\�j�RG�WCH3����n�һQ�]�[?����A� ��NTZ�#�%Sz/ƶA+��/�!\�S�����1a�*��� =�D���ѡ�0t9	='.B�q+�g����6�ł�۰`���4��DmE)r2R���� !1��� �t���D���	v:jY�Ao��=	ɕh���n�1�֜�㳩ź�3í�5�x_W���=.ͫƩ�y835�^�\�����pmF�X��w��ཕ����w֔��-5�nk�v�~�ԋ��`���|������6��H�tg�xH �x����{#��mZ��ؽ����>���n��J!������Dg<$�|t�/�GG�����#��l�gG:��S����^f���t.����׻[��mux������<�7�oN�ŕ�8?4	�zG�p�h��=�"���K*=1��s11��r�0(�}���%R�j��U��_�zo��"���5ۡ]�#Z����F��EF�$�r� �V�Xk�:��W�C��ө���c3Nރ�`]��Ը!�ʜ�,�!��S=v�֑��⫠<�p��-��b�4+;XKQN��Ij�oB��=56.yGc��	����HS��
��Z���P��������Ym���qd�v�zQcO��(vrNb��nb����p9k����6��,z���o�³�qb�2� h};<o�g�͘\����YexҶ��1&䉬�-r@��b�ڄGwޤ������_~ ~�	�ʱ~��?}�~�w�\Gyn2�t?|���
!0���"��-@
�>�����]�y��Y��gޞ�����Ӆu�^�<���ҟ��.&���ō�Ű�O���y[����0g��?'g7A</�s��*>��%/�����^tZ紞�Q�>�%���F/�L�|���m7����Qo��"�0˖9�%!�Ϟ��_~�ko��k�|�ӗ�űKo`ٞX�i���D�@�9����M84=����_߈/|����`��i�t�<�>}�'��������/�ŷ���O��{�0f`���۳��\a��4|����޸��;T�?���Ԁ�14�\P)��Y����:B%��9�UK3&L����Gb��9r4���t��ƀ��л� �0�z�F�!Cp��y�Y�VR5�*'h����ݠ�^@^A�d*��z���"�>}� y�{�CB����\�GXy�箕��P��M��1�I\IƿC��j�-�7�́(mA�~!2�l���-�	��.��,*����?J���vCR�Ҫ]Wn��llK�AS���a[���c�pl-$���0�T�J�wV5�\HavN�u=�Ȼq��W`��lZ݆�c�%����w��v�`�����&����s�`M��琗#@�*����^X��S�N���Y~Y��y?��� y{�w�z�l�V�v{o���	����A��@�Fl�܀+��	��u�!���.�x{�<�������m�<"�����!�{�n�k/ OQz��K���䞇��O\p���CP�]�]�9��AU���1B6	���>����O�i�H�`�T	��9d��,c�+�BW��ڣ�ܳ���`���̝f�� z���@�u�y�Y�#�ٸ$�>��ɽ�Ji�@�5+�
e[��b+�&o8�sA���L3�IRh�䁰M���P�T������0��U�� mX� x:�Z�&�DydR|s���G(t�:DQ���. �����bli;���1#0	}:��y�0z�*���f,@�acѺk_t8
��LGױ�n�24]�V�f�y�DT����z��U���Z{�q��bAF�8h�k����=�	����F�4��#Z�B[�}Ԏ�v�B��XLj��CjpgYk!u�ۋ�qw[nmm�ז����l��3�q~l".�M�+��qi\�NNě3Sp}n
ޛ��[���dM6>�T����G�'�g:���<�^�n֕������T�t[�q��[�]�x���W���
�YQE�������7�U��9exwzޚ��7�(L���qit~98�?[Ȏ��k*�uJ¦vqX��9%���A>���nh	wD}������s@��>�y8#���Z;$����X'D�l�F���:a�V!�V	o)ܬ.d"��EQ��B��q�RĩeH֪i/C�Z�0�a2)B�Rd�����΁�Xڧ�:s'���s�qt��}� ����� Jl�cK�=<!u�G6��@d�Oz>��)���d��X�����D��\���tF���I��V⋚��*�GAj���p�
,;��ݞ���h��R�Þ��ᑪ�~`�QM)zG�t4�� �->�>?�~߼�>����/2+��T (	M�3�gh2��?
��?VHӖ#�!O�H��ԨY=vvP%x��xt�>���<|�����X�`���@��9��_�������D�ϟ��ݥ�����^�<�2��?�x�Gɦg���@�KP����;^��g����� �!�%X�Hy�Q��.���+�Ǒ����=}d�A��=��o㗟��~��/������g?���υAk�nB^\2�:�~߸�vq��4�c?=��o��F�~�ǡK�����ꁊ��h��]�vAEz�08항�qe�����)�W��w�#2sRP[]�ƺ&4��ʪ&������{�Es�N�O����Fܥ�����1����!��9,	�gᏀl�������A��^T8y{���j�.ضc����޽���?��'_�ɳ�q��c�xB�?z�[�>�w㭻����b؄Y�!W8P�M��5@%@�J�8&Vb
A�>�_��ʌ5�;h&�d�Emh��k�Q�W�ө^�_@�����q�Z�{'�"�*%ȫ"��z��C��^��e�E���J��uh��yY�n���QZ�3k�q�i?�� ���%Ց�}�jx��w�����7�Kz��7��u�ڽ}�Kh7�*�n��q����W�r�I��E�Wg���Da��/�aA�����9�C�s�{��?B�ϴ��_~­KǱ�wg��
~yǵ�B��'� �����*<���.:��u3�{�ql<p��_Ǯs0c�cxugȻE{�lͫ�(��9�H�y��^���
��-<i�	�<��D�y|�yt�i�kBY���m+��+a�M7d$�!� q� ��@W���a[w�Z:�֪�8���;)A$[�DI[!J��\d�1�p��4�kɣyϺ�A��%w��{<Ԟip�j�S� 8�{6�?�y��!Pf��&m��σ�� H�3*���~P'��6�;d�%�x���;G�c`	�����A�QJǭBjTW4�4�ħ ���0fm@��˜���+�k�bfRLv�Ă�j>��o°)K0e�b̚�c��F�A#�o������B�����:��!��"�K�BOb��������>NZ:�!Xk�H��t:�:;���^g+�	
�r$�uP:��R�bWw��Q��9m�qjdNJÑ�q�8-W�ⵅT@��ũ�I82(
���G�"q�_(���鑱|	�06������\�fd�޼�]P��K	Җ�HV���
a���y�w-o�H��		�8*���D�H��Hp�-���]ֵ/����cY�?��bj�&d9bt�c�\08A�^�
t��Eg���z���Q�D��J<4��Ko'F���v��U�� ��_HC���o['e�pf���d�pQ�n���f�:�arrbe4T0SA������VbW�
�l$R)KB�J��!��R��瓣ӣ���k��|��p篝Ù�{���#�H�����<Z<��v���H�Z�g������a�H&d�H����� y?'��I��7����/ҥt�JF��"��hgo''a��+����Zp/9�z�s?,_�xru7�H-ao�@�� ^�!�!x��	ߖ���������o���3�ud�x��O��?}�#����\�g`2�{F���E�o�$����1�}W�o����cx���sP�_��������F����-��q�#���3Z8�3
	�y����<�1�1Ա;6!)MXn6vϲx>;�Y��¼�^�<���Y���r�;���y��~x&o\a��ǳ�Ra+C�j-�������t�=����I31q������:�usW�T4������((,��ވPwl���A�w$*=B�j�l�m�R�ж�5�Gnp1=S�蝄��l���9�ms
Q���&`]�	ȱ�G%5r��E����t�F'Oz��B7������/X(�7�!:�Mŉ�&|�P�'�����;�Y�S��QE���w���3%Ԉr�߸�����Dck'dI1r<v�>��c�����;	�إ?���@C�>�n�u�z���#M��S�����+!��C��t�։ ω�B��B�B������[�f����3ђԀb�"TF�F�o���	�:�p�2��� o���7�ݵEa]y
ʚsPV�����ߤ�:e�IAr��W6�|��jAZ�����4���꣰�:q�H*wAZa�M��J������~���B�c���H�^����5_�����B,s�@�1b�W��t� �,�ʐ�6&.���ӎac�|S��y�}���='�C�;3� �o��%� ��~��������y�^=��=;��E�]N�8��g^���)��p#��m�+�bY�,�x
��Ċ�����#L����B��C������b��ٔZD]J[J��^���(��$
�e�o�`����?O�i�)!����L�)�JNAV|�5����l�OCZ��}�^����u��.��9�1�g�u�?�(=� T�a﹤� ]N/�TX����i ����<y6D�4�����y4tv�,�$!u��x^��z�	��rO! ��]RO�f�&g�!O u����S�8��O�s�X�
G�:�<��&±h<�	 5l�k���@��1eA��!��k`R+7�܀��.h	oF�{.�]㐠�Ek�7fk#��!ۍ	ؖ���+0�����b�ĕ0uf�\�Y�c��U�0cz��IT������#��$6@r]w$� $6�
�H�x#�7�n��RsC�7U��.�	tE��9���C�@O�@?O_[INf���5J�Tk���<z��Lh���5I�W�����&'�����8���b��kvw
�����쇕^�ڄaIK�4�	Y/f�cFU �������1�̬)�q�A��х~U�!����ީn��)�U�Ⴆ G�x`B���<P�f�5rm���#Jg�pG�i>�^� ��
xkl�°���� E	wU�*1ְ#��(Ͳ#��Pů���F��UQ\�!h#@&�qS����j�5v���R��cb9�{!��WG���蹸Sow��֐[� #����,�VMr��!�Iv
���K����svC����Z����'�˧p��	���\8s��1�K���Z�"�S!�J�4�-���r7����2->u���nc�@4}�K���=>��)�8��6�^1UrevZd�eX5�/.nو��:T���kC#U~zhmdp�Ia+����X-����UCf+��@V-�<�*G�Vm�ޑ�x��5�;t�]{�^}���ݐ�j�/����5<�p�/*������(c��Xw�-=g=ڔaPǮܹu����߅��;�k���#��D=�TWW4���U�p4	LB��DTx����B�Ūf�?�� �E�������bic�og�o�@eq�򲜼"$�d�2t�>�{�>����y��"K����.[�2�Yb�1�Yܵ�/Ü�X|L�7����� y�>y��%ω�ej(�2���~G����]�.X��cg":>�F�H�.��H��d�rES$z�ţ-��?�r183m���D����t�m�[�FQ�.�}�0 6��G�K(j=#���$��(�f��������={"?1��_D��� ���2��΄�ZtwpE/'/�q	F7�/�{����\�>J88k�t����www��yx��=���	�J'8�)UN�+V�1���kK�DR�}PTބ���i��sp]h�^*��!V�!�J"�b�քCv��O��SqE�(߈9#�ܕ!�3U1mȳ1�1C[�x��A��{y֮]_����	����FC̐�	�J���u�q���
	Ȓ�A�8�TI3I�)�I�Ӡ̘	e�l��̃,mYs��]��Ф��m���W@����YD�.�<w	lr�A��69��,�(�v��a[�uG�o<���0�8�����`�M�E�0E�' j���i�U��z#W_ńE�a�l,��B
�q@Nz�b;�''�"��3gƌ~��y$<����ϸ�`�{����+�ݛ����ª��5�(�� ������0n�x�x� ������F�H�
��r4��W	�hZD�ƣ`�NE�����ʉz+�.	9��e�M�D�o#Yd����;>�>�K�(h]i!�a�QHJ�BZvV�v�K����� �e�7�^}~.i&�|���5�I#�A���V�yd�C��EC��[� y��d^���	��
�ñx� ܉�D�}�~{�Pd�&}�����i��켲� ˆ�r�E7BOǖzW@Ԁ��.%-h�8�(0J��Pl�1b=�}im1#���հ��L���-��1w�B,^�3�-�ԅ+0}��=ŭ!��?b*� 2�a�%�N�:F*}=�0v�B����HtB��E��(%Ыtӣ����buD,�R��H �E}#���ڹ����TP�z����݃\12����hk��+ڲ:o�*6bAٰd-��٣}�=�ct��CM�J|lQ�F���i�<Gx^(�
�4GR�H3h��!�A�h)"�6�$H! ��+`��ִ :� �|�U��Q�%*��:R!�G9M���Q��ɁC�ֶP��`G���tL;'=�l"9��%�y��)�s�r���}rN{*H�z��\��QW��� m��ch�(e0�R@d�u������$`�^�X�d�o���	���Y�ڣ¨E�\,�(ջ ��y�:o�?��'�����x��W��k�Ѿ��s�t�Yb�$8��q�$24�~I�xf��Tx����B0RdK�g%��@���X����}:/��Ѣ��u.n(��`PA.��V"��#�hB~`J"��F ���X-�`#�I*�w͝*�l��sڱ#Fw���a��8�u7>��=|����q�2>��>�9x�u*@޷T��������6�S��ş�yXg�":N�H	#=� g=�U�Q���;tĐ����ͬ�}��w����:�A�R�~�qXU��	8����3��X]D�	`�q�����O������eY�aP�X���xÙ�bǮZ��Y���e����"��x����@�?ݵw<J����r���=��۱,���Z,yz��ⱼ�|���7�#��ι8�TG`���8w�
�/]��3cۦ�3j
�����Hc B	|�ݑ�СT��.�hk�Co?���F��m<����݂��=��}|���5#��\���6�4�;J��QK��B� ��#��/" �Z<w���ڂlt����>|����D��;��A��"w?��D���ʵ ���l*��\����n>.�QY���
//vc{��y4,�=ᑶ\>����*!$�����\�l%�	��G�s�.�Tj;�<��Ȓ����'�\�7�8�b�� @ޕ�0g�|�D�"۷ Aut�!�k^0�I�x������<��X�BgC��VB���C��8~Dj�ǟ�4��Eu�:��f9�w�|��e�
�t��Ѷ�:*��iJ����}vk��=D>�	2;>�{���< �¾�a6�ȉ�s�)YU�q�b�V�3-�;m�­�Et��*�n���+�`���8� �g�Ɲ�"|៎�	�����h��`�;�>�<|��y���y�t��P��:b��'N��1�h���� ��m������=���!��|�!Fm�c�5?��zQ�=X5^�U�5H��%��^�m��BZ3u�W��C�Y�v���W���2�:���Hئ�0�DȊ���ж�-�B�rr"ey�h�]�C��p����_�s�kP���í�E��{�.Bߚ-砬8k�!�� ��<i�H�V��]�_ ﹻ���v)������C��<�7%C�C � ���Psx���B�������k6�� E� h��AU<��q�j	Q\?��Bӝ^�!��ڔ�O>���^��8ƴ����W#9�+�tsL�`mF��P�*?���Z�}�P��qX8`&�Y�Q�cƘyX6s	zk1k��^��E���^�9�=�^��e�����G<�xh���K��pA^�+R����W� ���:�ڕA�Z�L�)�^���aN�h#�����H5��~XUh�P��E���Z��鄎���oD���Y�e�<�	:k�ډ����F[�T"��*kA�j)9\�f���aPH�$��e2�
�	���%��^*�� F�	�E�p�%�R(�[�B�oΪ"��*l�D[[%��[H��	����a���.E-��]''rWнP�)l���q�Rl�������� ��Y'�D0�i?v*(�2�'fP�y-�a!�(R/x�܅���588�:{8Hi}�E�Z�&A���D�� ;@Ŀ��D�X�(�\�OW Q�H�G��<\ڻo\<��4=sp�_�����ǔ�#�"�JF�g�d�0�%:��EӾki?�l4x`k�u�#΅��k4F�KG��;=��L,yG]���5&�����Ҁ��P:���,���:�(4H��#Q��
T���<dR,�����p��;�u�%�Fbb�!X=n:N���G,�ݦ����k�C�h��RB}E�W���#w����?B�]X*Vۻ���Ǉ䦐SūE��\���û����0�[�nW�}	����-M�F�h�ߎ�*��-��-����၈L x"p��������^<��'YF�Z �����/g�c8c�c7./��|,�a��eKo��y^�"^fq�2�1�q�V�n[m�aW,�<ad.mg�<����Z]�✷<�֍~sN*%��7��j47�^������AzL:"�lKл����zGs��;WA��> �zl�kC�V��vt�V�~���d
B��?J�����-,��Q��~OΞ(��L�����&#��X���\��!.6����Q����W�3�<|�Jەд��/��0��5� /�3��(IuD��¨��]�]��[Gj����������t���v���Дԥ[7�5V��U5��+Q^[���bW!)#	�����	��P~���Q�"��$�ʸ��G��䝈.��E�1� //� 9T�d�U�߭bC��<�k��y�^}͐2���yT��ܶ����w�h�������%�g�D2#��&�T�ÏD��Bi���e�>4�ux*���1�&rx���f^��$��	lh�� R_N�9 �ҭU���������^��m�5���6�/���.b�#ؑ�O����o��M!X����o�o��/�}Y]��/��ؤ1>����@�W�G�w���cXZ;{�Ŧ}�c��p�!Flz��yMw	���}�][~⢃�)�B0�����S���乐$΄��Q'N�(bD�� �N�3�4���K3C�5�>O�(a�3f@U� ��Up�_�ҕЖl�:3i�eK�R�Ε��Up�� S�v8�o�M��{H��cГe�!O�x��y�B�n�2�7�i��N��)� ��0��^���J{��m�O�<��!P�����}���@W=�����]M�8W̓k�th3��ʿ� ��B�|������T�-���֐zUA�Y�؈�(GW5U��L�b�Ȉ-6�X!w�J} vG�c�G���cΰ)�0n>&NX�Y�`��5X�l=�O��!�����i7��=�]�����VG�ܨU�F�����0J�ݵ<�1���~j����ir@�J"��̢�t�-�+Ѝ*��J%Jhy��`�3��{P+��^�δ��^���vB	��K�6!��	tC�V� ��r+8I	^������S���:��u$G{8:����V{���b�#�d�s�������	P�j�R�J,�V-���DF?~�:�
��yj%6���s�����ɡ�( ���!P-��Z��N����
^�>.�e5t9�$�K����mU�r�*�uP��C�u���A I)��e#�Q����/8�������b��̝
~�sWLʭ���9�|�H��	��<��!��%��}R2qp�2�.�9�C�6����x��|��!�͘&@^ݳ$�� O�$��
-"il�;F�S�'�)���7��y:��w�z+�|��b=���U�������4��ީr�u�ȢgT�nB��R5�H����=A��*�zD�zX!6��C����&Ua�)w�cd>�����J|蜀/�p��'� /��G�)U��|����<B�Fhv�e`~A%d�:�]�0�cg��ֺ���t��$v���Ԏ ��4�B�P5aKIV4w\�"�5�=! Q\T^� �gYҒ�O��P��d�;��m/�]IH�@l\*��9
�A�x[�[�x�:�<^Ɵ�{��7���c���X59�e�uW�
�8�ze�+C?%-K����Z�%�eW-�Ð����
�
����Rw"9���r�31v��Z�������[1z�Ddf�!�`-�����|\X�D'b^Jf�aezf�b�1 c��1�?
�齘����ͤ�ʸ,L��̘T�
K�ڌ,J��ZgPp*��uuA�?A��#���71az��cGb���jl��Ʉ��p�P�F��k)��E!�f���&4����:/T;z!�� �c�T�x{���j��WWlٶ���?�w|�n?��[p��G�}�>ޣ�����{�Ǉ�o���wp���db*#�pѻ
�P���_�/C^<��Ů�8�����#spi�VL� �Ԁ�,Afh|M�y-�����1䱻V��,�'@��� ϳ�<9�1C^�V�+��.�i�(�v��Q\Q���Y�Tm�Ԗ�
jdJ���� �;B�$��B�6d�>��=_�/�G���2�d6�� UA��#�!B��C��" Ws��(�g�`�e��M�Y�kf5]���%��36�����a��Wpl�9+�O���ْ�I�1XC��izG��w����c�?��;WNa{�v���-t#�;x���+��ᶃn%W����8����Ŷa�q�{Xu�>V���3ހ��m��=&1�݀��&Q�	��F��"�%PR�Cd_
����4/K�C�,#
Wм����$i���I<�U�I�yfS�}�1�t]:�.=�д�D�q�uYzZ_GSg�:�>9��Wo��]d#�;y�>H#VA�=b�H� ћ!O����VJ;�<ώ�}��6�?lSzB�VI����&(���
��!�l����<���0UM�6�@6�+lsF��r�O�3򂹰ɟ����˟��Y�(��_=]K&�J�RC Yǀ*8E4�EU����Q�s>�i�0P��"f���Jb�
�k������i�V��æRA7CGM��	�r�v�_�#&/ ���c�tԶ��.(����&D&���'n�a��W/�P%��� �|�䀪8#r���k��E���_+��E>C*E��
�VyV�g���F7;-FSE>��]�J�H �bB������B�L7�v6y�2�me�ts�ɓ
9W������(X��V-�0e��R%�L&�L" �������N��q?DY�9�%#I`M�d)U23l�X4����0����Nv�+$B����i�����	N8���x��}�! c�[U
*Pi]���qv��(e�X,���rvvF``����aRO����& ���	6J����]�j:wg�5��b��=�����H�s��u�������5�8��n�9ݷ�����`��E�����2�J�=9�e*�@�����j=q����\����0`#�Z�UTq<#��#1'�=��8Ew$((�pA=3�8Q�fD%�k��/r���j��b@���R$8�Q�`��QY��ۂcɥ��,�3�=}���AQx7��Rkq7��%��i@
�	Jķq��+�QE��k0�sŗ:o<Q��15|��J� }���#����2�0�{w���{��1�C�����Eώ�3�'���Dz.>%:WԢA![F���Q��!�Ad8�s@cl��͂sPc�F������� �g��?''e")1CX/1!]����������`�t1|:fd���ql�3�^_���a�?'�� ,E�w����	�"���""�B9I�`Y

BTT���i�⅀�a�>��	���Ѷq/�bd�B���!��e�3xy#�΃��q�58���WFg'��������9�1b�l�w�ܕ�(l����Ri�e�9�����i~�:�9Tu��T~U���2�,� �������xF��*�*zO��ß�z���փ�s�	�e������	p������	sf�A��	d3�����v���$X(�ݼ�jD&���NX��+��^���ń"\N-ƫ	�8�^�!>��Wk��{RHe3�s��.��=�΢���
[PP�ZPvN�������֣���:�G�~�p���y�rN��
�Z5��*�<1��\�ER�x���w~�ƀ��8>w��]�֙M�wM���:c5A^�!ri���q�x��[��V��f����� ����ٰ��k�Z�� oE{`F (�X�Fu�Db�8����dk�����de�,����OD�R�Ğ�:��ΰQa-s�L�Fyw(l<a#��T�k�m�M��!���� �$��LE#�����v�,k䵧 m��ro�׮��}��5�p���K+^ù�qxT���p�3;�8b�j�˓g ߱��7B<�gF=��G����߅8y<�vG�����mRͿ@�n'�����䭨��]#����ʳ����C��w�=8����ޅ��ؤ$��%.���MĜLJ��],�q-7�<�m)���5�-�*��@��{.�� }�����a���� ��^ z�"z�N5�� ��?
Q6����@�
"���<���_�<��!�`�A� �ʯ-A�@�&� O�S
��:8�7@�S	���	�8|
�>���G�X���&m�r��6w<��*�AQ>NM��ִ	�V�X����HH�G����.AUp��6��a�`B-#�j�x�F �S�k)z�%��]$��1� o�Ԉ�Jo�ևcoD)f�dbPd��O�7}��ǨQ30k�*̘��f,Ť�1d�R4u���.Ȯh���j�g��/�Tq:�Q���T�z�lrB��9AZ;
V�P��J�J���"B�@�L�l[9�r.�I�O���>�^+���D�YO'T��B�I�#A���R����K��
<'g-����x{���/�s58	�2�dt|�10��ͪ�u�RfcC�F����%ȓJ��eG0F��8�(/��@|b� yv�*3 ��`��o|>l�cpS�� r�p����������&�6�7�Z- �?!���V��i0�u]��Ο===��d96���%28�9��v�4�m}]�C�	t.C�*�������p��u\}�vo\�c�w`��-8�{7>�uk�M�?�!/�Z.�lӥradm�{=M�ع�S;�}�����&�C}WdŐ��S�?��q�ணZ�"�ت�|Qm�@�m9l����Ȥ��s�t�eb�:i�Gע��1�]�2�s_�܆ks��m;�ڱ8�j^_�X���X���k�c�θ���	����)� /�;��ڈ�2{|���g�)�ᗁkQ�X��Zg:�&b|�vx�.�Nѳ3�����ڣO�&�ڕ���Z{�k�����;��#0{yT��0�3T�A��?<@��CC���o�)Coc<��S˾����!�S^��c����f�3������v��wx��!�ݳ<2����!/!��;�G�
&�"�$�3f1�ZH�F�h���H���
��B�ˀǖ<v�2��� σ`�c�ܽa��`j{g�=����]:��X�f-ƍ����pټk2�K���|�#�T*nW�ý�:\O�ē�j �&�ׇ ^1Bȝ?���1����g��H�/�i�5�Q9{=��Z㵊�؞\�>�$z�y��"��	��Ѿ�5���-,BE}=�w�РPx;�x}1kE�hf
�����3������\|�P�����(63>Ȕi�Lp0����]�<�W.����WA,���:���D9"N4@�9�����V(S|�9u����Rj�j�P,����1�q�!o���S���G��pt���=3[��/�|��k�C^'X�yV�������]x�'�@�7�B%|A�z�9�I�v�KwA^�6�s�* 5fC�Q@��J��6��$6%@�%�c!R�S�N�DP]N`�S� ����<�L�H2}V�r��>޼[���1��9�:�� ���W3��P+m^���Y�^���{���C�pf�e�(�������yS,vS�s��k��/�L���Q��^�<����~�U�x!�P�Ձ /ۈh�8w�c*�>u,ywS+q�f\Zp+[-��q��[q�.6����+n��7A^�-���"�ԽI���=�ɇB�L��ʑ@N�G)� M���2M��.k;/��&X�<!QZ�.��ʕ�ۅ������
���t�d
6��饦ح����*;Q�9aP�?-y�yV���r��7�g�WI�_�*(B�@��_M������(U|��	��&B�3�yP��_C��piZ	��eP�N�8q�����/ O�_�w��st��ʿ5"Bڡ�W9z���>�$��"2`��k�~X���ɭ0+�����X̜���N�ؑS0s�,X�3��x��!3V���h�VtAl~BR��E�H�$�L��ܠst6[��]�튤@g�Pe�E���y����Z
#��781�5�,�r�D�𣂅]�MV2��1\�F�R�u�k%�#�f�B��uLJ9L*5j�i��[�c�_o�<�B?6��G�V�F#@��,���T�tnf�3[��0�+d�=�`	��u�تF����ԩ` R&�-�b�y=>�ˠ� g;[�X��˒�\��%��o��1�q���(X�_�5�E��;A�-��kHVKQ��$�W�ܪ��:��wn��Gwq��M���E�/�!����`��Bt�%c�����+�e�J�8�>��O�	��`������ܒg'�X��C^���������Rw���L�G���ct�)	�er$��p��Hg'��}�>���:�hi��k7a��X8o6m܁�wa��c������������[����x/����[��r/O�>�Hi��r=��	�^��	\5(T��FKU���e@���ۮC:���.�Kޠ��пk3F��*P�bBOS8ֶ����np�;�� �c�1�ED�/�j����5,,BHƩ��x��%�
[�,�4��Y\�<������e�>,߱�\h8��KGDP�D�M F@g�ޱ厡��N�ǟ�-�w�'ȳ�?����$�5Y�����Y<�� �]�/C��w��I���8y"��׀�8�ب�K�?�θ�L�#x�0e*z��޽���];$���cB��	Er{t�8c�G0��8�5P����`�-�����1��ޗMI��+?���!L��1yX��B/:~ogo�2��!e�>���ޮz�'�bh��گ�w�.];���!~�4��F㩌-����n�h�����#?���O�|��:jYi�:M�z��@�np����ҫWp�ҫ�}�Ҿ��چ�hۮ��ö��5ʫ�_R���BL�6�w}��2���H�`��8a��򍻣p��Y:W���A�������ԵX:r9&��F�G&|9�5VS�ږ஛ yR�c=�B�҅ ��<!w-A��i0�����f������ �`+��v�&��[��_U!գ�ˠ�Z]�F��6©n� u�*�j7@_�v%+��co�(��B�8	�(�?�xR/lD��!�>Ф�]�0��G@�9��P��}�
�»d\���>e>��+!��Q�a�8Xs�5�t~�_��e�a�ᇘv�C�N�=��y��iT���pMg<�� Ȼ:i�+����ؒ���!T��낝��&��̐�%v����*�ƚ�%�?���� �O��Ɠ�0z�=���֤�[�i�!l�ށ(u�/=D+�k�$��Q4%�f�|i��$2�:/w�d��K���Y^fY{��Hr5˚Z&���Z)$k6���<�g��}�:������y�`Ȗ>yֆ���4���4��xe�EO�[	���pH�' �Oq�y�Z�B�2��q��M��f!TM� ��i�,X�M�M�h*f��8����K�V[�B���)��l9l�&�����2�����ѯ
��	��zb�s��`���Qؙ�3b�1�=�Z��ɋ��D�9s�Nǚu�p����Cf�Fm�)H����zx���-$�10��	i��?���'���}MH	4"�K�o2	b�u���eT�;�	֌NzQ$���*U"�J	o����$(�`���6hE�A�9l��]�4Չ%B�q�n�B�sH���1���� G�^p�r@P�p1(11�Y��y��e�ck�����<9�ٚF�Ik�g ���2!���%�A,v�K��w/���ek��,�c���߬x,��r�z<�P˝����F�+�eK@L�G��T{��/�E����8�o�~|o��&^�u\��-�,Ga��՘4n,�n� X��`��d��D<��ϓ�t�j�1*�?�x�H/@�T)��XJ�|��#��'��8a
A'#����BsC��ê8�gRM>(�MB��JT��!'*�����ak��Q��<�|�rq�=w��R�݋i�o,X�wVm�������x��ެ�'~����/�x������W:�j�L��E:+�@/�F�G;tn(���ѷC[��czt����1�c�vl�~]Z0vpO��@/w?���.�YE�a����*m�1`����DGG
S�$�t1����5?6�*�%&��.E�g7,ϖ:=^���e	.P=�6iw�!
B`H A_0�"霢�<��� su��X���X��bx4C*_OXxM�R�w���E` ��cQ����-�d�`��?!�e�ܴ�!/��%� �!g�u�C����=j��`��~���ʯDqY]�u�	GS��T�����H���dZ)�Lu�&��[�_����/_y��|���>��ǗT9�@���,|�X�A6:j�Z!Æ���wE�_8�`
�E݇M�=d���*��{��&���A$��uuG��;����g�ǃ��ᗎ����\�o]	6i�ǀ,���Q�io�ْǐ�<���vl��Ͽ��'�����q��S\y�:�S����g�y�������?�?�
���@UM�dj(��B�D��[��`!T��?�J���xGl8����SVb��ŘM���+��3J�J�\�C����<�/ O�=
"�	/ φ!��N\�����큼b��{aS{����p���0�v�u�p�A����z\����0��	�>@���v�
��o���p�L۴>%�C14�k�!x�= �6{�ֲ�M;I���z� c+�o>C�h+�CSq��U�b�I[�e�[t�70t���p�3�V��S���d�0|S+@��x��y�ȿ �v�_ ���q�<]{�
��!�e�<��[A^>u^�M�8ypu�!�jZ����b�{Xq�>��}��;û���M�z��� mx���p�C�D̩�y{��t���zw�H_�]DZ)ά-�υUT�g-W(J��̹��G�0tIS Rx�s��D���Hk�&�,U$��A�n4�Ow(r�BƑ��������%�@���j:�sw���V��a����P�)�*�f�[ǐ'	m!��y�@!.�=�6�m�rL��tzq�'@ٸ��Et�ªa�53`]B-��Q��'����,�*�|����޿ N!0D4�!���հhDBDkt�)FM�؅`��	��<�Tl�r�X�����nH�i3f�[��S�c��)X6w��،�[�b��Y�9~!Z^��6�]�E =�$���Ra�O7�;�
�w��<���$B�1j�ɱ�|]�arC��:��ưǱ�<	�|i>J$F�D��Vq�J�آW%��`�-&�l���s@b�b���Z
��n^p�sD���Iyq�y6Ag�0𱕋�aH!��k�����m�.��<v�r�{{��e���܊d��	�;v����yY�[��YF��� Yl�c�cp�X
-bP�e|}|�|nN�,�]�1��Kkk�WWD�ufh��G��qN��P��+���s����x������k8y�0Ν<��v`��u�0f4�<��/_B�I�e���)��#�-�wO�O�p��a"� ��5�j��08�%�c7U`yJ[��!Jo�W'�:c{�A�фt���=��]u-��2��@��Aa�M4�B�?|�>r�d\��ד��f�����YI_ܜ�_]��/v����|������/�M��������Y��Ò��3 �Kђ\�X�$�l����]1�sG��ܖ �	��4`Hg�}����ZaX��XU�nT`�s����NXP��*l���D0VHA�yH���rI�+4>.Q�2�1�񔗅���/��)T�7���ֱ@��������be��]@0X �eሎ�Bl<mO(vղ%���şY<o�M�1###���3!2�·��P�p���,��g*�H�oG�cf,,����85O��<�_�2x#��3l+�<�mao4
�7oޏŋ�c���� ���v�c�N��t���	�:�r�5�}���)�b��kt����'1Y�9�ߤV���z��ь���eh����2�����
�L/B�{���P���`�{Ç�IAA����Jb����!���U�hg@l@$��5��f9ѻ�R�?C��5H8��#� |��OB21���|[���C����;l�4p�￬�-=P���M=QߪZ5wCs�^��c0i��.���m���-n��d�9yBi���l���;PY%�mf���=g�8*w�ɤB����Nƴ����C�{�`ɳq� X��.�!�0g��u��ڵ;M��/��@�~8���@2��9%��$gDy[`��������Au%�_��*����4d�� ��hΊQu��ٓ��� ��jyV�ށu� �H����ڽIC�Rs⦫�6rD�KP��y�1�ÐT���8�U)�e�Y��{!*1M�.?	{
�.CR��nA��.�}���c�ѧ�~���g�����/,yyM�8g��jzo_�0����y<���k�p�w���� �5�_ o./�+�kw�9�M��cչ��~�&�| �~t����݆U�{���
�����i�o�4c%���)�}�68��"k9}���M_U�|ئ̅m��Ҥ/��剳��c�R�s�@�2��I��L�$qlR�A�6A�,m�)��@7ꨑ��"(��KB������Pd0C��̗ �+A^��3�)������}x=�ՐG�Z0�q�2��~PDw���	i�xX�π�� �� �i5D�VBNmK�'�F�H�_<V)# ���7j�\��<�K	��̐�U��Zć�B;�<��Co� ��q�+3�-��c�1	{:M�јh���j��?S��䉓�b�,lܸ+֯B�acѪ�XT����.�^����a�)DXb�b3���G-F����w6"�I�Pg�MNznzH��BS��N"��
���x��XI�"Q��
�\���')��^$�x��5�TI�@뿠�F�@�¨�rVkB�����8½�Z�<��A� ���-�����f$K���d��~yj[��8����wO��������e�,���x����q/C���,�3Ȳ,n�"0����f��X *�	�_[��Z�O[��]˖L+ڿ^!C��]���A��q�¯�J��)#p��>\x�<.�u�o����z�Ϟ��SGqh�&ھ��!����p��%/^L�gm#��e6�q�J�1{|l�;yO��|� oA_(Ua�J�;T�=#�:�䃶"j\<QAm��3Z�d!-,�j�:8"��^:G�L^B�h_�;£�����#c�AP������P�w�ķni��-�Y��.��g���h~>�O�j?<���C�+)���J�_���1 +��,Z��#&�Af�T7w����x����1�M-4ՠg]z4T�Ws�7�cT���؊_a���]�GbӐ)�w�-��y!�Q�!�/w-O�����Τ���a�;��1��<Oy=^����y}^G�@ h�<���>sV�P��l�D��OP$'��q<�:�j�����ak"%g<�!*C^p�Z� wz<5�F6���/����ˣ� ��{�,����F�䱻��+ ~B(WD����$t+�����C���C�a��M�4b�L��A={"�ۄ@/O��B�ܺ��qf���cG^+�6l�Tv�;Um��0�1q.u���G���q����?�N��NC0#��m؇�f#�ل<7?�'� $��-_wj���������l0R9���oDp$�	�jKkpl�Q��+�Lg<N.�o������nAx��O��p?0S=�����m��a
�n��Rl�1�a�}�HVT*i^i�v�2k-�u�,Y�r�Vq�w�5�9�2�[�<RS9�Me�n��#V�/s���왴�:���h\�,����7R�<��)E΅u�b���m O���ܝ����[���T�����.Y��8�M�E(Z^���+��\�u�y�[k�A�p
6M��o�WJ��a�D��IʏATz���q8���dUz��՗`]s� �@�3~տi�[P�z��a�0rӧX}�3L;H���6��<�cY��ix%���E����i�0�v�%ț�L����_iC�ݫ���O�� ��y>�����q/������;��~>v�:��{�`����q�.&l����!��6ĵ��M�H�lS�*�u�BVqZH/"���1�QT����8l�~Y�c�ge�RW��!
WӃ���}�	�����j=��]�); y���)*�����]�~��E�\��|~	���w�:u/���a�����~	�	�J�Gȳ	��}D���UB��Y ����p�
yBw�~'&��7od�+	��C�f7�"�m\	eo�L�+	��C�1
��(������b8�VCC�%����W#&�-n��io��~r��`��	K�ܰ���}fa�EX�S��n��T��g���)�0q�0L�:�V,Ĉ�3Ц�����!��8d��آH-jFbJ�CA�IJ�B�����
1���,�R*�K����?A�r�#�A�/ACB��Je�9A.@_�H�BR*�:�u2(���n�8p~�p��?�7@����D�:\3�1��YvaZ�0�S���e���1�qxv�2�1����]kO-kw>�u��������z���Pg�g��ˀǲ �e4���j�˸_�Eܗ����e1������v����V<�?z�"�0�B�X��XL*	<�b���cP��رg#��;�W߼��7��K�q��\>r 'wlšMq��A=�W/^Ʊ]{ap��	yk�9rl<~��UN:d�v��@��C��u�@_�T��,��Bz�+���C�H\5$�bX	�G�b�B	]C��Jb�L���jt����]��="��8c���H�ErD"i���p}1�
�S�,8��.ŧw>�'�_é�.xlJ�oAx(v�]kg|$q�'"=~;�{�XLq��k��a�̹)��թѵ4=Z�cm&:�g�[e>:��]I.�T��Cez�4�6;�N��5zcڈ�1a:U��B�ɮڠ� Ãx ��.x[�� h��>[���c��X�#�b9���׍�}��e��ej�	�&h��<j5:�b�_^ƮP:=>W�zFSK<�<�U�-y��tt���v�/��"?��ܵ-��-~<"��כ>�;�Y�o ��ܵ���������zga��3�s�
{���H4{��
5����]?��$;D���T�Il�����c�����)s����k����%8�b�ؽ��߄�w1���w~yxV�B�N8��8�ߊh�;���l.)A�� �7q��F�zM�����x_/�H��PZ��N�Mn���At�'���=w�ax��'����	z7$�l����&x4��mp%Xl� Q�1x�3��A�!C0h��'���9)��.^�H�NBqM�|�w�3^p��/�;!��R&E�\�.!د�F����e�k���%����y���k[�<;�y�Pa��VC�C�8�'C���MPP�����c晗s����/Q�%�_�:���a�J�¶p�� �ILH���Ӧ�O�u�"ap����My�Waͩ̈[8�[��g�=�@^z6��aSt��k�T�I�kt\C�Ʒ �x���3������}���`��[83�$�g��Fn���e�$��z�=�\�����O�s��3�63C�O?��W9�J'l��vgl���WȻK pi�.����]#Nb�:�a��{���&|��O�w���$y%g��)J/�Ҽ0؁Ö2�-<E�M�ri�[ɧy΄�	�y]�u�9�!����$u'��U�Qzx�2�@Ӵ��7Qv��g�����B�w��6��sA�s ���}�� X�ܵ�!O�l�<��_�'�%ȳa�˄�����&��*�=�]9l������TqH+��g�?��qp,	Qx��Ym�!-���t�6@�r�Z{`�H�K�i^
q�4j5��R�1����!OHkRa�<�"��j�S�&�$�fK�&l��C��P�5�.k��ĎA˰�'cmC�.��LĔ�ѱG���3fO��uk1f�r�������hN��qJ�{#��F����B,&T1�Q��#�|�U��B,7�E���KKB�����*x��:�6�F��%�B��
�*{�kݐNpǃ08�T�FK�' ����-a蓣����n���x��C��٢�&đc b0b�c�c ��py0�%�C�����g-�jun�)�v�w�!�X�j֬����4����fٖA��o�����g���F������I��/���s,ww��I�׋ʒݓu�e���j���I�&�E��7��|�����o�Ǌ��k�f>y ��z�^��sǏ��=kW
:�u.�9�[��ĥ���v�$$i�KP��P���X����jt�H�B�gK��na�Gn }'@�D��x>��C�0 ���7�BtV7�Kb2j22е�
�)��LI�?z��JL6\�/讷GRr���nO�����s������;5R�oBp�;�FO�ׯ��'�b���g,~7��S[�<G<���3��m���*���	88o!�A��n:L���w.��m�pb�J\>��مW�ƅ��qh��ڰ
c�,�e�q��QPۚ-�/�r��a	��H2�M�)�S	��cH{ْ�S[�X�L���@�\lݳX�}�̐��(�#[�x��.$4�X��$�䜳����!Ӿ	��O��08*N�ǲ�������yqN��MF��y��X!��r蟗ϛ��b��)�!��!C�0`� ���7*��ܞ��0 O" �/�@��mQ]X�vU�޵/�7�ŸACpp�,�=y�^�����ٝG���Q���գ���w೟~�;࣯������/��	o޸��N���>å��ѱ�e�a���ظt%�h��Ŝ���;Ə��+����Cرz%V͟�Uf��m9�N��]�#7$�
��tuJ!��p=<��'�S�(�r	�}�`ɻ����HQi�����H<g*o�|=p��y|���x��<�����c|��g�������hl����߶'/��>�[7_Gqe��-��N��ߴ0��F!�u�T6�r��z����cW|)v�[�M1"���K�^�{-�F��������W�y���
$�ˠ ��>xr�9ۨ.�"�*g�YY���縼; *�I�!h��@]�Ҥ9��ȱ"i*�{)��$1� I��W����*y�9�Y�A�pf����� � .�����ʒ3P��'��@�IPWL*%��=#�[���U�w�+�|���`��;XM�wn�I�J�OBJ�ch��%c�[N������-�������?���^�?�h����/��޵��ۯ��'m�����q�����c��@-mn�����xe������#a˞���}�L�y�]���� O\�>]�e�����V@�Ux��]�<3�-./+21�A1�eU�!;���0��'`SC`V��Ut��j	 =@¿9Z�3�����=����R�x�p%��8��pǲ��C/�n����l ��4C�<�a$�.���`�հRC�*��,"Y>����ɣ{C��v��AX��z؅��8�ⰶ��Z��)�卆ut�B�C���1t��	�WAִj�<E�ݐ5����@v�[���qD�`�(��g	V<��� O�U	��NHhBC
�چ�"����]0G��"-;�`a��X�g)�{$b���<й�FL]�Q�a���X�d>��ގ��`��%0y5F�߉!������:d*�Zu@^Y-�J�P^S��$*h�=��P_w�tximlp�����" �~>�bu�V*����+>	�	"��u�h�8�����(��R�I�KD �a2x����� �C������ۜ��;������#T���谫�A�!�⮵X��*���:,a��ݭ�K����l���P�rL���u��K߳šm�fL�9�5%0����� ��-�W�sxdk!��9`3octw"Ȥ�P�������E�i͜fy�,w������1!�MCMc	R����}��B�A�3 �%�a�%p����t_��n���}1o�d��w$'l�Ƀ;p��!:�۶l��u+�k���8~���>�����j4�]Cόè�X�([���C�$��h!�=i#�C+�#���-o��c$A�I �"}��;N����ǁI����)ؘ[�Z���B\\ᡱ���_ma!jKJa'�	�~�bx$*[�"�~aQE���()8�T����⫐4|��kY��f�\��z0�{���_8z�k'oܷq��$����3���E�ļ�1p������oO��O��W��Ǐ�Qi�-����~��+*����]\��c`�!��s��Z%W�b	�b���x,v�2\Y�Z	s?9�G��	SK�a�Y>�ִ@�%x1�C� L�>�9l�_2K~a��y��,�<�9�Ӟ���,�l9��te�͂�p��<�� ��9����/�➵�z,�˖�0�����%@���$���~9�7n`�u�/���~��\W�B�~�:���r�����qz�4Gg��H�4�ti�d�I���M�����O^�٤�8�ښF�e��ڝXO�hN��@��#���#8y�$�����鏍0�_���7����U�˰t�&T��`�S(>�*R`}B��G�����\Bp'0���n����v�BW���ʛX�v�K��[��RU6c��cx�����ї����'���;7�t�vt8����P���g��*�@a�Qc��2�@W��XK��q�Q�k;��w��d,�ȵ��F�<k�����l�s!�s���U��y������C�7��!��	�4˦z;{�9��6�0تg��빫����J����9d���� N)I�1���^��Iˌ|$�)��*�<b �	�̠����W��~B-��Qv�8�����UX5�Q���n���¬͟b���{��ﻉ3c�bj|Y���Rq�ʦ��!8a�V��=%�P���a~;^��W�cO��%y�_{� o�\��v�8n���(�͇���X��s��ʼ}�T3GG���=����#���o�S'�M��jo�]���
�L�g`�{�ܣD�^��������M�Y�o�1��0j�B[�W迧�^!����&ء�y^C�<⬅�-�v���n#h�N���\C:Ü(e�ݾ���e�!O�b����;�ټ�<zY�̐���I�؝Z�_l	�8H�*�#ı�R��D����%��<u��BɛJ�Jǭ�e�vhZ�ºa�賶�n8�]���B�eE`d�yP�
�X�b8�1T��ƳA��C�眈��@�U����/A�3��XEZb������2,w�2�=���a`L�����`�X�a3��ڍ�vb��U�0{&�ߊ36`��K1i�
�\B`8y�P������y�Π��?�Ѝx�u�B�C��Tth���ﬃ� ��e7�� ��J�p��"*(��Qck�<���ldHqP#��'XfW�5t$%'�FO�9���D�.#��ٚ������*��`�ֽ��d��>m,�8�x9�Ý gVV�rކ�e�cH�ܲ<�����2�V0�Y\���ek [�,!Z���ot7���!���q��yz�P%�#�Pc�c�%'l������ xy�i2�z��L�ivͱU��?���Q'��*�HK��C�r���]�v���߅�[W���58qh������fm݀}������ػo+.n^��zcah�S�c��@�Hkml#�,y^$�wH��'��s0.S��W�B����|#��^u�F���~���Ř�X������L�PM�Ї*.-���
==�D��� �D؄�	�"s�6�^��B��a�	� |��?|��G*��L�m�h|���La��3 _S9x_医2'�����
��<������5DR.�[R����b��~7r fO�Es�cڄ1�6i,f͜L��:�\�����_�~�w8��q�i�����3��{yj��7��ς��-V6�g������Y/��e9�۲��}�S�����E�%
��"b�MǢ��D����-`�ӗ�˲|��9��b��,�Y�`���xp���'��z(�b���qp��C��	^{�&�\y�_��ӯa��CX�a�n�!�:��Ǻ%k�k�&�D��;c;��G���op��gx����`V��G�ѧ��3���O������8�q��X�8xS�Q����}z�{1s�,ݹ�06�݃�a��#�7w���qG�<9}�u��]GP���� <�)�'^Ix���X|��/���a@,��R(���	��Q�X�D$�g�4]c���	f��hij�R��g_{5MO�G`l6T���� �Ձ�:�i�,ՙ�����r�sY��C7WlN�����ў@2�H
��y��Ւڙ�պ�5���l�㑵/A����y�%o.���CT�Ve�y�)�@B�g��^��q�/��i�~ؖ�8i��1�tb{XI���ZHm8-g�c��Py��L��T������t���9k��@]}�ʓU�K��㐖�4��+g�3K���k�����C������[�aÁ������$�ז�eK�e�d����̜�!��033333:�����4���������jG����Ͻ��<5G>::ا����*L?�K��Ԉݸ��?�����3�m���YKH�`����_����y�j7_lR�b����{�k(����&O���m�4��+'�(���ϰ��+4\�ӷ��g�%���'�W=����'�:ӌ�D�'�Ir�C:$,v�ǒG�WzVe���[�!0q��VNBO ��?A�/=4Z�ŒV�#j�J���*s���5˥�K@)I�Dи� ��/y'�[���@^Ο�<y>m���,|+`�]s�2X���mbwX��y�P�e���p2��'@�6��a0͙@�,j �j�Y���b5T�6��;݇�%P���3mo��DTҰ�)�C`lI;
��&�ݵEp�m�D�*��E��ʓ /}IC� ��,���u�Ŝ����2b���zL4$�{^�<�����E�n�l�u�7l�b�9�6a�­��tV����m{q��I�i؋9sga����Ծ2S��p꘽|���1?�ӛd��!��.�J8�&�'ȳ�4�����D*�Dz�hSSDX�#��U:{TXꐫuD��#�U���5sy�����p1�qdann.Z�h���8�ty��Y46�;�����0�����ߟ[�����x�B"C�q?,ys���%���sp��N�QX�X�f�yd4�#,<�4!����R(\�n'[�\�䅘�0Զ�F�V�b?��|�5���ɟ����X%3A~|,����`��M8DP�x�,�X17.F�έش|�/[�#�w
9ְ�7�����qo�����
���5.V�A�T�P�g!�Iz=�\\ќ�wk\��]� �G����}QH���QQ��
��9h�z��z�� �k�ѡ��9���������'""C����{��|���F��'�%��rs��������O:�J
�{m^Y�k4>�q�����n�c�÷�|'��g~H�l�P����'��	>4PzK�`gj'�3�-�b~W�@���ek ���f��\)�(��1����0|�H���W��9n,�'�g�$�E�T�}p����AO|�i�ڳ�C��������?!�?������?nA�O�f+����(Qf�@~.�'��A
��=� �H��G�C�"j�Z�0��ayȏ+CzD.���^% �������_zQطy/oއ��l!c{Ýkq��e\�v7/�ū'����G�x�.�|���o`����O/D�Y�+f,Gjh"���:!�=1^��
FeX%��ʑ�w] ��螹���> nMuM�g�iT��b��^Ǖ�G,^����1L@'�~��~�6�2S�������9��ج�����DU�Z4k�QT��)�BÉ3ض� s�������e"1�i�%�z�������8�/��ܱuOCJ���<�WL.�����x[A����G)WS��C��RC;H����t���	��x�#o��A��'�S�<o/�[	��k��x;d�a^�	��h�tL���xΰt�Wx����1�On��
�y�@��m9�5�r[�3Ii7��7.z��U�ɘǚzX4%�)><U��[ȓ�z �N9�l�
����c/�x���c���2|��o�<.kvi�b����������pd�p�u��S[l��!�!_j��B�'QUx?{��؉����m�����c׹����5<:]�I�a�cw-C�,�4A�q������<�<Y�iȊN��cy����y�*H���Vܥ܅�C�T�
��[���� �h	����}\D�"�jG�b��"�$���l��O�c�3.E��B��(Q�V���搨�*s�(��:�ey�y]	�����VC��h͓��<���^�����a_�P��4y�H��ɐU�S -�Ӛ5x+!m�������RhKfC�5��PyUA�Q;�28�T�!�\D�2�
���I�eh�E��p���yb���%�$f����cI�yX��]�U��F��* �ܓ�-�5:��^�Wb�ݘ�r7Vo�ǡ�i�l�vk���ҥ��n���Ħuk1k�D���@B|4��KP[[+2����E��N��.B&^�+A����y���UiG3�H�������J�K!�m�D��d����(tpB��e^��������vN�S��E�U�{j*

�h 	�Ǡ����Z�5�7�4#ȱ{�-xl�3�r��
��,�����1-{�·��`+����1̱Ŏ��nS�Dr�/�����ĤX."HD 8���*�s���v��@�D���:{nz88�����:��e/C!ǰ���"�VX�+2ұr�Tl\��W/���+1{�dL�<+�����a�
�����n����qxg=vmX��f`_z�9�a�G�+"�q�\#@<��6'8���æ�s�0m~ڼOZ��c���Lˮ��lv-���%�q�`����x�X��j�)�H7X	wn���g-ĳwQ۬2�R����ؐPx�=Q�s�Z�l�DH ���0Z���$1~H�����G�sp��^�雋+�Y����i8�������:y?����?�"pu�&L=�Aj{�Y8���@����dd�F";8Y!�(�NA���=�'�pP[ :�SFND��.N]��x1��q��8�1f�b c@c��o����N#̱�oY��R���������A�1e
6�Q��8]��¿1������yF�����J
G�~�F�|�����?ݵ���ǐ�Aj�
g�9R��$ ?��Q"P[���Rd$� "01��v	B�S �m݇���&2�N����ǫ�q��K��k����YZ������ؾ�(&N������*�v�	˧/A���i�I�E^T2����㑄^yu��u"R�`'7 �)1�t_��2�_mOl�y� /�u>xW�>�x���x��v�x���.4Z1�QKʡ��*jrsZ�={���w<���O�\����;���).ܾ�c����8x������Oߣ��i�օ�!��x���<���j)�V:ؒ2�B���L��iE��s=�L�i���J��g9\A��.�!u�@P׮���H� y��O�;��c��g�������f�۠(�E�dH��Pk<������8`"F�^�	�bƊ���j'f,������s���2
qiUԟеq5�z���'�Y��!w�ȝg�1EG`ZuAL��A�E�G����M^aڑX��N؆K1u�%Ȼ��=y��V8����y��������w-[�"/�Z:㔓���>�Ԉ>Aއ��qn��,%ܵy��D�];��k��E���V=�I��� 擄�)8Ȃ@K�Ap���u�U7�kv��ͰIS7j��v�g9�RI���Z������rk"nS/�<	��h�	��]&L9b&u�E��*w�� ���opg\*��B�2�)�9�ܱ/A5BK:M	d6��T��x�LZ䵄Yt�?!��mPS�F��5�-��[C֚Υ��~0�E�I��0�"�#�3� ��M�l���AU���<H�Ò�q˛�O+X�VA�_ǠJ�rt��<�P8��ٵI.Eha�NJ�����qrG�! �K/�B�H�o;�;��/lPH�Yf�M�N�����q�XT����	��p�m܏%;�a���X�a//݂%K7`���Հu�7bҘ	h׬9:��E���0u���1�{�@�!C0~�(�h�� ��,�D��f�ӫ̠"�Z!AOP��
xX������);�J�Q @�D���!n����9� k�x���$u��ƕ08p�!�]�mqjvF�����6p�ʀ�Ѫ�25F� xb�q���^��Gy),pX{ƿ�=ȑ�))I���"xIGBb�ib#��il�b��i𸺈���Ic�"�YM�Ga����q��h�8l�c��ؒ�VF=o��9cGbɜ��7{*�Ι��'bᨑؾ`>�oފ���b������������3�93��q�=[]���D�P��
�0m��<~���f-qj�"|\�{⒱51WoA����k���ÉE���x^����hC��N�X�@�9��aJ�^h���&1I����ዼ�8��{������ġAB"�	����Ą��E�3=Q�^�9ӤV�������}���Y��xD�y?<������1� ���5=xA���٩=��O�V(�LB�:��T��/B]Y%Za���8�� j��L�;a�4/m+R^�]�"@�s��%�XSV�ݧ�U/#����7C��v�0��6�~@�����6��Y���������-~y������O���q?���6Z��V=>^�<[�?�k���<���7Ý����X��-x��;��|:Kx�r׼ � }:�l���2tnS���Z���͊������[`��}X2v.b\C�m}=��>��pd�z�$���X����ܽ��|�7<z��}�+�����{�4�L��f5mP�����cᄩ��ؠ'�����a@]G�,#�<��zĲ���
/goثlP��	��"����v%@;�RR8B�vp
����kGܣv��!_>��Pk����jo����W�"9��MQQ��Mۡy�hҪ32��j�eM;���=*�vC���'C T���X���:Qh��)졐*h�C��>|�J2��&#<�\z��5])$��E�c�KO��Nbn^c�E�?!�k�2䱻V�9H@���xH���4~#�y��`�s����yI=8�¢d/,3�B��&/x8���I;����d�flܾ�����1!l�8u�&N���W�c㎃�7d
���m�i����� +�-�����g�����S)<�@�'���I�݃E�$�~���b��'�v�n��s}6�:1�w����;��"����!� ,'������7��[���������񑣰�;Mm�����_zD�k� <��&x7k+.N߉5ţq`�n1'o�7��{�����<�Y�cȚ<��9�`N��Z���x��*�<��.¦x,b	~,I[������DY2��'�b�Q٢����>CѢ�P4i7 y]_;�H�d����)���DA��Se���n4��5[lk��O�H�L��� o��<�CH���5�D]L��E��L���y��A^T!��p/�ڣ��������.�M�]�0����q���<s,�r��包4"$3!�X
U�*j�3D�U�pX%��8�qsQ�Ӧp�]@��P��A�υ�K9�Z������CPG�7�@y:ݗ�4s��y�fai�<1�i�R��&�4��~����|�"�;�G���c�Rt��S�l��+1c�Z,\�	��l��ѫ� 1����Ǐ��y�0{�<,\���ى�խ+zV4A;w�R���D�2�9�妈$�2��`��T��Z�YM��noo��&��K�e�8(����6
��Q�'�#\S�];��kgr�C�����]˖<�=#�1��W��oc.k�,����X8�݃-ȩ,��cǖDNH�/��vF�c�1�Ezz*��r�1���ii4��2�E	�3Gs�נ�wԋ�zVZk{
3��ho����X��	71� G�Vde`L�;�fN���a��%�8k6�nڂ�-[�s�Nl߾��mŁ��P?y"��%b������m�`8�I�p3�@����BC�~���[X`ٺׅ`���e�1h,����k[��{���pW9bH� �_X�{e�����$jT�P��,gODZX!�T�7)4�g�u�AJϓ��9�R��c�c�"`"�!�a���\ǘSۘ;Y"$%m;���5Kq��|�_��?��P��u���l�q} >����o|�� 4疭øQh?
D�0�o��	�A~HA�����P����'$aɔ���J3�����F#6(V@�{�(pQ�����Q&xl�3Z��~��>��-d�u�i����|y������f��X%C|�$�����?���؜��s�OK��7�,����m��l���3�q->>�6�%'<�+N�b��!��x�9�"A3G5�X�0w�dܼzS'MFMM�u銎��(#@O��*(èA#���#,9�n����D��}�sܪ5��{��g.���sX�a�q�0x�,��33	$6�݅SbȐ��ѽj�j�|�b�;Q�f�Kw�V5��NCuA�v�C����?O��'�aH�.Ƞ�{�h�#�Ϣ"!c	��F��W^:������ڇ�be@��
.��}3�;�d�"�X�9��R�(�i� 3���\m'���Hђ�x S:�xj-���{CC��4Nb�C�Ԛ�C㇛������qS78�}Jj������
aI�w��y-!��[�K�|y�E����K�����d��O05L�k��'O��Is�	������}P79����8���#`N���}�x��ٶ���vlغ����عw�܍�gN���k���>.^���n���7���+,�~���q����jhL8� ��ʀ�p�Z�xE�	��BRz��F�O�Swb�{�y��`���8�s-nEt��E��/g<�����A�n��0k��=�}]�~�W������X����Z��ԋ�������@�g��1Ux3c�����c�0p6l�'����^X�L[<�_X��2�l�!Ȓ�C0�;FԽf�= �O��"�n G�8����V1h�$lڵ'.]��G7p��5��rQ8�8��0����WLm���rX��@,P̕��.�e���Y����'�!ȣF�'�q���� /��|��u��,}+�;���j�K`��1`����~p,m�`X���x:4%s�,�E�t1/OU����Y0%��p��S O��n"�2�/�nǐ��y�J$����S4�thk��r��`�D�i4�Nr�t��%]�b���*�Vb����	�63�v�����:�5C��}Q�k$Z����faش�?w����]��I�&<r�̘;�ǌls'����Ћ�&V�hC �Mf��4`w" (�ȐF���^�&-I*�X��9�ng;��uª�&��-k��:�Er���
�E�g �H1q1x�Ο���2��ّ�I��~�9r�F5&6�c�cX��)Gg����xi��X2�'�s/^bR���VDc��`��O�c���A�8
��q�7'��A����r	.��s��n���4���F���8?NS��e��k�%[�g���7�G��s�M��%��k��޺����\��+�~�[�}b�R+;l71�	��콰�:��2Yk `�ż�S�p��:�=�����O��f��x0bu��݆���^J5�hК9tN����)��`偖f6��: ��D�U�V��]K�&=>f���pQX���\���� ���{�	�b#	�n��z��Q�����4���ce.;�_~����zB����7?|����k8�r�=�]`2fz����زi7R�����A-�ЭU7T�V�&��֥!'"��e�شj
�к��2�P�[��cfb���t��%=��ե��̈́'=W�z�ˑ!�([�"E�c�+n�GF˗q)����՟���Ѫ���%��n��:CS�׳4Z΂h��k,����b�''�\x;>�q�����m��Xy�ϼ��1J����ݹ��܊��+� dg�s��)1�h׼-zt�����O���ܮ��Jұytj��:v!�A��&�
Ms�q��%9y��_V�\��;c����̑30u��4#������1��XL�=&�ǆ��1g�|l�\�c'ΠC�:t�i�I#&`ܸ	=z,��[���b��EX4e����	Է�����1x$��ޏ�(���X��Ge�{^�gg<q	�y	di@����\G�@Zz�Ց=�P�\��s�Fg��#l�ppw��V�^�?��+�o���`ek'�[kgب�Йs
���B�YX���f����R�+,M�F��c��kR4	�乴&���kx,wC�����{�ĭ$n�qI�A�f�<N�v��OY;8��Q�5=I�$�K�ԣg_�޼������:p;a۞=�R��v���S���>{�k�/�����>�y���.��n�|Ҡ���T ��Jb6D�G�&n��CU}��t.tN���3ȓ��O�w����}0��,X{����ж�.��R?s�'NX��9�	�;ǐG}������o��_�僻89v����Ff���8��.��yl�{�o�o��{��|2��% o�78x�{̬�Μ�:$� -��? Ϭ�nD!��]���m0	�m�4(LUHɪ��U[q��S�z����£����}���!?��������8~��!�?y���F��}D#���i�$����}�1O�ъG���d<�ԭ��P�	&��@� H���3K��ђg"�y��O����y-D��֗�˧�"X�W�&�����2�4��a�у��a�N�e�lX�΁�l��3��0˝A�ͅu�,�&��ll�@�
�
�O={�;]`9lC�a��r�z)ː�Q�f.����Z�H�2�C��Q-&�4��i-gbY��`��|�W�w�I;Y���Z�-�䭳0`���]P��V���Ԭ���.��G�A��s(�:�A��1�:����`�܅�5f"F��a�����JK�Иk��+0Tj��{-�3� �K5�@��l�oᒕJE�� Nbۘ��D+3sQj(�Ӈ /-�P��0'7�S'f�s�VJr�S�'7��t6�t؝��=c��4c��Ƃ�4���oY�{�:�,^6N������9���1� ��8I�1��Ѫ��>�w����c0$��%�}��|N3��+������-Cd��^^>�w|-�=�,�#�;[&MdRX[h�43S����z��[�H��kز���c���0&��y��M�<Gj�z�jO�� �}`�{F��S�7�t��]����ӑ:{�hQDµ4�4�G��`yZ���,Q�]۶Uk���%�2	3��P�B�4G	�6�H��!�N��S��ō��g��u"@'H��l��H°�<jsA�t�I�B	$h��PF��ٓغh	lP��#���g������Ob����o�s��5���{�L}�G�Lq���a�p��-�ןĥ#Wp��-\�'v]�����o�^�m8�]k�qp�A\:v���wb�M[��[�aɤHO
ͬi1{�d%&!3)7���P��	�h)��/X<gwWQ��S�9h�x.�c2[�?sg�H^� 8�Sp�%?a/�Aρc0�ܒ>��>�:��������.� ����H��O0I F�I�	�����b�>~�<��8w_�lű>m�l�V.oƹ��z/z�h�@�e��x~_���+��{��gV*�عa�ƽ�L%0ۼ|�x~����='p��%<�|����mسn�l;�����=o�k/�Ɩc�4g#n�ڀ��7���z�Y�/hy�&|��/l�ӹ$K�qkeNo:��������xp�!���&����xx�6�8����׽��q�5<�{	﮿¥ӷE��+w���L�6ٞA���ŝ�L;��=���'��} �{Ơ��"�<\���E�K�<C�ͳ����\�מ��NX��kop���=�����_s��H�da����Z��I	���x�6�qV�julu�F{o��w�uX<:v���hDX{"�;V����TG0��@��� H�����Z�� ȽF䍂��dHA��M�Ón�<�敜�y�qX箦��5}�����}��j�.�߽[����}��>{\d�p�
�}�g�_�͇w���8}�&&.Z��Y]���j��SQ�d��"�i� �~A"q�󮄶p5,��5�p#�q�߂3�8���n�=���!4�"m�#,��
��?¤��1�\���k�cH�I�%�y�~X���s���	����$F�c�m>�?x��o�@ud�h����ɐ�jlq���<��. mb�*��nť�XY1��ņM����K��%�nz
���D
��!O�G��u��h�=�4?�v��E�	Op�PmSw�w��-G���Kܼr�^�����[|��;�Ϟ=���Wq��ٹ��!8t��?��wEB�Q��PB0&c�-Q�Y 죺õz�yt�ĝ���,n��$)� O�e�
H�'�D�R�ΐ�%Ϻ����`�"i�k:8Y��w5�"�Â@�<��>��.��{l*Dy3ux��:�2��r��mc�,���P��i�x�s��N$����	P�%ˬA���]r'���S��7�]h��s+h���.��� �95��he�vV���Q���`��Z@�D}涝�ݗb�>�X&�b���	�8��j����Jk,��}��+���b\D"F�c\y-��v��n}0k�P,0K��~#�r�L̬��9i�BP��H>.uc�fG�7� o�]O�	�+��V�P�1E���f�T�	�������NL�5�������T�� Wg)ꮆS��L0gOZ)g�OLJ5>�82�k���J���x *"� *
���HOMA��
��d�)[�8P��m`b���������-�ɇ݄����'->>�kc���r�Ec�Ƥ���偎�;X[5jƜ���m�y.��ݶn|섄a%�}����aa��<@�`���*�?��u<׋;h���-th��G�k$�.F���_��W,Î)�e@,��Ƃ�4�u��"+[���c�R��vI�8K���\BPC@�e�ؒ����}{��Љ ].R��,T;��fu�j�dlM.�V�$��X����%eX:t*n-ځs�n�����=ZҀ���!��`������w�`�'<�6�V�S�Z+V<�w�yy""�qn[����F�ɋh�@̫�k���~���߿��7o���{���!�M��`|E��_.�)$�,P��y�еM?4������-�Y]ʺ�ku7t���{�k���ܼ�Vv@MAs4��T%U�4�M��8�V�:D��IZ.=�� C����
��?냲{�gN������.�p�ib�vB���`k���H��hO�GkN���NԶ�VЙk�n�)A��VzLm�aE�uv��n]���48���V�>�|W;��W��hu�VcN��@�`��'|�����`K
����Z'XQ�S[Ӷv�bN���	Z��H�ĮSK1����s���8Bk��9X���"��N��x+kQʐ��H}q�$�N|�5#�� �� ���fp ����~�~�ݼFt�)=�bz�q��s,����ٽGar�A��u�tL�Gc��)�I]�bd�@L"Y�y8��Ç����	x�| �7郟�N��-��mu|�펿�t��_[���֓���z�4C��(�~��po7C�Ĳ��x�z<�V=
h;?����]11�-�4����ѫ����B�w"
̽0�>wc
�]P[p��3'��䋻���҈��\n��J�8�
%�����b�E��?�G_�g޴��st�4%Łړ��?8h�X��FK�V�MK�V\�Q)/UYc��7��b��?���bX��HKDG�x��ʇ���f9񄫶���$�v<��x���k�B�7�����B���z�����$Y{�G!mq�-	�|zx&���(��Q����z��ߺ��bg��;������.�ғ�8u�"�����;l�sm{NGN�~(o;������F�X��w�������̢��ԗ��4�O���a(k�J�
O�sKJ��*�CR����jwœ_`Şw�p�&|�+n�|��x���g	�;����D�ŴY��h#d�7�Z���B[��[#��y[L�^��O<��Ck_��
�W�x7�!o?�W�Ǝ��i�]l8�?`��Wp�N�ZM�Wu��C^f̚��C�+�o���vL�b�Z�����W�֝�r�qp�>�=}����������/p��Ul߶k�nAþ��t�&N����g�aǮ�ع� �LYHH$&\�J�dJA]����P$�"zL�7C��y�h����d�] �v�<��)���M�a"K��<�BH}�C%,yz!�DRb�B�\r��.��o9�Qm`�������@�7@Ա5Mk=ӬQPd�m���"͊4ud�á�%ȣ����MR�At-�ۖŊ�_��an��A ��<��-F'�l���C��C���\�)RLr
Ŝ�3���"Le�# [,�b�B�'䭔Yb���%
��Az5�ȫ�c�C02����C0�?��14:c�#1*.	�Ӌ���x,+�C��I&jL��O��b�D��3L��LAo�Ą@O��
	Z(MPnn�<�S�������NJX�vvqvv("��2Pb�C��%�hs��:=�TRӳ�D���p}<���j����"	�"��+�d�[�@]��(���0f2���(<bF�-C�����\	 	��SE
(c.��c�4Z��zǖ/O��93��b�։4l���E�A�E #������>� �k��y�E���x.W ����PZAof���Q�XT��-[b>]�����]R��O�D��s��^m��&%vJh0S�I���BW�p75CzX8vm܄�3f!���i4���\�pϫ����q�M.m������%S�"4ח�ĳ	�1T�
-�Tv(�8!���4Xu)����3�,��V}���mN D�ǃ{@���<o/ @�y!���[�X����K����1m�x�U�&x��*����޽{8B�����q��5�8�="���Nx��u.�h灦*�삐��&>�h���V�(Ѹ��k(�h���G5i�M�P`጖�嚻Ç� J�;3��]ަ úv��.��鬇��'JV*Lhq�(��������>
���`'�wĜ� ���\-����J	JK�D��a�{�4=z���[ͭH��2�$�g�V�.�j1e�`�����\݅�����lҘ.(., �&���1#l[���*�����+,D�0NX�I�S����	];�B��<?�H��S�1,M-�\�D��%Y�F��W�:���5\)���"E��L-,�fԏ�ktέ0q� ̘4�Y٢���=���4�C���̝��#��K��⬜MۄȭJ}a��^|��%��~NJp��z�⺵�;����͆��6#p=���X���� <K����D�����~�'br\sԺ$��S<��Έ��!X�@�=�J|p�1?ڦ�k������ 4'�"Bb���N��R;c)�u�X���!i���sO�u���^9��_: �i4p%h�r���3���-r�A���K�� ����ۋ�ĖP):R,l�`�#h' d��H�B���T�tQ�	�TEc����8b��Ƹ|��1U1��B���Ӊ$.���u�̽�.x,��	��@�7�������.j4���� ��p�n"$�K��mVt򒣐����7�,��*aɭ0g�Vl;xPTlZ�a3�wű�P��GO���Kp��e4�>�%[6b�ܙ�2b,�Z@RaD��ENe?t8Sl���'p��+<}�;�Gr>]�\O���2��:�l���A����� -�L�G<$ �)��¦�M�Lz��{����5�,��3-��A`s|뗁B�q�=���qБ ���� ��+��>��g�H����(k�ii�佻wG��Z�x��B�Nn�����ax`�{1x;���mr ����3����W������<N�,�?i�Hr�
������^�*s=�x�07��%����6f�؁}�/a����?zG�Ǎ�W��������_}�/����ؼ���n?�8N��a8r{��#gP��Z��+�6�m�
M|8�m�EN=L�wAC`G�'�'o�4|$S u��5<kj��ma���̔ O�I���"���Wt��x��K�HV̐�p/�6����R2֙C`�3ֹ���i�P����,{"Ls'C�3IbH2FC�E���:g8�������60�o��ZZ��uhG؄w��(���s.B�!ͼ���35�H4�Nb��
��f�}��������,Lq�|Z�Hj�e2,�[c9�J�ZXoVJ�XL�<�9$,��^e��*{,6w�|�#Y:b)��C`҃�oC�	��rA^8�i���w���Xآ7��h"E�	z�e�AA��9Z��_��A
u�l%�%��T���+Z�Pi�E�J�`�\|��t���v�NB^jJ�(q���7� a�KJ�n=�;59	-��'\�F,[�Є��E�s�c�,[�������vjt?1�1|!�#f��������Q�x?l�n6vQ10��qx~���(6��b�KJJBJ
]-� ����������||>���J�����V������ewltp�6+�r�&��䛩]�P��U*��m�r����y�r3zFӮ;N�?���aJϑ�1f.���m=������t�/Z�)�"Y������mƣy+����
K�hlQJ�\Bں!���A��pp&�� ��Z:;k-�CCL���?�w��������������	�H�M�g��}{�γǢo���|/q��#��}뇎�Y�|���c3Gܵv�Ǆ|�S�۱�x��_���ᛦ��<�O�K�uY-&�zd:�6����x�S������f�d�]���\���x��4>���Gw���(���L�|TG�6�d�2UJѳg|��)��ϸp� ��]"`����TF��䪷���K��_>●�`��e���E��;���ќ޳J[[�)"YpDd .]8H��_���	��C���c[q:!�Z$q�@(�?ݶ���ï?~�7�~�V�հ���B���� Ϟ�m;R���0n�`������w�y�ʋ2��s�)��6	R�U*q݁�nX�b>���/��i�z?<afb'�<)�<'�Q��%�#9�W��Ǉ����5{
�{3��#��Ń�П 2��$����1����F��ɒHזJߧ���M�?GNm�$��oF�~xw��8pﶟ�+�T��ܾ/&��� ;�;�bKv.�L��<���5����t7εH��R	�c�DR?؃��k�T@�?���[D6vЉ��(�B�D�b��%��:�����On��1��蝽��1:m�Ĥ��ZG�Y�ps2�@�<j��r�
q4����?�98
�<s�sy��8�1[��Y�~����-{JKK�`ݕ�]��4�Xo��!X��y���6<}=2P�G�&���;��:H]�,<{�,�`H<���	.ID�Y�W���I�4(27AQv�r��vf-.C��"$1�!��Ő�q��UQ�m۞��}� �<�G���ś"���c�1w�Vt0���PҢ'���BZq;���ɳ�c����;�����紼�7.b��t�G�-G�s�P:n	�*WBUM�Wr���d�W`Rv�X覘��hs����d�S,����?�������
δ����M�-yF�[i��w�3�3ɿA� <�?X�o#��y뼃�!�`��%�I{~��oSJ��/��D�Cޒ���2� �／���W���Ϳ ��_�'�=�/�+8
}���7#궫$���0r�r�~���~�[bƲ�X��{�^��;w}�<y{��x��K|�ïx��[{����wq��=�z����cŚ-X�q'J*�!��Y��p.�]�N(8�K�&��%/e���aJ��>r� ��yN^{H�����ɔY0Qd0�Y�B����]a�f!�!�ȅ�-/�V��-�G5T�ݡ��G�i0ѽa�8��a0Ii�8(�AU4KbX�̓�p̋�A]4��Q�c�C��
��m�
��:��Q}�X�A�\;�8e�ܐ�Z�d�t�B���L,1�:��r&8bz�	��z
�8`�̌ OCp�h��'m��U
���S]H/�f�[M̱Yb��k%���j}�P��@����&`u����5�DJ���i���O��ּQ�e3��mت��޴�.tN��ȐN�H��m|\���%;-�3�SH����9w1��G����)��EGD��H�����,/G
���a��T+��Cnv��[�ǐ���o��O����<',��K���dM�c��&��f<'���H��p!Fȋ�&pK�������>�
g��1�5���Ǒ�I�	��� '�zt^�d� ���4���=x@�}�qx�[;�i�o��Cws+�*0���Vz"�9�s�1��)��� o'A�&zkI�����<N~�K�,��Q����V�ā��Ӽ�v��px�2,�δa�D�[���T�_c�xG/�)�ă�p��`�ѹ"� .����|�@�!S����I0�iw��Vp��ؚA;t�jژ'�_@��q3����<ó)5A��ڟ�>���c��x��[���?�������_?ǺA�q���xl��]���O޻��D��H9}��/�����>z�	����v���=T���w>����&�ҋA��L�,Oo�YY�UU6��x�����B�漢�B!���f��,�M0vL������x��&�.�t,�Sfb�"W����pO�&e�����;Q{xX��ڶ=&�`���m�/4١�HOK��KG�׿�ó'W�u�RzCN�Қ*`%���(��l	>{�k�/�?��?c�qp�����v2�p㳵�Ve�� O,�7��� �7/�SmX�u��M`O��0S���NJDx	@�u���E�ٷa��P_�F햣��TVq0���U�"�㱓G�ptA�4�$"�� *���yp%H$I �&�%I�7�� I'�ﲨm5�v@+'d䵍-��qi�ql�7�1;�D�=|��-ֵ�;\�<�8s�ÆN}������x�v f輐OכK�X�_=Z�7D�orW������`��;:���E���r�~A��!��Hpq�Y��ԧq���޸��/c��mxN����,Hc- ����8p�s�3
G.sZ&vъ�{�?ݵw��Z;�Z�F���-m�q����ݵӜB�;,[B�0?2�+��MT9DW�UpSX�+ݵ��Z��Mk�!��I=iu'���'6�r)��*a�s�T��[�,j8�r�ô� 1�D�X��y�q�G8����%�q��%�9qG.��ޓ�n�A�Y�7��Щ�P�<�[�@i���{,�N[�i�6`�ҍ�x�1~�x��=���u����n�>��c{�p�(���AvQ)b.��xA�ɂ,~�(�*)9��]��	I�����]��(��K�������%,��-��a`���<v�2�]��	��:g�9�?!��hi�<�����5Bށ�#��7�l����n�x�T��2��Cx&n��MY��3�aa�,��+��ƊOE����å�k�;bNG�Jr�}��s��݀�oOǌ�4��O��c�����O?/?�����m�L��p���8p�6lދ%��c��ؽ�0>y%
B�x��H�K|��o��:h����`��Ť����Q�S	A�D�ۄ�p� ���
��������e�:�C拚y}{��P�BiO�g��^�'�c)$~y�=`���
��up%�^E0q$�υܻ9�A!	&�%�+�Q}��y�p�'��x��װ͜U��r'�4o"��#`�8 ����sI4���r4�Ļ3,"�.yt�CaL��T. /ҽ�DT�&�CJ't��D�
ST��*5y��R=3[��d_̣�~!��h�^!��J-Ub��D�(b�H�-�r�D-d�ĂD! `iӃ�����`�*��A�O ! ��1_��l��t�/[G��Ѵϑ��ao8 ��2��)Q'7C3��;�uq�A7;YPǫ� �:�`o)ܨ3�����#��	�b�5�'�����w	A9Y�b�g���ϱsq�B���`ǖ0N������jǟy}^^�(���1�%%1�%#33[�����2Х��Ս`�Ӽ?�P���ow�`����K���!-55�����6�E�n_v��k������L�u�pus��s$���fP�=5�Z#�B�l�R6��d�F�(�����Xci�M�Z��7�s�N����fz�k�yl����y^�u�F��?!ϓ�ax��ڣI~1����)�G`��I8�b'6u���8Q��=�c׌�0|"����S��j����Z���^(�����A��#��Hw�D�A�`;"�l���Hg����VJ+��6Z�����%[���}8�8�R{a�"�I��\�?O��w�5���?aߘ�8l�g&�xn�(��>U������⹹�j<qO�'r;���wJ;<4���!���^�]s��%a���H���A%�g�Gb��	X8���)�ѳk��bEm[tݴZ�8Ck&���X�p
�����f	�g���97A��I�aK���N$��Y����ĩcѴ� ���`����K	 �m�J�[��Ic�aɂ��<nƎ���H�y�`�@�����z=�*s4+,�ʹ�z�b�\����-�d�<H�ru�g�/���v�Ђ�m1�͞��s��0%V��������V������}�w���4�A{����@J;GW{Q;� �tt}@�O(:4i��{�M�n��l�ڄ,�̫´�L�HDG�7Z�m�F�C�=	t�9:���7U�����!1���!��b�=2d:��3=�x�OZ���9��5G��,o>�¤5Y�7�pa��J(F}F��5�����m0]�RN8���ݖRk<v�Ï���&��c��H)O�qF ]#�)ZN��kR:^��}�R�GN^x���I8P���NÛ�:�q�D1�߮��۩4P*K4r	F)�E�"P�8�w:X�Rgm�Ks;X(��V��A����NИ9�zږ���
9��J'J��U�s�e��6""�j�buF&�aTuT%T�Kf+G5�¶� �@��f�l��2��0��5{���Tڊl��9�6�J���W,���2w�~���$y�`��
�J	�<���{�àɳ���۸ih?|*��@jM7�T�CJq+���L�7����-�I!8����ԅ˸t�6.\��C�c�8u�()`o���{>'n���s�Ѭc?�O���!Q�@>MAR|��J.�]���$ͯA��:l�\G��/�t�k��s^�����x��D@޷�2�mu��!� ,w����3���Z��O�'Ҭ��L����������ľQ#�я��Yb=�.�x����qxD���r���g�⚹X?bV켍姞��fc׿�kכ�����.`����F�3kvv���%X���w������H ��ǋ1o�vt�;�LE�~1n�2l�y���b��]�Z����a����ɫ����N]��W�cמØ4u>��\��c�!&>��ی��V��)^EA�H����=�L��B8��%$6�jŐ;��L�S�dH� 1#85˄DGֿ5�Ѥ����2�#��U��
��� s-�Mh[8$��uR_����"�?,�@�6���0'�S�M��`��3�&CS4[X�4�SaUL玁M�8�J<�Qc� i`��GѺɰI���l��Z�R�L�9�ap�E��o9:�1�����k�IMF`z�1�h�94h�#p[B����(�i _.��yyH�]G���h�B�Ѹ+e��D��2z�G��am�a�]�B0_i- q��d��<��M̅5o�s�cBџ�}nO��L��<G��
-,MQ`E�9�e��_I�L
':GO3��I��r;�>Aư��~�4 q5���Ha�a��o�}����Xzl�c��;���Œ���h�c�����e����R3��o�B�,"�B�scEE�����K7��ɉ:UG;�Ƒ��J#%9M�s�q��R�A���q��1�2C"�%�H^v�ry3�G>.[5�b~���a4�E�*ETl���fR4w�X`xk�}�^���[IA�'�F��/>��mr#����D��K�nO����3�e�bT��X6b&�߂���q�5�h0�פ��ǌ����Gò��:�u2gT���h cY��^UU(�H���)����HF��7�2�p�鵶�ru����U�n[�0��zx��@ �+ݣc08"}}����}"�0��������+�d�&l/��)K^ĽP����I �]��8�G�θ-��.��{�?�R}G�'��[?|�) 6� ;��Ձ	��A��e�Yyj��D����=|l��E��N�JAP0��]*3Afbztn�^]ڡm�JDS[��Z��}�vv�$Kpv�/)Y�ެ�����уѲE%-�h��ѹ������ؕW�zW]�����ܖĖm���+�vE���2:e�a�`e�#5i߱���Z��Z�G��ݑI
�Nk���tm����LQ�J*AN|���mZ��Y5"\�rd��K!��z��t-�R�?�8=5ehQU���4x�������k{a�u�>�K�G^BR����H�A+C.U��}m<o�W+��R~3\˯���&�S\��%5��U��J��*�����>
K�����y�в�m��s����58�X�oRp�+��IqY�;:LĚ�������[��=&sv��ȅ��b n���\� 4�t�boz�Z�ux꓊�mC���o"s����f�V��sh�}���wN�x-�%ȳ�]��zqS���r�4���L�pTs�;�l���N3�� z��r5dԟ˩�7�w܌�uS��
^�i�L�3�mL4PQ?�s<���*LDNN����#�uh����X�i(�6���l��I�h��ɑ5P8T�����
��88��w,T�� �{�y�B-5GRh2cR�2��D7�p��A�9������SPU_�eI$>}E!������(Fla�s*�����fȫ�.C&�z�v���g�mO=v5ԣ�a;��َ���s�>8~�/�kL���)^}�n>y�G�c�3<s"қ�JD� X@�4l0̫8_�	1'OVB�S~� �
A�������l��<�Vￇ	{�c�ҫ8W=�+�����A�2W��A�G����<��H���C�����ŋ{7�w�p����:3�����] ���u����Et	���W����E�<�V�g_b�ů0zͳ�	y��ܵ��遜���4�E+�ޛCb��cp���L���?�����;~��<~��O_Îm�o�8������������!���m��r����T�v���c'�iG�N��q�c�ع�i��vԈ,!u����J^B%� /����}bN�i�x(=�@������:H-\D;�&��8H,� q("�k	it(c��o;@��
��0hA��Ж���H`���:���A�CX�i#�)�K�1�IRƊ�Zy��a0�z�Ƀ`�<V�C���{A1
���N������M0J/�6S$C���G��m{�ǜ�1�l0:Y�a��&�1�ff��ɎޘG��B���,�LF'Sb1�z��,��n��@��B'N��)WLt�N�df�L���R������~,�u�@�p,R�	PX ��T�ʵ|�Bml���O�H���C���G�Jmے����]��1G.�]���j<�l��4 �*D����U��֕#����l�e׬7Ql$�@p�/b��D鵔�8�cH[!؋3vw�4΁��� ��gt�2�1�}k����Ǡ���)R�|�I\9��_Y��g77/TVTcҤ)"ipNN��̱���%��]�y���(�5���s�9�
�G9r��O�n\c��j������nA��^a?��}���RD��c&.�L��^X�揍V.�"�b;r{�MLE�9��/ۻc3(�%1'χ������p =S�)����Ҝ=|/��n�̷�П��(+D��MZXᢻ/i��X�vF3�h��7�A��rr�W{�\��%���H�mk����3����xq�����z�>^rԪ?�mO�\K.��L�&��Dpv���;xc��/��E�tp�[{��OH9z@�]��͝pKA�̎�π�.�.�!��	�3�wyB@x��{(����x���rs0�� �%�9B��H�AVR4��p�,��+t	�Bw??tF��Z��a��K�PײAM�Nr�:�`@��	I�N"Xş�;һ���-���I)�ҒD-��\�N��4\L�B� Q�&��9���*,@aF|���7����(��E��@++�H!�w�<� -*��$-��\h�RWwt�D��8���@��֥�(.EeV>�C��L�K�C�' ��w�ϛՠT#�/%��(L��1�5j��H�q@���Z;��Tp���ai�zo���O�g
�eo[<��ҫ�<���D	�[@:��к�L $��m�J��Z|�V��hK�M�K�R�����ơ�8�`nL��oV�Ç�'pj��*莇�����Wps�n����x�o���#��TzkLR��J�A)�Q��Ց2��;?�E��wQ����SZ�wÃ�[)�ϕ:�t�ss{\����i_W�A����æ�Xqk�����B��[��a���X4k"V.�����cͲi�7c&��-d���ܫ5�wk��[�W]5�jKѺi>���Yi.�4-A��2�j����3ЪYr3b���_��2�1��0tk�	����jL	+A����4Am~R"[�̩
}+��ƹx�~����i�$(=� ��@N};[���I2�A���ܯ���2�MR�I�A��
lJvC��ޅ��g��Y����j�e��}�X�_�����Gq��a��شe6��B��6�ɦ�=��W�|�������`���l3��Z�����8x���DsM��pH�i���yb������������u�<⡶wa�������O�7��1-���M'�w)�!��iy[}q�5��|qv&A�ߙ���oF:N�'��_�O��o����?�����_��+^޾IZ�0l��x�J�-z�w�;�>:���σs��ԍ�1�0V�[��Ob�އXu�5v_��V?�K�D��!)����;�	����i3z0�\S.
�dt�׾��L���4[��_��?|�#�޹�U�7aݮ���9���bˮ�ذ��V���Ǡw��Y,[�c&���)1a�J�4��\�L	iҊ��P��(�Ɛ�N���� �5C&7h��u0��\#"�X󑙹�����O����:Q�VڱѲ�������,R�(B��6�!	m��ΐG��E�`X�qd-W��䎇4g"�i)Y II|oHb{A՝ ��hD�^����"~:$1��H�˴i0� &�m���N�琍d�\�wY��{��̑[�\�1j����Mq��B��Ԕ��Jouj��YF��:��'g�#��d�<oݓ�toxN� f����8�2�!o��Q@�B���b1-��E ���O�ƐG��A�A3sk�rpB��VJ�je���B�N� S	�fpV6}�2���J-\zg7�X��
,[�h���EZj<R�ch�(�.9�ݴ�"*��]��yvqKz�7�k�x�Q�u�V9��Ԕt�O�6�زƮR���b��+2<��t��+1q�L�4�EAA��$���	L��5�d�qTa�fը���g��Pǰǐ��y�8�ϝρ�\I��{\�S��Hx¿A��	�,L`fB�F�pP@���	F���N낵2~���ѳbw�	R����5�h=[V=IB�R�<=�&�  ��F���F�!8]Q�M~8lBZρl�of�N�x��%j�	:�(�9���E����-bÃ�w�����e��u�И���D�
��g�ּ��@�q�m �O��u�x��=b�$�?��U����H<����7L]�F�{R\#yh�F₻z{O�.xe�{�I|*w!���$�B���� �婥+^�Fb:�'�*a{[tD����bÐ����@$!�@��G �G$`'A���hTi�I��r�FVB� ��(��>|�tv���E�����p�����g�#/%��>h�AZ����18���|+j�	��<�A�O%(<Ζ*x�Ub�`2�?��.�����,�������l1X[Q_ㄉ������qF�X��X{$��In>J3sD j�w��3гΰsA�Ιڣ�m�0Gy��,+���p�}���d;:#���좵�!����6�CNr�+J@����������
��7�Y�!$?��>	�1,���w�Y�20�G��%��%�x���J������i�����`ۖ��5o=��X�/�]���װ��6t.�ř�X1j,����.��d�=x[�����b2��M���X|i遷� ��L�fgo��k�$eǋ��:�j[<���SR6�ػᦽ+�j�q]���4<2۲������[�����/��xr�<�}�^_������ח����{y	���������xp���9��wO��ͣ8{t+��݃�7N��㳸uw����6a��NyuY�׶Ơ^ѫC����Im0ůu)-����J{�s��ʩ���$�+�3-{��m8���!s'ȓ;C�4���-��$�� .4\���7��ypJ˂�4f �8��s�-�����-Em۞?a:6nډ����ޮ�"mRÁ�X�z)f͙�9�`˦]8t�._��;�^���p��k4�������m��J/ELq-��z"4�t�M��)��}"�41t�yf)P����� ��Ϋ��%�!�����/ܵM����ϱb�M��� K����qx�Y�����&$��0lr�/ؒwn���_	�� �I�����<��!���x�(���wo��煷���_��p�6���D�
+��8�mC��W�Axd�G�Ey�qc�~,�]�Mc�b��'Xw��9���<��W �yI�-�J����蝆4�1�BU{�M��K �z����C����{q�������-{�h�Ī�įx�����k���8w�>.�->~;���J"�s�a��ذc&ϟ���gb����1d&==SI�m�"u4��p��%���2{Ta�MH��w/���	�d0% ��.&*=+z���y��̿3LC�C��6����VQs�a��	�b��"D���a0M
e&5�P�O�*g2,�$Ȫ\:Ǣ�B�sFC�4��ˡL_E�R����a�9��a��5�A��L���E�į=&Ģ?`Ѫ3�	�� :���~�U;���c���`�TX��v�i aa�ca�ca��J�Ub�]M�*�=���\=����4�	����yA^S�YD���{�rp�z0�%0�n�����2S�2�b��D!G��,�Q��@���:k��������2y<_K�֘Ƞ53�=[������2;;���C."eJey1bc����iQ�"H�a��m�A���U�s㸌G�r�V^����S3DZ�`�H[�`��ՔLa��D������ry)NZ̮ؤ�$�>7���_`����I���x�.�	D�7A"'��\ٴ|�7AtT"]W(��n#��9𹲫��"��6&j�9{�	���	��Z)��j�o�t�
�k-j��7=Cg�Wǖ�$�����@����k�o��EO��2.\������-Of��u��,�eh"���2�G��;o\s�9k��
�a����;>C�<S�;z�e`8��ء��g����."����B�w�s'�ss�Vc/'����~>B	�g��قɖ<Η�� q�$�H�ڢ�9i��m�p��P|u�,��\�Ñٸg�7<����[���P����C�A�i��jO�1��+�+��^�r�����T����xc펯���R�Tj���nFg�?\O7���ey�Z6Cynz�`kD�����l��I�2�0���������Z�C��"	����FJB�M��-|���G���p�v�k�Ҕ8��N�D�p\uy�;�b��3j�ȊAfZ��C�"�`ڝ޳l�Sl�dc�0�rNgd�6D�[�Z4��y�V(��D� \��_��ovD�axbڤ%�YI!Ǝ�������������ƚ�!F�=��m�R�S�L�<��uF)+�*Sd�g����C��6�9_��KKХ{��n�H�.��moWLr����t{L�60���\яd�{ 9�c���lC�6�)�w��G�(����#��B���lv.�?�;sC�r�L<8vy��h城��¥�PM�w�g���j���5,�9�
-
��(7w�=d68aO�Ǟ���˰Llr��n:QYJ��S0�;E��ϩo}��GJWܲƑ��1�+у�`V�.�r�o����׏���c�q�8�\:���v���z\<wׯ��gp��iܸ|W/�ܸF��~�o�{�q��\�r7�������7g":�o���UB�l^Q��5�1�iw,�m�y�M18��F��U^'D�� �k!.����ސ���k,��>�5�6App��mZV���lE��#��p�Zۊ�0�;I&�����l�:m@U�H,_�	{��;�z��nݍm;����r���ص�����q��m�>t{�\ł��Ѯ�tt�?-;�FBV�(�ʖ��c���l$u��5���g�$��!� �/�+�BRy� �4$ŧ?�k�B���mnC��Z.~�E��a��;��%N9����֧����P=����~�<� ﯿ�o�
��5>g��F��')�w��!
	���|���/���=�?��"�Re��֎8���[�@|��'��x��o'�ƕ9{����uw>�����p��]����'ȻA$K�����Ue�3���L� O���h>y=zM߆6�b���j�S������?������B����>Ε���7�w����+�nag}��ހ�kv`Ƃ�X�n�(3}�
t:	�ԸH�6S�@"s�$�;d�; ��i�>H�wA�>&~�P'.SY����j�=R3H�+,a�q�L�,�ݚA��	�.�u�<���`�n_}�����qhC`�1�t��!P�����,g��&@�1^��2w<�Y#��.�"�挣�I�rHS7�,���`��ʬ�t�y���C�{r,��<�C����|�m��茡���$mPX�������X@���Ă��D�޿ o�
�WЀ��:�$��yc�Ⱶ��/��y��}G��b����b��y�Y΢�O��	���@Ǡ7�L�ԉW[���V#��ε�K^��N$[Ѐ�V(�	N��I��B�U[��F_owl�������oWy���b�p��ċ��d"U	������Mǀ����;�`��Y�G��2�E��#:��,]�����i�:���UX\���&��K@~a�u쀁�����Տ��kOQٺ���"���cW'��y���|>PB��%p!�$��4+�>��9WԸ��	
��K�����ظpDFBea"j�r�s5=A_��M�&HK�A2AgSRT�Y���&ZZc���L�����a�ߗ�=	�BМ� �1����F=~>o,l��&#�R�q���c;/y�h=[��t�E��s���c��H��%q@��<lH�V��`�������ھ#A�?TrS��� �1N��pq�?ݟ/_{� ��Qt�C��E���Q�2`,�^��'vcOF9n9���K����'�k#�1�=37๊�O��=����o�@�r{1�TK�ǐ��V���'�-�Q@�1�@,��ZTvɠ�4f� ,�;�gL@�v��7��cr��1ǐ�  ��IDATW��'m�9��������+���3�X��v���dRJ��hm' �Oc��];c���w`�tj�V1I��k��x���/nvغ�X�AQj/��������(LL@ ���w�S���D6����L���D�	���:=S�	>\� ���S񱘔���9ؿs+<���Oc�����Q�����3��ɰ�����N��������˷x��!�u�$ /C�C��#�T�ȥ���6K�uvvm�,j���ף$>�ڢr	|���4:8�hsPE���3���WVIQ��[���|��O�
��2�����јCm����X:}&�t�0�=p��Ե뇲�j\���[��C~dJtH��?�Wܽ{m˚�}��%RF���v�E�P�r�eɾ���/ڛ����C$��et�7���1�M���*/u�" �Aޱ�"��ؔR�^�ص`&~��[�~{���ąS�q��E\�x���鳇q��I=��O��˧p�����,W�����i��8C@x��>z��l؎���b��~1j�u���$�+��̚^X��s�0,��a�h�WG}fs���5&B�g��k?�z��{,��Խ)|c+�m�(t�=e��Qk�����:e=4�xD|Ӣ8V7 �O�ڄ-{�~�a:t'/���}q��~ܻ��x��[\��k67`����:`���B�ֽѪ�8���ޭ�ؾ�<v�;�3��νG�������̀�-��%re�$ɐ�������#��k�A҄��w.�n����XJp�������'�����x�Q��s��c�ތ��� ��d��_	�~�������o<�_ O
Pg�u���������-��:	h ẵ<��(i� @�y_;ⱀ������6`A�9X�	�6�|�}g?`����s0)8#��J����� �b=�rH���ǵ�a�6c�-ز�<v����f��������;���F�3��������b���_���Sشe��������k�����F�Q3о�X�V�Y�q�!�E�6(�`��@f̲A�G0���c;��	���r�e?2��O���Gd~I:�4��=	����]�
���� ��N��IR�@�:D̿3�e�H��B�7�1�6k4�� ��)�̂y�H��@����E�$-�$c9�2�,t�
xX� ^��$�ht*��+o`��7�q�����!�)O�ycr�Q�\;F$6f��B����m��R�� M?	AA�ri#�1�!���!o1�㱭�Hy�ؒ�y�b�$?�<��M��b<uvc�<f�-0�T�&�HU[��U��sЅF�Bsī��5Z�8��9�7O�0�U-B���q������A�c�,[�DN:_�Ƅ��&g'Nڸ�,�:�Sx��	�7��cw(���䚚ApԻ��#���;h ��`9j�P�_6[w���K�m�>l�w����{��^��h,���$��tZD�ƢK�^5r���@X`8BC�c���ym��d硠�	q
�k��FJR��TgQ37�f*�ȥƠǓ���ŹȜi��^�\�{{T�c�@�\B�@�J����`�L3-VJ�qP��5� l�Ψ��e�R�(=��mS�`7����z�n�mq��{d�I
���乑�|�yf6�A
�#� ���D�T�8�mm��g\	,L�E�\{+�]�+
�[Q;c�'�de�H��U{����DjS�ͭq��7lpd�$<�rV+�`s|���7/tyO�nxb�*�A��@�xc�(TN����-���N�mj/�.��h��/ɭ�@��k7Q||	݇2S-�t67�'�������/��_?�̵�hѩ�33q���p��J��C�I�P�w��y��3k���a�^S_�J��.�j��N�vvϑz=m���W��üi�HL�0�(ܣ��;�P�v�� 41x��������߿E��"x��}�wAf��B�gs�zٻ/~��g���蘞���Q{���ϯ�}p63	c�#P���O�o%��:�3����C��6��G	��|�8��ʬ4<�sK\������6���M(��F��3R�=,-ѧcG<~��F�����(�ʁ�����Wd�"���F�����L�o�H)+%E�@i�"��^$�B�}uN8���=��Ɛ�K����/�v�nD�#T닲�<;z��>Ƃ��	~v`�;X�� p+�5���g�k�	䄦 Ȝ�͆�A�\0=�>�n���7�@|�.����hK�<���~����`��c$^*<������ܲ�Ѩ||6{r:��s(�O���_=ǫ��q��Y�?{Ν�իq��9\�u	7�\��K�p��\��^����a?��[���2�!稽��(%z��	�;{;�=͙3GT�8y�2gRʓ��� �Ln����T�V�Eh��a!�0u�i��1�9w�ԥ7I_z&�!�� hû!�j<�j&" g0����_?����M�i��RV�ƣ��*ߏ�^G�m�,ذ�yr���_}�s�����Ǒ�1c�>��e��!��*	λ���V���k��������ƫW�p��E��x��1��z����P�%F����H�bSNc��V#��I)W�8-j�J����݆c���]���Ħ��`_#�]���C�[ȿA�a�����w</��1��~�0��i`b����7�����A�_��;84n$�E%`���m]p��[�`|p�m�7�D��ڵWĢ6�~��O����=��]��!O��8��6���D�&1U��p�>>�{���_�q� ̬��Ocݎذ��\��o���}������w�
��0���>~�_�{��#ǰ�� Vn���������+X�m/z%
.K�.����u��P��4c;$�k`_�A�W%�qt�� ��@��Bɥ��i����-LT��Xq�(��C����N��t�"���}!����̣�<a(,8eJ�@�IdIC`�<��;&�#ż<�;i>^�(����Ȧٓ`�3�YөM�4�@1a�I� I$�K_Ӵ�P��~���)@�S	��`�AL�x�w=��_c��El�	Z/�o>[��G�;̓�a�֟��	�>��%Թ2�-�/�����v�-(l����\1���o�7�]���	t�񴯉&j�����P!Ri�h��h��5G�5i��*Ҷ	@�
x�I��"
LI�"�6�yY5Q���|�\����=Ŝ8�iױSk,X4�w���1C�e����!�]����"�Op����Lt��I$N����S���E*���h���gp�@iY����)uW��8|j?k��0s�"W���[z��'f"(,F̯��DzF"�����6`���h�wkVm���#1a�`�Z;�ԡ�<��U��-jQS]���$�� D�'k^vf�>a+#[Mi�d�Sҽ3Fűp\^�$ ��Рgm�ږݭ�Rdi5h�ס��=z�i�ME��34������@Z�E��y���0B��Ծ6(	~,�p���C����δ�-yys	z���b��]�
	�v��x���2�Jh���h�����9j���,l�d tsjwo�zQ{ @a�S7o\���\\�O�Ն�x�tv��{e�y����y,�i�\�䖹3.ʬ	���D�[�W��k�%�]S�3��z�^���1$��75J��"0"�Zo����p���߻��/E����RY�#��iI9��Hŷ�e���L���c�	k���g0l�D��"��$I�G���HH�'8��姵��p��i:�%��!',㢳�:*?�F�s �ƣ����L,�� ��nG��-(JI�==�$��r_aq�sqG����S׼��É3�1}�ldyyb<�Cws
�KN1^%g�d�r��IE��c�Ǯ�m�N�l�Y�#������fj�K���I�wx��A�8y:/^���y�����[hQapGQ()l���L�\�+�mĨ)��oS*�	 ]\�B�@4��4�M�.(!���BL)��x���V�" ��S�i];�
��k�\<n> 8q������3 ER7,�O����<e;�\�1�v�n<�#k�̖���,ze�D�ʀ<�Tjd�{RD��X�7	�u�Ɨ6!�28뜼�F�B����A)R�0�=w��s�(=qW�F�Gm��G�s��й8Q�]������R���ꦭP�S��U�Ь�)Z�h��kѮM-Z�6C�V5hݮ%��茮��0�@zĐ��ۣ;��u� ���Æc���ٽ+�v�&M��C�n��o�R�Ej���,�0˒[c�W>��=k\��]�)�ȃ'1t�Ե� =�J�e $� �'����_/H��A8��'��N2��m4>�I�I)���}0-ڏ�.G1`�q��?�#'���������9�Э��WtDlA[4��~cbѺ�8}�9n?����+^���+�n���x������޽������+��f#B�[��2R�(̉'�X����]�W�T��}r�!��}��ޅM��h>��y�M��a١WX9�n��7>e���St-��u��Q��1���ԙ�om���-�/+�߈�����}�G��{���#ɷoH^��g�wo�?~.�77n���QX���j=�ٹ
���'_���U ��U�ͬ-87?�^�u��9yy�ϿŸu����$͞ȓ�^�4'�.8�.;�v��KL	�B�Y��{����زk3i����+<}�
��_%���������Ϝ����~�_~o�������<��_�/?������������_p��5�_�))E��`��y�z(swA��f��aS�
����˝- 1#�Sj�o3<Z r\�uL�s��:�<x��n��G��ehzl�c�2�d������Q�J'�Y�a�SL��h2�DH���'��4eA�x�ƍ�Y� ��} ����%P�l�Y�ȃh��:m.�Z�c�Ř��6&l��)��`͙W�6|>F��ָ	+��6#0��si@�'3Q���1��y$x�+�cw��$��2�;b�}���w�-��y��3�l�E��I2��7Cf��4x��N��L#2�'�: �N�d���h��rg[9� �kv�)��}s����
J��4֖�pr�V1v�:�m�q�Eii1��[��ɭx��N�ލ�b1�/1)q�4`D"<����l�4z"'7]�:
���!ȣ��#c98�݅j�F���
���a��=��`-���#�c����+*��.������,8�p ETD���`����w ���R�:#��B���x��&�]؏ISF���L����FK�]+��@���PW�E���u˥��4@�p�<��DT-�D��J��,�5�͕��8�"����Հa!(֨PI�ϖ)���ņ`��3̹K	��y�%�-�A
)�	�6�r��w�>�%���`�`Ȼ����1X��n��Q��Hq֣�'�QgJ�欝�V�^��z�f01U@A�K���Ha&S����Ƈ���A�qy�r�O��������3x�x�'��C0�\��y������E�K�ib��jw\2s�U+ܳ��U�]���:vy{�C�m��ٹ�]P<�(�Y	 +$	P��bm�<����4m�M���<-�SR������N�
E'�C���E��v��ж}G���!�/i���l����lic�pj���he�7aZ��F�f-��Ug�����P< `�U�#*k�f�@�6ѿk�ef"6$�q�h��2O�������pĻ�
��ۏ@l�\ħ��Sg@1WT���T���a����<$Qt-ڵǒe+>Z����OT����EZ=J&+�y!"�1CG��]���g+-.h�fvRI)�wB;R��r�о�Z�SL���G\��wZz�P�S&�F���q)���6�K�A�`T)�9���UjQf�T�Rh����oǔ�eD��j����e�x��sp��=^���ݧ�xn'�)����)�8q>^v���8S�+�y�����	�蛌KNḥ�vfMJ�>�Ұ��o��1�Q_YA�yaxj�{
RBN�&��C0p$*o�MҞ�䞀� (	`���n��'��m{X��wKG�S[q"���R+�3�л�F��fi�/�8��B�7��`��7�4��Bm��&r�킼�Lo3�;bA`)��S�f~7R��!Ϲ=AC^g�]{��ܽ7���!��4a�!� �A��u�4&��!YE�n�J!K
AZF`Ela�م�^���8~�")���9z2k� <�=����� ���;��٫����[<�O��������;yǏ�Ľ�����sܹ}��=��SWѼ�4X����:�FO,	y���n�I�Qb�s���	�$U�	�B��.\��F�ɏ�p�#l:pk��Ŷygq#g ��,�7���	�֒b' �����/�4��
�xL���K�o8�����W����?����O��_����׿�8�v���	�V���6��#�q�T��vl^�چSbV�EX;�6�{�m���������1�;��<��������T����b/̂�P�K7I��
�a��c�1s6m\�3���ų8x�8�]���O_������.޹��gP�n��7_~�/��	_}�~�+]�t�����_~���މ�2�?�2�SӪ�$I�ԩP��I�H׋R)���P���FH�C��Ő�	�hp����@�)Q�TM@��>R��^�`TG�׃ �?�lU�'ʰH}h�_(�:��z&!{�U;�ɐN!��e���g��j6��g䍇$v$�C	�C9fa��h%�K:��`��]��<�4!�<h���k��f��y�n�[{��ƪO0u�\����8�'�ՎŔ6#1�ɍ�N��
�.6���p�<#�1���TBx���]ː7� ���h,+섑v�����>#�-��<�o�AoZ�&�iО�gWJi��tnl=H����#�^C�*�l��S#�B!�Oz���ũ����u��2��Magkm��s���6G�^�ѧo���m�нg;���p�r^9Og�
5�����vXi��w������k,�Ő��4�tϡ��霃O�Պb�Z��c��/��E�$���V��$��Lop����3�N�HJ�9�R3��\=+K;�|��M1vB_��ȶ�M�����qvz��w@�Q�-[��9�8͊9�T.����l9X�T.�q�8�>*	�_i�J�<zQM�.z�' -4ء��o.�zo,u&�k̷ǖU<Z��%b����yl�%�<'?����"��dZI�)��V��=zVT
�3Xi��*$��Xw��6JS1ǐ�l�����"��C ���?�������>qww'�	!.�	�ݥ��������;
J�w����'�w��y����Ϟ3gf�Ȟ��-k-Oo:��ȉmys��N����<?p��#�p2.��vA����S���gyOL��o��3�����Qٷ�ړ��R�����؁;|{�n;Jel�=���<y/"��e��F���f�PE���+R�Y8b*+筦{�.Ļ8i��yUСz�
�����O�3�u;61u�8Z�
|�6R��ںi.Fʢ��׶95�ߠ��Gw�i�Z������c���kso�����'�9�h͛�f���ܤ�;��F1�s{r�}�ia]e�`jIiH8��v`X�~,[���s�HZ6hCa`�F�d��%�d-y_�&'3f� �|W���Q�B�N]�V�H���(�m+ in#����v�X�x�vncĘIU���LL������L�=��?iڄݛ�is�@�:�Ҡ+�Evu}¨�{Wn`K}#G��z�ml�^s'V�q�U^�Ć�"ڛ9�P�O#;iԸH^ԧ@�c��˔J��^�G��<}��׉%|�X���5y]ȗ�*�.��R�����)܍��yT-^�g�E�4^TO�Ip?D���!�k�w���K�֓� ���)��ZO^��W
�;G	�J�A򧱫@��ߐ���.e6fY|��&��KSo�l�v�����[澸�y�i勿c ��}��~F
G��$�`��E{��F�4�}�<�#｟W�Y���F��Z
F�'ѶafI#_���"�W/�{R}:w'<�>�.��~m��I��ӹ
�����U����K��==�1�'���.zy&%���#\��<5RhU��.s/2g�y��EVq��^AS��YKr��C���Jx�����,|q��--b��K�w�2���������{��oq����Y��9o�d�ac?tr�eX��Ģr� �pN���yM�a��6~�n�t�S�z�ڽ�X~�e�e}�+�������!�pVH�X5\��6������5s��龓T�N�Sz��?����o�Y>���;~��������yT�H�j��#l=8���g��|��M�j�L�ϳ�[8>�S[
�=Ɔ}��|��νdԊ{��P�$��_� ����"����qn��8!t�D�p1w��������#�Y�d�d���gɢ5L��H�okV�f�ڽ��{��go���Ev9�Q���Y��(�w��������*?�o��wo9s�
M��/�C!VEK0�؇.}3z)�1�Z�.y����`�X#��*��M�K@g���YM-2���T�6�k'��Y �;FQ��$�wǸZ'�[kaȌCZhú��]1J�i�8���`P������D2I�������$mn�.a ���J�u\?��:bQ)j�i��K_�u�v̳�a�E�5K���������|O�Ȝ�X���F,`�C�,4�ک͇1VZ�� [,��5u6cVU��EyU�2��؃�,k?B���լk�����N#��w�`���y�7o��4CK�jaE�T�av�Dx�����|�IЉ47���� �=M����fK��1�z�&j�V9����@`O E���H��J�ɑ��
��tʈ��7� ܥ�T�--l5HR�]jXS��H�%R����T��z�T�v5|�z�Ԥ%��T\O3#C��̵yb��v�JAm/�����x�9@H��r]�����,�h�|�clX��X*J�����X-��,��V=�.�h��Z��b��h����DZz<5�ⰵ3��T�S}i}�p02"�ŕkͿ]� `��5>x�hʕ����,n�+kFG��Q��IkcS��r�5��.R���SC��1�=5�d�G�I����\5�#e����~#R� 璉5��E3���w����gZC��ie	`������B��#�V�DZX$ �~�M����b/?�0�E;�7lL�VMܭs�����|6a%���ūq�y�s�S�8j��-k_�Je~�B$����W���x�M�8�P���>W��$:d�U�w�qt��I@ϥj>��#���@ϒgN޼�Na�������z=�����]��4����u�Z������C���6d^��"��)fB�^̚2���������)�o�(lH���F6$�cdA��D���ɮ��ٲm�\����<��3�ϟ�u�P^��p�;�*�/\�J���S��ǧ����Ϙ;�?r���<�l��ɓ��k������/��+��v�jEĒihJ��(��g[�5o���ͧ_?��8{�'�>`ф�$�Z�(�O����WCr<�8�g;���ĕ�Wٲ{7.\��������,fK��)5�k�7�o��|��+m�ԎSY}x7��\`��a����S��r��pi�\G+KGU�iw�d��BD_���pd��$����Rh�H��O�r-S\C8W���
��/��~���ϴ����w���>��o���F>ob3y��98�WR)σ�x.0t�z7���/���¹o�M�ڵ:���i�
�R�m4Ëz��+��y�.��,����TVn�
�e��.�Ur�Ig�_���M[H�i �8<�#�6����_�,oL%?[�Y�y�d狷���G�VF��U-�`�j��g�i�FK�5�Ȑ���qw���;���,ڴ���~c��u˳Z0#0��Ջ�Ґv�]�
o��{�*��j#�l{�;a������vֆg�{c�?�Q���u��U��.f	��[0.܅.k#z�0*;�v���pfI���K���d�5���!\�~���#w?�ѫ��~���W�j��'����;�z�7>���'8}A�{��En}�-k�ޢN�I�
TG_�H'��$��a8V�ƴ�	<Q��25���k�@ �.A]��v�kV���]י��1��rF/��e�}@_F�j�(6
�t������;a=�Gۄ_߿���Sp���"����?5Å_��`��0{��evMʲ�P��JKP�Py���Ep_2⃴�|:�
�TO��]��)�ϼb�����&���*n	�]��S��/���=�K��8��C���A��8���&,�x�[w?e��̞4��w+�gΤ��=��}�2x�TF��ǖ'9��F�O_e��������l1o�Nn�����o�zú]G8z��Z:�f8�Q~v�����̭�H�I\.��ÀI�����H�X5p���}	�6����ت@� ��<����+���S�5�a�d�������<�5f�
�Z�WM2p��[�8L�g�/`gP{6�es��=WZ(�$O蜈^�0Lb`�����XTk�}D]l�c&뭲�n�<{	F!��Yg`�\��$���Nۙ4k9�^=G�`�>��8�8����l43�g����l����l�@���%d
�K��ܤT�P���C�B�q���4�E%�Xlb�� O�
s��d�3+mh$�ښx?2C��K��q�:RE�\�h�cO;��S�lJM=�t��X�U�1S�0m�rts������z�l
̍������.HZ���a��S�&�T4�*��N'��Jz�gy���`��r��TUO��� ��2Qs�LM4��&8ؚc. def��������&�@Q_;�����1��|VC�JFgz3�V��yGG{��=G'k@3I-���^�B�Hu^j�����Ԁ� �ܤR��/�mnTՓg�O���bJE�P�-�嘵`{y�����r��&�J@�R��G��3����<��yʿ�9Y����~� ��>�'_�HEF�����d��h������R�Z�i1<U��4;2���L[{ͪW-״��P���G�"���څyQ�L�M���qv6d
 e:�1$<�	܎�͙���p�>@����g��c%�ʷݧ^<5�ȓ���$�A};�mM�"�����n�5���z
�u�#C���ly���À(ڸ	0�l�Du9V���x!�t���{���\?z�XkK��Z��*��dw/6͛��ΗOs��9~��[~��+�5(��O��	�ުX�e��Z�%?�ē{�9wr?�	����;�,��e����O0�_~ǿ�������_�����~ǻ��b���ה���'V���֮��F|����>�R�f�q�-�����hfH��>�۵@��㷟��WR�(�	�1{`jXK�ӣ�ԁ\
<�ٻho����Ϟ���g���O��z�V)�d(�6P�l&�dF��
>�u�ןƓO��ۯx��K��%�І�v����zxfԑwj�{gS�Yj�M'��^���<O���0Z���(#�H3%RnԒm���%4�S��\���O$׃c9/�s�/�c����\��
��4��c4���hD<��G�#8L�����3�0����c�_�Bc��3{�<s�{�ƹ��F�D��1�M3'�����8����}F�;:��z������[���iKi٪+e��	��!04��D���
���ȹ
�U	��_`O�P	䅆����bq'g��N͔Rjd��SDe�f��7���W2i�t�uƢ�fL�eX�|z�5�U~"`���5� O�KA^�*��S���A���y��1�)���N�e]���MnG�����G�{ ��#�6ި1W�ߌ���s���=�䙽ܸ}�k�nr��E��?�A��s9|��/^a��9u���q�������l9q��CaQ�ή::�@�;t�~r-Mp-\�S}�8G�N�dY'�y��5��Q���w�K�E_�����u���f�1nf~��y55�S=y
��E��-T o*��V��6-MG+��A�� ���e�O)(��6x����T�ߟ���<�}�]����?T
dgV۸sP��s��9�'֑�O�ϋ�[9���;-e׌�,�&'y�]��1������\�m*�W(����UbT|�
�%��l����*���.�QV^y4�8�'op��9��\����X0v!',d�Љ��1�Q#�1n�2��\���X�v'+�lc��c\�~��w��q�	z���i�7#C�md�΃��,�Ǵ�X�oA��C2�@^�6Ls֣�>�`i-x�@ϵFN�1vc+��J���04+A�X �,�C��.*4Gǆ�=�Eu�z��;��V2k+ɜ�1	h���EX{#�z�LҧbY����0�;�K1*��a�lt5g`�2�艚�;9�MX;l��a�_�eDcL�b��bܮ�${!�Q�H�"[2`.�5{а�2���L�.�ɔ�{�,�B|��SB��t4���d����[�g�E�Xcd�jCkV蛳\�L�*)�Z��h1m�Ja�T5\[y�-��Ζ.c�h��D^�^k������<=S�Լ<w�"��r���+�*��o��b螚L��!t����ÝXݙ�I�t�r�M�5u\��)��b%�'p�,oݥ"u42��J�ի��ej�z��0�S�zȩ�ZsFp�t[:}=�T���ߐW�NO*#=�N���Wi߉>�}S������S�Ī�ȱ�1X�
/$�g(��O��:W���y�٩ؓ6��i�ci#ki���
af��<3�b�B� X͆���dJ���nF�s3����C/;�|���s �͎D[�,�27#�Ƅ,Gk:�{3�֓s��<���r��RaZj �o`�^(8Ss�"��ޟ"��u�n\������f�-�\�#�-0��i`�|�X����K01�bp�JEV`�L�@E���H��P��fe+� mb}ãAѼ�����t:�
�5Xؒ�g�H�{�����S�y�r�-�;��\��S�>�SNg�[�r�Ȗ��|f��=�V�����Td.;N[�kֺ$�Y�@ﮂ;#7>5��΍7v�|����R�Ba�jZ�j�t/�à�յ/�Zv��N|R�	�մ�a5��I������o�n|/�����x�}=R���)�8N��Yt��uef��mՃ6�k�C`�ʺ���h1�
����_Fep!�.�[лM7>(�Ѩ�eyp󎴐{�e�E��%���r�l9�S�£��@����w�0\��mj�A�r��igN��4>��!��v���o~���M�LM��A���9�rO���U
|��.�҆��lC���۰-}J*hCm5��N�˂F�<;%��-���9u�R�>r�i�R@��\*]����)��!�P-�6�Lt6��kjVޙ&�r��+y�I�<���2D����)�[*�~������:S�șr��Z��V���0s����,�i"��fvT���%ǪTY�Y��ƅ:�6Z>(��'q|o�w���::��N4�L�|"�zW69�B���x�ҝ�nܕ��e{'��u<�d,S겯�������k���/��Çw�u��N�d޲U��7���PX\�R2�Ν;ҩ{gʛ�%�Ni�6�C��m�ݨ������צ�^%-ڴ�G��7�+��n���^��A��m��y���+����h]�o��7����yzj�ֳ�{�>w{��v�z��6d��^�PF�Ћ��a��w	T�D?�j�6O�Aۉq���I�����L���Ws��iN\:�9��t�/����3r?������s���#�Nq��-.^���Y�-��i�l\c`���y�/����K��z8/�����@��_���/9�^� �,�J�	�A���;�$��z�}��PY��6S7?a݄S\���7��|��S���#�#�Ѭ���ؙU��N����G����<-��޽������*����%���z�06��HA��Ϡ�!�U$����h�*N������8<�2��<f�7��=ʅ�mãB�w�7�/V�G��W9.,TaH�aoǵ�A�f��B��i�y^Q����=����a�I�ҟa�1v�x��̔�0vc�/`���,_��)�3b�d����C����5N|F�3�^ڎ��68E�@g��zu(ڂa�Ft�[�e�yy�0�Z�~�l�'��5DΫ'N��bh�^�P2�U�!O�4=���	��Uů�U�ATG���<5<�B2i��Za�Ө�����,e<������.m���(tIC�̞�U�t��`�8M��5��mHk�B�b-Pi���^�e�E/o>����&/�u-�j��XyF[o0n�t2�R�_��I��1��K��y��j���T�
�l�����߀gP%���B��ҮC�j��B�G���tY?Q�AR95�p�\#4�cty6�;��}&�������|����^5��	`r����fC��y��Դ2 �ژ[-��� �)�Q>�T�SkB�V���\���PR�_��>WY�~����aO����jk�25ɲ�T,J�"�o�9T���T><�:�Z��%�y�h�z��L��r��giD�����3j8[��fE��MC���ʐ����`xW�'��#ޕ��4�u����n�d�ڑ`cF��E�����-��YCwzű�=J �Bs��c`�Y���uTV��2TO�:kw�Y)�Zc����[
�f�����/��=���i��@��Z5#�ؚ�R5��L~[����rl�n�k5?��T�w|� 6�kAI�L�T�jxT���r�e`�:x��ړ�Z$��־\���#c�H���mKG�I~T����r�=��^U�@N9�p�6H�g�������=cn*��Ь!��<xc����'�&�c�@-+��s;w�|��"���'�Η��d9�'�d�4�j��H�FX#��4�|�v-jʵv}X[Ѐ6^�!�&͐T�ϔ�^�N�gi��D�=RC�C��s,!G�!��2Q��7�W�`2�ɛ4��R6���If�����j`/PbJ������	��kҙsEM�]�=�veBX
��*DZ�4>2MLɶ4���?�e����T֊ˍڳ�N}�88QdnA��-E&�J#��Ɲ2;O�̝ɶ�"���[
��,�)3w�����u�:k��{�V���,�)����20�0�X�����h=%Ϟ����oZ�V����V�=N�`OP]u�y*_��)�Sý��1��,]%���<�w��R��8z�-�e��o��leM+9�\S��/e���ĉ�I|m���QC�+=�hf���H)���v���x"��M�c�t���r^*�Ł�>4�ݵZ��Yo~��}���w������H������w�p��1v���Z�#�v���U�ݼ�ӻ�9�w7�֯e���?���gN�{�f6�\Ζ�غr-��o�Ў�ع�K}��U�iq��v��?�C�j��;���-i_o(�՚�y���x!OI��)��yu�,nu>]��k���D4]���<xy����+�9�S�t���W}Zv��փg9~��o>��ݧ\�yK��Μ`���8|D����Y����;�d��Ӵ`��*Bg��4=yU�5}�B��&��x�{��`Tr#�;���U��~�S5��Y�x��Cb�������y3v\cƶl�t���|����I��ms�� o�����̪��UX�O�S�!������!�I\]L1e=K[��ؼl���u�_p��Ƭz�c���.hõ�'Ϡ�����B!]弰XҜ���=�{�mF��R.K����	����;�{�"K׬�&��ٗQ}�1��dF����Ә8q>�-a����:�.=�ұ�(�v�ü{�t���0��Qn���M3��+@��w36�m�@R��k1�؈i�r��)U����8H+ö%:�
��"�-
�25�3��
*� OŮUqiUx3�ĮX$t�8R2oh9f+���(�ǯZWm~�� �2�P�gmb{��k,j.-���>�v�,�%V�Ͱk�E�r�c�a^����0*���Wq���4U`4��~����m�3j�T�<HO�������9C��d��<�ֆUz�,�e5�Z���<m*�����B
�Q�il�:N����*]jj'�����e���}���z��3D�e���t1����P��1�c	g��������I��é>1\^��#�8?$���b��&������ɨ�Uw�{��}�h�nL��>vZ��DSC���z��SZ�
�<i�)04��`��H�i,��J���T����O3�_�ro?�L�T<��+��}5�lc �e��I��I>+(R�f��p���5է��	��C>�4���u���l�`ːT{Fe�1�Б��,i�����n����m͖�,k�˜
i ��1�ȟ���4��N� gj:���b)���0���	(�5���3�9�<9w9'w�*�Z5)�a��d��um�V���U�[]9�E+��W�W�fJ�y]Z�_��s�/�f5ʵ���_��C��H͚��ڑ|�*�޽B�8U��%s���T=��N�����|n�`�Ήb��@����ƫ�$���n��u'_�9rW�ಙ������x(��=;�H��
t\�<���}�,@�U{��{qG@꾀�s���R1?6u�@�?{�>չ��>��!5g�-�1�r������,�<o�Iu�}ocK����^�h�� %Gߔ<3:��p�?�W1|�Λ�\���0@��D�ɶ�Ռ��j��#��P\]I�ȑ�u�������ܛ����r��D�^̋7�Rr��2$o�	xճu�� {�� )@ֿ�*���Y���jI<����o</YbE� }�4�2ts�d�5�k��η5y�&�Id�����؊�*��	�����bC#���UH9P[=k�.u���]���GGy�f�����SjeKS9o�Y�h�4�47�� �-��aJ�$�`-f�I�����y����|f��P)pU`&�sG��>YQ*PU.yM��\�9���c�H'M�5�r��9�9�d�/G�W��=5�l�g.�'0��y���&N �+�������4v,���X'���n�ܒ���4�Gf�<3�ɩ��>�#���0�_ρU�8�^ l�~Nm���[9�t��آ������a�Tv��˾ɋ89o��*�:v���l9�Mæ�o�B��[�����=�M#g�m�|����nC94q�La]vFz$�Zη[V-�{�L���@���_R�y*��@�γ+:oI���z��7�ߐ#���V OA�N�swa���Z;��y�����ǡ�a�KVc\�:�bk��[���^s�Uγ��Mv_�ξ���v���f��Kl>}�E�.�k��;`�"�} :C't�����bT�:�h�ca]��~�>�������$�}Æ�1ns�.7����=c���L�|I��m�.r/��y�z&�EDMmN��m�v�{8gFOp��f5��?����/!o��@^p�yO-#4�{<n	�&�bA�	�y�����c�{�ԍ���z�jZ��+��=�.K�.���G0�?�q�o��Jv�\�Ts?��
�1�0b2�g�t�������?y&�;�_�toݛ�F3z�Lz�O�.�i�c,�̢ߨ����:`�"
����%
CHy@�x�Źr?�ʷN���A�jt�+0L���=�	�u�H�k�����M):�\�̳�7IGϸ�@^��,<�9f	�m�֘'v�>�'�)�1��(��V��S���b�=}9�U-,��R1��z�U9��F�(h2��Leq�?�7�9����k�����`���^8��Ǧ�,��'� /�mMt�ev�ŀU�]s�.m��lbGJt}
K4ț����{�VA�j�����vK�Z��䉖��L������W�k�u�)4�w���n��[.�F�)8�2��'�}�����ʶ�Bd�HW)ܻ֨��OjsmQk/n���ٵy2+��s��l~6�/����Z<_�ç3��7!�K�R8�5��m���<�����0��žL(�eT��R��aK�`K���P�`Ɉ,gC���H�Q���V�� �@W���G *7 b���&�(����*��(�J�k�G��g{C2�ud8�Hqԑ�,��fH������T[Y�>Ė�Q�qbD�/���]/��Mr[U�ۑnq��/�!����9:����71��S�y2����qwTW��ql�@_�(6����L�Š�(�Ey��lI��9M�m����&��Kj�O�۶H��
��o,Pg���S����$/m����@�=�O��o�މ*�ZF�xp�#���x��)��Yk�0Ҭ�h�Do�Ԝ��*�w�Td���:��ڙہ1�Tȵ���w�ܪ�xEr����y�͗�a�xSs��	�ܒ����#+7����������&y���<��[-�k�ޜ�p䮏o����4����Y����]|*��g�"��6\{�'��Ȫ/ۦ�[��oF���户T�|�@T�,g� �oh����o.�-����9/�^�3��CO���@�xs'2�?����_iC�ffd�-y-��X������1��Ï��l��hE���ܯTcc�-�)p.�����L`ސ#3�M�H�w�X~k��?߻F�\�OzN���d�A ��H0�!]�;��E@Ֆ�4/\���$�otn��3��>���*�7"�ڊ2KJ��)32Ҥ��׷��������Jer/�,��g� ph�A^mȹ��ZR_`�����\bl"�(�"��70ЎQ����u6�|y3"�ɵ��"��x]�Հdz	h+XS��'�^haO�����e����o�1�֤��
�UJc�����_R��r��r?�$������1\ލ�R��,��"��z:���hjhA������ֹ�r_��ΞOM�yn�g��\�
f�s(7��9��4x6���e]�^li7�==ư�y_����a�|H�cmrD�}�{���5��[����ڰ���,��umY�ל5�-Y�ӂ�����me�֬�m���J�7`��0��+ڰ*�>�}�kMk+Z��Q7��~�1t���</I}z��$�����3R�������t+����؉A�~a���H]��t'��Rwbh��O|Cb���;�ݰ)��Dxa}&Ρ��C�~S��o���ԥF�I"�3�.p�-�#�S��sh��fr����(���T�Z����D���s�\Т}��|��K?e��GL�p�I��}��v���|�ϫ���C�a,uѢ��������_�S�i�}�2�Р��[^ߺ������WV�yp�;X��ϝ#4ȻU�3�sv�V����Aަ��X{�G/}%T�9=����J���Ũ�QLr�p��k�U={�D[���������M�b����'4�&uS��`�#L���1�2y�\&��� i}t�d}��a�̍�������y�<��vB��Is^l"/�N�.��ֵj^[�3[2C��3V��R]�f�䁅L��<�N9� ���ή@���E��c�jj�F߯�-��o+ik���u�:����1�j�9J�������Ϻ�94�2�g/r��9mN�ᣗز�4��.�9�	��ͱm�yxL#�`����8��ǥV?��F�Pg2����\]^�8t��gw���M����Fm�Vpz-��c��#��}��p�e�[��B����[c`�õ+�����Z%��G)�[%�:)��HKz|T:;��cyiF;F�V*�MR���3�z��ц�~���5�\��9r�i��i7s���=��}��%�S*����Gyϖ7��چ�Z[��V�lE���|���׫Jx>���s�u;��׳sy53���S�=6V�'�[�%��q��$�]���!�}�����[*�Y_�����)�ge�-ˋ��SˈY�L��cRMS��\�Pd��S�Դ�ԒI5,��d�I-O�iŔtf�3��9s,�Wd����;���k�z��a +*�U�ň�7ۖu�~�i��A��S�c�2$��2x85��3�x1/�/����Z|�������b�����֕�ӆ
�����Ԁ��6���z|��!�%�?����F��Kec�,�5N�CB5J=��mhco�2O�H�u^��G ��T�vc��� �py��bT����(�S���z��A�p���z%Ce��F�L���o"�g�6�1�b
)׷Ќ:�m(�s����o�S�W�����o6�ޣ��+"�8	Y\�J���i��&��6�<
���D>���?^z�i9�q䍅��;�Hޛ'������xa��5��oDp��:Dr�$�31���pӆi�0�䕾3/,���+�J��G=7��s卉7_�%q=*��1�Z<��^	�b�O���9�Ņ�2����.�&����H�FEGYV~�~Pª�'i�7H�_5�KY�&��TCoyƆ���jICE���ֹ�{2���. "r9d�[M�L�C�*�j���z��z��G-S+"���z�v���[�q��!0���P�Z/b��S����*�_�K�X0�����h���l�|����mdN��Y���
E%�����9�k�9���个'�Dʯ�zV��� R˪��H�c*�0�c�cP&���{&ʽQ�]#y�G���(��Qy���\�$$˹�!�<����89r�49�J���?�\9��˓��R��Eir>�Ʀ�\Eb��v:FJ��W�`.����B[;�~մ���
�ָz�MH2_��@�yE5����p�ƍC���!*��1�|�"�ubm�F��jh7�r���� ���e�L����ˁ��Z��mO�s�/EӉ����sȫ�|R���N�8�9E��=��n�lr��b��/�m�Ye[�Yf����7(�����o��[�*��h��]�ÿ O������T��VA��o8�������8K����Uֵ��0�ڂ~�r�a����]�Y�"o�u���x����Cg[K��d���H��;'y��nјم�/��3V@��Tx�R�T�Lt���Ƶd%6u�`*�+݄�_�t?���;��r�+ȫs��KU^���u���&��i�o|��C������cŨC�I��ni|�ǗQi�m��>)����sf�Xa�?D���B������q�C��gO�g0/�x��A���:|6e'flaq���q�����ا�;��?ã� ^��B�ra�B��r�0L?�~�Qs���8���<e������x�Oĥzs�����7w�m�	I(�Y�������#�3k�F��^#P��>�g�}�4z�C���H�h�kp��t�b����1�;v�kЯ�KH{�6O?uz�+D��I�K[/�Zt��%�D��C��!����ʃ���!����a
��ymXĴ�*�5�ͱ�m�-+�3�j�axK<��!-�%�J�<=��81v�2���7|��.�9��]�9-�7y�Z�B�c�.�k&�~3L"����a���,�p�ð/�s�@�bbl� �KD�n����S�R�S�7aZ�NLpve�TZ�� o���@��UR��j��+�,�2�0�o���n��
ڔVJA�ZZ��Z&��R���:��%���X+-�M��VO��UC�J��S�@O
�i�V�6����%M��Z'�-}2�:��zO�W����|��1o6����r^�.�Ŋb�^���뵥|��6�m���Me���vc���7�⏵��.������k���
~]S�w��x������e~?����9��0;������|3+�����fj���ʫ�i)�/&ej����y9.�J�y59��S2�jf_�N�y�|;?��d��B9��~^�Ϗi��)���D6�s��r{���ȋ��W����"�Y�*x����k��z����;���r��W������J~��o6�C���p��ȇ���sI��Ӯ�<_U��9���ə�U�7��&�ラ��NwW���k �I�뤁)���X�D}yn��!�ИP�6̰
�Ԝ�R�~���f�pG�(��Ft��jH6P*Lգ�Z*޽N�|�ß���Zɖ�ꛛk�O����*��8T�����r�m�j�ȣ�X�Ƨq.0����0��2UYb��s�}(OC���9��f�< }b�Ml���1�N��iA�oDgr98��!�l��ai�;��}`!+�İ$͟i�H��4�&�|�9��Y��S־\���m0Cy�ƫ�l'��$����<�!y%���i���iě�V<�ӑW�p�V#:	\*�p3���s�+�מ�<s
���,��&�L�g��E��qc5�,4�$5d�TQ��^���+S�����s������F)k ��mhB����[jY)A���Ί8�*eP'Z��σj5\���Z?'kV�F��$���<s'Rͬ�/e���t>�K���<�N�Ь��X�e�D���<?J|(��G�W��Qd�A|C�@�:R[��a�B��3��Hʳ;o�l��m�E���>�9�g'_m�\��}�@P����_�%�	-�k�+���$���EZ]VG֠�݃ww��\d�I��;���O(�n!���Q.P^ϧ���jK#!�)�B�j���5�R�Pm��=\��[�lb�Y&�	�Eh ��Ԃ�������ɼL�g��/�fFD)�uC�'r�������^ܗ{uU���Sw��8gd�	����ᖕ<�`��zs�ҟ��[ƾ�4�e�`����HM��"�k-yV��l�5i�_���IHSN�qDߝ�r�c�~��0�b��{�̼�m�����i�"�P���G���O))���p�7��	���Ӥ���<57Oϧ��^�*��A�I�jk	�e�G?}�6�^/[�l����gl��[գ��[ l�u��T���aX��[�3O�����8A��4B�.�
[撉A��G|�}�\|��î�2��-l�]�:5o�f٫��/�+=�����ߐ���6?� oڶK�[��#s;�=߻H����A��'O o��/�%/�=J��W�S\��C�6\��Ｘv�����'��&N,�ve�{��i�����ɤ����ŭ�pp���b���y�#W?���q����Uސ>�7��y��CB�0�ٍy�.t)4
w������ڼ3C;��{��}i���R-���f�6�C�z�H�ݎ��V�' �yH�a�g/���32��N� ~,VE;0-��W��SWa���i��Wc����j�R���6A2�d*�v85EgS_T&�'4� ��B@�(�o�3���*�%�񭰎n�mL3,�T�[S�"�c�Z@��67O�����L	.�LY��7�?���9z�5��s��1&�Z�s5y��m%��J ��&��V��u�9�nE�p*�kn�c*1��V�y,	E�0h�^���ANj^��lږ�}3�Ói�U�7�� &9y�@
��&�ӯ�Us��40��g�z�Y����yk� Ϛ)Q���:�U��'�f��=�廵sj�VA��zUΖ��S-~m+�:��4؋��ތ)�g{�\��ǃ�żY[�o65����׆J�g꫕��jm��^�l(�_������������S������@3�Ӕ?w4����P;8މw�Z	�Smx{�5�h���yw�!
0��/�'���6�[󇀒J��k"`�P~��7�~��?�7�}������|8Қ?���cm���s+>n����qsL
�����W����2�}�B�n],�Sr�uyw�	�7�\�҇#ͫt�%�l�o�Z�ۙ6�z�����Л�����)�9ۅ���/���|�HfG�hf6��Gz�ռ���ISwZ�Y�G�����V�f�[ e�|U����!�$���	�}��2��-�U���'�9N;�:�#�_*���W�����,XUT_{��c~]��fRjkM����>E���rpѤ,n��ώNdX���Ɗ�B� 6���	�K��f��p`j����*��6�͏�ޡ�,�6a|��lcgW��WV���90yG&-����,�ߟq��d`6��Ĥ���ׯ#G�����ul�3��}F���p�t�Fs�ljؑ���p��'kӛc����awvUv�p�VnҔ��r�u�uĩ�Yݼ;{�f�'�դ��t�]�v��h��&m9�e0w;�d�\�֟��2�ASzU6�iQ!-��h_^N��,�ӳAC��nO�Vh_����l�����?;t�\�>�mډQM;б�1�4cx�ތ�އn�[Ѻ�>�˛2�Ig�����iŠʖ,m�A��[-�q�mN��Κ�m^�!]�W2N��5d���fՄi\������x�\��_̙���0h2���`����7�哖�d�|捙ɬ���?n'�`�ة�=��3��h�"�M����+Y>k9�f.Ѵt�BO�˒���"V�Y��i�Y:u+��b�$�n�f�^͂�8�p	O���錕|1{3_������Y3��cӜ�l������N�k�v6����i�ؼ`�ɶ3Wk�Y�Y%y`�ʝlX��u�6�v�mݚ�Y<u1���iSڈ�u[үeG�6iD���9Ѫ7$�\nӋ����mF���U�#��;е����>��=��Yo��#�[V�<rP�纙��$��m �%ϟu�傕Wm}5]��G.���EpO���Na(��J��tE�]w��"���	�s�,GI�y�j�;$�o��>9��n+Ov	ln�tb� �V'�H�f��/�t��p���{5��p����y^]�����<ߡ��G��,c�@�F�ti������UI_M��ݬ��&E{ѥ�v9[�,ۍ[�N�r�`�6�؁Zp]h'���<B巃:�rLbF`�2ǒ�8�>V�s��SJ@�x�u�bX�]� _���x*t�^�q����U\@W����e�9��-�Yr���_c�旬z���m��9]3��&6�c~��� ϛ��ޜ7R ���3�S��O�S!�~���_�ȁ~}Y��c{�X;��͟g�Ѽr��M��+y6u#'g�ce�%[t��G����Kv���1������70h|[HW.0�8Fy'1�9+�}R��ݥ�U�Nҷ���c�>e��U8������P)����B���)�-���Q�}г�t�m\1�����] �Y��� �����p�cTzF@s�@�*��Vb�����씒����X�ֹ�A�(�С�? /�]M��5��)��ȫ����&�� �)�%6Q�5г���vXDw�$���:JFm�εרR&-X��7�x��6��]b��=~�9R@��
�y5�\��$\I@Od������w�H����7 �(9O��r�5�Y֟�s�qR�]G�ޠa�A�T'o�~L��	=Y(��j���Vxf�ַ`����ç��Y�#���V���Q��������[��S=y���*�,����)�|��kboG�@o�'F�"ȑ��>χ�s|h"���jC��m����uu�zu߬+ ,ȫͿ�7��#�:		М�gD'��G���@k+Y>ށ�g���A�`0<���z<�?����|�ח�7{��^�ODK7e�CD��Z�#�ݑ���7;����v79n���/��/��~GI-��'��{��R'��؀��8=P9��dO�h>]T�_�ԓsX=و�U��i�����T;~��ݙv�?۞:j�y�;�n����^r����u���ݵ�~9؄/�WpZ>��d��m4*���K#_;�lԼ,G�l�%P_G�e?c�+�O��0W*x��[��h��
�	36�z|J%�l3S���u�����D#�NE��f`JuSK�WO�o%ya�TP���y˷%X���Y&j����ZT�Z"�*�s �ܘv�܊��CroU)��7���
�����i�z�vT��_5��-2�{�9��
���|��[�>x��#g�|�O����[\�rC�J\1b(��`��Q\<v����p��#N�ȕKw���nƳ��y�l�-�����ۚ���� �-�����]�n;�:.:��w��'�:���G�rv�.��ëϸr�.��Һ]|�T��y6���C���/����ɓ߳�kg��ٽG�<��/r��)�:���Ϲp�����mg��ey.�ǦC��|�n<�ڑs�8q��~ůϿ��;\=v�'����{��s�'����5��x�?����]��}�~;r���_����~�9?�/$����9v�ow����+���"_�5�<x�'����K�~ȣ�ϸ�->{�%_����}��#�z�*�o��r��Un����3��w��}ʥ��9{����ک�ܽ�X����}���r��}��y��w�~�.�v����|��4�m>ɋ��x(�sl�qN�ƕC�yx�)/|��ұ\=r�3;�j:����K�/k��ж�\8r����st�I�l8����}��}���8��gw��ɥ{\:q���6���m|;}%?/������|�>�y�k��qb�e���+�6v.�FN��s�3J�yV�	���s��~|*xF3�qᶗ��墝��}9g��o�:�s�%��6>��Kg�|5���^U=�'�NY�sV�Q�G̽�c��N3����N~��d��3Ll�h"e��m�YhD����i�M�S-�>B�g+��Vx
�԰�Է�����Y��	���D���Rw�D/f&�A^�Z��5U�\�^�ZLJ�bX���uU#s1��)�!�����dN��p�܂S�5ؗ.št1����Qo��k�)چs����ۅ�L ��~t
��\@IK ����C���Qs�ʎ�W��lϢ_��@�%tM�c��4y�Ni�ˎ=a������k��fdk�wJ�o���އE.>U��^����@��{��?�E��?������~�@���}���:{�ر�;�/�k��.��lbx�Pɫ�[91q7+�-��۬>���g��ʗ_� �rQ-nc��ƍncV���3r��	A/OnL�6�b�ԍ�n���`�/7�x).��b�����:�I�Asy:G�=�cg]%�:c_l]S���#��	��a��Ǽ`-��;4�Ǧi����RW��5�t	K�������Ga��AB�̦A�p�u�,ga`�"����y:V^u1m�E�����U��y�qMj�cB;,#[`�R��S��>ۣ�-�#�.ӗn�闏���-�\�Ī�k8v�$���?^����z������&�=���~���*�s�x܋GbU)p��!����L]|�K�S�����MZ�g|��Lv�`����`Z�>Ls�c��%�m����z����6�!�n��/�Y�Nό���l�
s���@^&�����V��m��kW�v��LYil�r���yzK�VHŮ����1�܊b*"<�M=G#
m�h�ĸ��4bW� �OK�يZ<_�ϧkr�lM-�-��ղR�ZW��66�mxw@�� ��}Dj
�Nw���ּ=ގ?/��P{<>�?̀���ϒ�2�J?���_�^����i"���x#�~1]>��ë��f�l7���F���1�{3��_�q��핾�c)}7�?�� ����۩�|4�]��ϧ��lM�//⋕%�������Fy����9�y���w��ϵ�r=�0�)j�$�SPw��v�ݱv���1?�+�-���\�ow�f�E109�vN4�5�����}�51&�Ҕ75����C�X�`̈́���o�d#��yy�FU�HLm4t�2$��zN<��Ly���a�����''���Ƣ��<
H�u@?�j���F��Sn'R�;;?�]Cɑ�&�ܚRgg��M4㄁֜��秨,>���z��|�sW.Wr�����K=����Y�h�P�G�pE*���vиvc��ԥk^}�̧Qz!���!���a�4���SHۜ�6�^F)uk�f�)ܸ���Ӗ���%�ks'��{��<N��eJc>Ol��5��UJC^%W�y�<�i���f��0�#+�z�>ږ��k�洫SA���.k���2I�-�ˇ�^��p��c|v=z�ңa36-^�o����m��֨��k�'�Ѿ�.�s�q��_�Kc�\މ���|�+�1��9}��g��L�<��=�0�qOF5���}�ߠ-mrʴm�5�ʹ��|�ׅ�����O*:s���K1�c_\�����!��i�i��+����څgùZgsc+��K��R�%Ӭz�#j�&����'���K�Cet.ݓKi�&��b�����>I��O�Jf6�]|-�Y7	L��G�}jm:�ץmJmZ�Q�?���:��4��[u;q��9���b���OoLC��j�&�,�'�g�Y�Dg�$&�B�we�_
����Y�����J��+�
���b��-�p���+��M�qt�qf�]H���)j@?�ףK�2&����]�T�E�O�U��R*�^�.ͨ�oJ�F=�8h:��90Q�n�<�垓?�l��,��~�0�↜��ۮ�\���<[o.:r�9�*u���H�N��s�.�?t�ʛ��2va��#�m}9 @�Ǻ�o�w��'�L��(8�����ٝg��tC�sj��+�$��|I+P��#o�gkM�~F"�^'2�k��;:��/uq��^�tq30��+T���үB/KA�JmڕQV�=��9{��e;��*��Z/з�J�VcT��8�d�֣_�Y@N`Q�+����jC���f�[�Ot@ �֛�I OWGE�8!�w��9r�Yt.c�����dή/Xq����g�glt�[�-yc��/�i�ص�����2���������m��9y�Oޟ*(�ߐ�����_9������o���.��v�y�X�'��qf�V�_���7Y~�sN�e��7�X� ��y�n���&���`X~�jn� �.g�fꬆg?B�a�u
ܩT'��S��0Ls��Pk.���	�N��nx�6��3s�,��ecV�eH	���L�{�X2�b���\yHٛї�1LW����0J^�~�2j,�;�(�䅚��G_��;����b�,s�7�4L�43�:�4�4��6OA�� �Kb���`����Z�<�i�8��%������ꇗ���1�.�e���y�2vA%��=�p���L�ǵ�4Z>Dz§�8�kOƵt6��,�e�Yw$K6\g΢�`ei��~\7f�6'OA��ƽ�"�7�!P3�P���zVq��)U��&=��P�w�l�$��,$5��׌,�G��#�l����R�.70�\�(�\%e�� S�\�o�j3{&����ʆ|7+��x1 =�:�z$�iiF��=����U�ʎO�qzB2Wg�qu^��K��\�.)���2M_��䇭-�}o�Q`'�sZ*���4}8с?$}A���ݓQ��J��_3奚�og�V�ǻY�~͕h9��Z P�_�����Z��+��%��q&�*���@�/�Ɨl��������������<-���g������7�x�z"o?����yw�3o�5緽��mG9lo���~S>j'�N�����r�ӭ��6�=՚��6��M�vw�\_�oח�zE�g�ss|��kͲ:a�J���}l�ll�,K7�IK�P LQ��W5�~��=�����M�W�p�J���y��
��&�o0r�e Wt6���`�w(�t�\�H3�J)F`-X�ň���)�+��4O�?e��Xq=Z8h��4p&��Ssӑ&��smw�~s��br�=�����<6���5p�#�ŏt37J��RA�smi�ǁU�iհ��3��I�Ւ@ɻI��$I�kd����L���-6w�Ig��4X�3�X4}	��.0pO*��e�x�Ә�Y�x�Ք�&O��5�Nznd4�VQ+N�jIw�XF�Θ�p7r���_�eu����Ľ:]�"�c��]�A��E�������FE�<������k�k5_2�̒ty�g�%q+�	#�p/�6�,��(Ҟ��l(��&ןf�L�TN�K�S�1��+j[v��ee_�g������v�D��&K�m�ż�s�ڢ�O��p���c���K��0uO{�b``*�V>�y�+`�"{$(#S���si���iC���r>%4��]Cȳ��.�����u���H�X&�����kϐ�*N�(e��e�B�o0u\Y�ېo����x�}$�?���v�S4��>RN%{�p��Yt駹��U�v�Ԗ�J��l:�ȥYL���kҲzZ�$S�7�B+/�����ł�3)K*��؉ S+B��I9���|1d>�Y�O}��ۘŬ.jJ��'����L����5p%��Sk��5���W4�=����Ukw.��p�Б��^ܲ���c�6T{Y�<x�\�@�B����ygm�ݫw��[3�Q��q�v�s��G�9jN��:�j�7_����f�K
-����+��O /�/��Q��#��y-0�i!��@Oh���~@;�^ /����yS�%�NX(�\Xa����Щ:=U@N��q����Z/��JٲN�#��
�j	{��C�!�"�;��K��o� O/_ �� zE�4�pz�{
�j�R�c�=�~��O�8��H������9��=� o��/�1r?w�!�w���)C�Zv���+��Nz���!�����/����ym�v��V�/��倏�֊��1�'��ܕ��9m��b݌Sl=��e����K�-��c�3�]�2�(�-:��2%�W��Sn�v���HyF)�0��FKk�ͭ!7��Zm~�Q�R�
��^����p�����fNƪ��`��fa��ے-���N[�e5+���_s�1�f��4]�"t	�I���-�[����`��z�s�i���_�A��4�~����
���cݢ��B �>��֛g'�<��@�����6ֆk-��3f6����~|����پm7GO��S���e��^�Y���Vo.0�����F5�"��Ń�;׺S5+[k5\k)��Gv�1�<��k�b��L@�۷����Ō�u`��;S��eJ�~L�B@E�X'0��.���W�^�ߐ'��Gț���n�X[օ��Q�)�SC���-Y�o�|��ERѪ!�RQn20a�T�--diCSi`���(��~��T8�j֚���44$�łV�mY�������ɝ�<[^����ܜ���Y	ܚS���3y�(�����k��i[c~��D��	��l·y��� Յ���;�?��������q��:G�l���̔��6Gӯt*UЦҟ�~�i��"��b����w�}XÇ?W���"��9O��ϒr��￞����ˋ1��l4<�sx�������.z-�eg#~�֐߶5�wu���>��q���hC�?�������b^����ܙ���q��+��ã9�'���Y�$�������`����̵a�}��9�Ng�yf*֬r{2X*�snո]=��R�+�
�	Zh/�d�HSKB��K�f���܉[��\�Y��?����i�W�O��r|ol����@�1�Fz�q[��U!�T�'�~�Ӗ�饴��\b��=�R����*�*y��Z����QN>�O��b���g���v�P�L��+�b��)�
��)�-aߎ�7�@�krXu�L����c�ڴ���E4.H�c�\�����]Y4a4��M�m�S;�&%��,:��8Z���׻����g|��v����U�7���rt�"�����ׯ�?��4
K���-���i��|��gb�~dFD�:?������',nۚ�sfqn����ޝH�&/9�o_��g붸��PT=��}�1cH:�3�A}Vv����,�WT��$&u�Đ���ط'	�Dh��@+'���
�8m!武o�>T��t�hίZ��%��s�(_?�ͣ�в-~V�,�=��r�>��bc�ǟয়yq���\e�ֵ��ڎ��[2n`���E�9�h.�c�(��ō��ҤQ�V��[�+W1��4iBݜZԊ�A����kҖ����O��m�]��6y��((��X��Q�7�VO��Mٗ�={2i��Ŵ�9e�ƌf�!lۺ���:�'�vj�1�w�C��5u�C9�|5���d��,]���K��`�R6�\���Y�|)g��Ԗ�ԫ�MFh�'̣mF��,.av�>�n֚��f����?��M[�u��g�d�'=�է+u�s��s���
`*��s�\���i�ܳs皹�A�9� �%P�z����i�w�F�=;.:����� �}��R��O�SC�gl��ړ�������-�[xH��F�ɻ�Zޡ]6���w}��7���L��kAn�0
h�.P Ͽ
���[b��\ ��-4�S�y�}��o{٦�l�]Ht�C1���?m&fY1�Z"p�L��g��I�W��&�~ڊ*�S� O�B�@[�?��d_���U�ݢI?o��k̢����z��Z���� � %
�D��ʏ`X�@�0Q��y�?�*�7��b�.>��%G^�t�f�W��}?��໘��BA�N��y�pj��"n�?�<���	�����ʀp�b^nc�Ao_��^;E��!��5�x�pgם`���l^}�-'^h~�v_|����qn��k��
��R`w�S��@eҬn�`X ϸf�) 3�3H^�I?IR�2����0$��Η�����i�H��겕ﲶ�C���/�<~	&�+4xT�����d<�.IZ	sqs�E�B/i��2J�[y�=�$��4A߶R�2��B������)����d�_Q�4[�¶z�Z��,���VA�@�w	:�8�ve��S��t���72�*f/]MA��9��īC�l�bX�E��r�X$���O���5��g����rNa��>���v�c���8�{SPT��3��9v��"���ͬ6��b�y�e���Y
��y:͒vFd�? /B�RUO��ϧ��6��죌/6I�\*11c��5�<����@��-����H	dPv��Ri[Y�!�)��jX0�R��Ӑ��,���)����QI�ǹ	I�ϕ�IܜR��32x8;�ϗh�X߬,�ե���!?miƯ�:����=ە߯��ã���b4�χ������r��a���4��y���W���\-}��,>�K�Z �(�[���.��t��voU/����� @���wr��F�ӝ�{<�w6�������v��u���v���۝�y��qU�ގ��������;Jy��6?o���kK�bY>/��dn.�&�qfx,G�E���u ˛���ҟq�^�s������%�<�X���I��:Uӆy�Kr�%��6,�pe�O(W�k��z
EB�y��'��J��nlB�T�!m���[e��+7�	��<�-�^� #�[OG����B�H9��?�*�����!�TY@>����F��lG{�`��K�T=4)��d��+P��� h*�"c����f=�ǔ�u���Oa���fe�~���-5���%O׎/�𖓴��K�)�Yy�<}��ҠV:��dӣi!��	�U0gT?VΝ̹G��ΫFͤ<4��'�U��t�����;�o\e��a��ؑڵkS��}`�ʥ�<s������o�Ӷ~������wC}�����I#�$'���(�4���O:ѽuC:�l���Y�'���/�<�/%�鼺���kaE��@��!�n�G�6�l۔Q�:ѡ��Z1m�(�6�d�������� Z��T�)E^�7l�����d�@Q�zhZ��I�F����@ω�8z�(_�ĄN�X/�c�T���v� n޸ȸ%��>y8]��q�vT�oD�-�߯'k/��s���ѣY	5�|�$#۴׬��ˋ{��0j�[��A�
��i۰)�:t�{���$��38u� ���`[�N�̭�)�k�&������4��VT�H�F^	��[�U�	��ΡA�U�����N�CYr������<@�o���/����~e�մ�7��}�ӨcW�{1h݇a�@���Oiߨ5�)�����Yu�w`��Ґ|�왳hծ=]�Z�t�L��()oH��\z���;�Y�r.�!A��s�n᤹�����u�J�ɗ�V�\5vцj���i�)y׭�l|5+
����ey�i����~��#䝰�ᤥ��V�C�~i��f��+[L\�$����U�z{�䭳�g��/C�x�P?��э1
��.H@O`O߯� ^c��b��H�NV>�4�3���E~*Th/���-g�M��rnu�~O��Q�rL37hQ�Ls��i�I�2a���k�=l������k��EM9�T��Qsբz���BQ�t��E��{D���<epQՋ'��Q*����it�.b�����e���=�ǔ=�W,���A�(wL��*�;��:�py�=C9-� �p���)Ë�R������ū�90p ��Y*�
k[�z�j/>s
枴�D��x�t^���]wY��!K��c����#6�µ��]�y��/ݞ0;$ԫ� ��9k3F���$��(y%��k�`/ML����R���ŉ�����GN�r����vi=�5V`����Ř&-Նf��d�d��ę�
�՘�A�BIh�%�w� ~f�O�.���a�=�'�bQ-t��|<==�+ϩ���^X#jt�\ �:��@^3�,#�����Ԭku�-%�
4z��ܓ�O*�i�!t4�v��Ұ�'dW����y��Ļ�j��Pf6*���<�>�qM���w�h��ϔt,֑u��|���Zw��ჷ�*��w`(�����W��;�q6N��Ŝ6���b�6\��\��3g������N�F�f}��P�z+��U�
������39�},�jwf�K$���)+ܕiی�4�yZ<[#3%�c�Ƣ�)���3.�R;JiW#�AY�4�"�� '}��ߡ�Tt�T��A�tMp�O���G��y�Zǲ�{�%�b914�scb�29��3�x43���c�|^
�e�fi>o�iָ��oƟg:��U����t4<ǟ��>��gcग़O7I4^����VI���xY/����G��q��6�x����w��>|8/�y�\j%jg[�Ǒ&�=ؐ_v��ǭe����������\M�.O��)|��&߭���l���\���)���N5XѸ:s+"QL�� :&{�4ʅ"/+RmM�16"S߈�nn�r���ƅ�v�,��g���\�Xi��2/��'�0�:��	�7��b��� ����$�U�7�_������8r�B$0u�#���i*�MA����6��Ԛ�aI�0���N�����O���Y������P����T�
@Լ�D3��<ҍ��5������5^*�L�^ū�^���qY�R-��a	��`��;��"����D���\��]�Iޫ�vt
���Cw��U�u�@VL4풒蔟O�|�4k��%�0x�Y���2i𤅄�}�2��Z,�VN��R��R[��X��TнmGZ�l��a��w�$�[udx��,:� srcB�׾iQI�GԠF@uZe�2��9��Q�F.�sKhע=�V��o��tkԁ�W�1��p����TZ��sҭU�֮�kE�t�͸&�Ծ7�{�U��4o؂��2�m'�<��vӝ�X6q2�.�e��4+�O��|�&f2�eG�vꮁefz����ގ�ܘ������l�nt��W�W3��P�
*�,mJ���Tf�R��E|@()Q�d��Ұ~C�ϛC�&M��rv�Y�T�!\`~���'��Q�f.*�S�Y@YJ]*�ѫ�-ͳP+:���xZ4�d�I<�ۋI-��V��X�l�T�΄��'�0������)���y���}�N�S��t�oBӔ���z��m���@W��ʪw���4lӇ䜺���S��e��а'�
��]F��)L�C�Z�X;s����7i������<'�'����RP��p�H¼�i+�8q�j�H$�ʚ0i,�9�\y��3�P�8�inR��xr��v��<�;p7�|�l��kMW}�>J ���s�~K��S�O�M9a᧹N9�ܧX���Z��K@p��'�L<�a��� ����<�b�MK���'�&2����Bʰ��*�S�r��*0	��i`cL�[��j2	P�ρmd��R�v�1�/a�g�z-��˰Ȝ�]�"V␿���h��z+�y�f�sq.߀K����²b��6c]��F;�e��������]��X�oļ�@�ȼ�f�l���v,��Ĭ��Z�xۅ�|/�2���yy�G�5>���0P�Ujy]���{�Z����|��C�?b��,:��e��p;�	�=��% �o%���b�<�䝟6[�Mp��B�)ȫ�*����|�����.sx�VH+{����m9���k)�_;��HZ���s<��k��c�	��}̢�Yw�+V�xC�Yױo~Q�V.��%���b�d�iq�2�P]��kt� �(E(:e�h���*I�R��[5��:����0V]�I�HB�N�&��(c1��0Hh�u	q"��*)��%��d�"��LC;]����g��d�o�C�u��y�'O@OA�֓'�T� �ĶXD6Ħz�*ȋk�EDSLc�]���W�󮏞w)z��Xe�U�wB)���x�(�"�&�A��{�`�]�Y@9�����]�FTb��炞xT�£�T���2�D ���/9�ك��#�I\�t���ɵ�_0��h�ۺ2�ɇ�1�I�8V���ӗ
V
�{��'�3�� �o�ӷ`���? �V /�C=��y���<�:�{�,�* �F}6����<V�jĩ�3虖B�j�T�:�>ޝ���4�$��w#c� �"�W��1�Q�͂�lu����e�;�"]����\o���gv��
fe�@��
�@�0�����Xn�O���4NM���b�YV�76����y��5�p)��3]��B/�]���˽�T�Õ>p�/�e��s=5q���?/v�݅����E�v��tމ~?ӊ_O���C���p[~��ZF�׶�|����֗�je�-)���|͚���ۣ�<��έ	�\���!�ƁO��3����Ph�̆��+`hA}2�h�Ee57R�m��s���խM5�#�̌8y.ʧ��u�hfB_#C:Ȳ2�h,����}�h"��Bʆ}m����D��\�T8X11!���V��1��r���rn�xrIg�y����ŮU=y���$H��Ԗ��󉠳��~azz�aF���v��R����G,�Bk0�3H��P�����#�Ԇ�<CK-������7f�����L~�㻠�L��|F���Yȕ�
v����y+8ݺ?G��YB:����XIR�������s��N5�|�0q�$&4���$��i��[��E����5Iu�MgL��+��!�{���CVp�́^^���i�:E�%�:����`jJ����~D��F�{���T�Ր�P,)A�}�a�$���B�٨3�_�L`m�R��R+*�Đ0j�EQ� `�J��Z&	d��P��K�\�ڦ4&�7_��)��� (�49� 7��<���%�/�ڲ�u|
�b���LQ���LjԎm�{��䕼l7���9ռ+EA�D�ǓX��I%�O�%/,��r���I)DV�NAv	��Wr��u�
,��o*�n��a�l��É�{���O�ܿzGR�?[s��:�+�������B�eU�&�_gOB}��%0�k@K�Z'R�If�Hb�X��.��;S�������� b�}�����k ~!�8���F�{4Ѯ����"L�;^�x,5*j͚ٛ�/��TM�!NKN%�Z<q������1���
�jR蟁��;�����%�"y$�Ι`s{�?�\'sW ���=���kC���}��7켸n���wY�Zza＃�w��|����������}A��N3i�I>�n�������f��7r�B�!޿:��ɻo�V�D-࿁sMݲ1���ȷ��1�h$�c�*1򩇱w	��y���I���i@	faR7F6E?�)z!��XG�P�!��)��O�IT;L�f���x�ۆi�p�rFa�7�Zcq(��S�D�'�-�VE�R����l�X2��)xם�o�r�����f|�¥�^�+�a_g+�[�p��w��d7>M�S��Y��^%��)Z�<Ą՗��<�֜d��Sl�6�gr-�9��_�D's<@E��z�T���S�
ͩ���Kȓ��] ��?�՝k�>�u�l�ٰ�Ȏ���q�'�P���3+�V�brs����-7Yx�%��|��}��>�6]��]AW*��Bz����D�t�|��Z%W��&8JZK�MM�����8������K�&U
���%�)v�j�]��\ �UO� Z���)�R��*)�S`�� ���6�S�@O�� 5����}�:	�)��
��
E��,��7Wΐ��ZKɀ���kõ�Q���i�C|��<��F�6�b�j>�Ѻ�<]R�w��y���x�p�V]x�l[$0XW�6	����G)�sHi�{i_����$S��TZH:���p���_����]�;`�����,�?�)��,�纨�@f7��"y�[�l�԰� ���Yh��7���'�����N䭵Tû:Ϳ�r��QŲ�7c���Z�&��J~���ji��KO�U��b=��̸o:�Y�am�����j"�g �g#���4�w&�ي8[3<�!��Tw�#�Ñ4og��ܩ���u�P:gGҿ8��u��Z[��y��VgO�xvO�|�T���ƨ,��L-|�g�sy�8O��S�� ��.?m���׭�����l�t]#ފ�Xߐ�
ה������^�pS(�^V�WKx��H�-��3k�p����|n�/�҈<NH�p�vwKe{�t6v�ɪ6�,k�ȢƱ̮_��u�S���`�d�ѩ�/<�H��H�.#T`.ĝ� B�p�2��!�Ƅ�}L�2"�֘4s��N9��57 ^�Ր�� ����lmX/=1gcC�'���\���bk���fq)\=��<5"�]E+Xc�E�����S0��"i��r��ܬ�!�!��
���8.'0��M뵈�7�z�{�k�B��C
_�,fu`�r,�K��F��M"Y Q��R�R�e�).Wb��)�X�n�f	?G��W���ŕ�|?~)�*z�5��a��%�ӾQvjΰ�-ر>�ۗ3i`+��hİ>�9�+��6&�ӋV��<ouSJ�sO�w��vl�jfѥ��.%t)��g�toז��ҮMjtf�2o���-�j���	��ܷ����a��,����c�ѯ;�{u�o��tjVN��E��)o�Ž��V�/C�]=���0>��Yq�ɉ�Vb�b�H��<�HeZu�RH��Nb�N�&VdY;�"��bEv|0�9�����O��d9F��ar�x�����A��&��˂u<�<���Y,�Πc�<:6hŤ>�Y>u:��/b��e�<���g��n�"&�B���3�$���G�Rlэxb�ݮH��[���(ap�ƌ�ߊ�]�1�Kc�iD�v�hڼ�\W�ܼ�%���<_�j,���m�p*k$ж^!��e|�Lh]�Ȗ�nS��r��M�iY�)"_��u�����ܟ$�hiD�g�ѳG���n��2�o_�������ߣ�:�d��Бx�¤l捞M�%��)#�Dw/��BI&�݉/�����r������4(��$�K� �+�`3��2�Ё��a�p�涽7w�t*�Ə�~�ٗk6Zl��6�����j���������9#�wR�sR��] �m�UI�O	�a�R����д_�O���#з��W���)l2wc��;,��g���K����%��Z`l怱����0p���=U��<�KDR?J��^�T��"�	0ꌝ��uТY���љ�g37Y�X�uC_$�虸H�*�Ef��9Fi�-�ݓ�w���)�8LE�NqX8�a� r���E䖨��-	+�dl=j`�Uo�tb]$O��&>�q��ɭ�@j�8RK�QZ4�fɽ�'eA|7:'��w�@�Odh�l�V�fA��l���C2q�lV�����n�����`~���$ND�E�Y�^yj������?y�ܻ���cX��2i%��vӼ���W^Q�q⪹��yX�{;�`�����x�)3t��/�I��/�jp���9�y�86<�[�ø�T>��`T�����ĺ�F�J�bX������(�J&9+0�_�e�U��Q�Bs�b���쥘d/�(}&��1I��I�$ӕ�`�6�T���	&O�6k!���SwN�˰̚-�LC/q��2J�ί�d�6�������m1��^V�X$cd��(J2X��a!0XO3�����>���&�j>��+1m%�������e{�R���}40tHm�}N[iEtƢFs����o�ŭ���d\_�E�(���vx��z�\+'`W��@C� �xu8��o�>��=�?|��ϳ��u�4f2V2�L� 5��ܺ�Y�R�M��l�e����<�����
yۥੂ�L���Xy�@X��)��
��|��R!��uu2�a��=�\#Y�]�>)�tH��4/��0�4���.��[�,��35��N*�<w+����bO53#�N/WW�=<���I��/�\�6�"���D_2�5�+	p�YuW:&x�+͇A�����E�̨��z�X�:���;G��k�zTgo�Xm�P�$���C�89,��S9�/��}�8�?��29�+AӁO�4��Ö6��m�,h\����Y֬:��D3�aˢY���X)$B�F��hH�HoF�R?�O�5��P_��|=H�����'a��x����@�,�����ꂙ��RI��:�c뀏���-P�*��"
�
��p�&�ޒpK3�T�i��ݹ��K�J1����H������nn��
�;@�=�Ba�	`)kO^j��׌ܸ���[(�=��R��#�aױ6n\�F�m��O�"��g�Q��z5���i+���#��Q<w��79��ۂRkgm��q��,�4��B{��H�ƅ�l�Ή�>�.��<�<"y!Ǻ�͎�
���ʞ�	I!�Ӆ�ݛqh�J�|~�gO/���)�?�/.���|���_\g���}.M�`޸���,�GO��y�l�?�O�^��Ϟk������~��s���|���ܸr�Q]��àv4�>r��FF�l\���K�=~|)%������7��|��&7���������W�c{1�k_�噇�Xҽ~!7�n���]<���k7s����Ń�x~�8�No��t�W�`S}��t��9��/*��yV�����݃���"��{yx� �Nl_Ϲ-�ܬ���l�N�����-���N�'�������_��WO���~�U]�����Wܹw���F��Bf|"�wa`�V�	�Dڙ2�kc��9��o.���a>{r�7�N��W���g������3�n[Ĭ��E��.9�9���8Y8�?��ϯ�]�g�N�����>���'Gy��4��?��>](JNa�tm۝8GOͯ���y��}���	O�]����|��?|��/_?���|��SN��AzD8q�!,�<�ʚ�ے��F�uX5}�7�����۷����p~�&v����]��2t Q.��\Ȱ�#��V�G:C �Wun��sK���hs����:E�[�Y{ʲ�&�9���@�Y'oN;zqZ����}�|'l��y��4}�=`��^[�<kvX{kN�ט:�F�w����]� e�
I��ܩ�[5έ��7���T@��>
#����� ��J�a1c���b���%˒%Y��%˶�������L�c�N”ĉ�8�$�̙�d8�_k+��9�w�{�����kU�������,58Zkq���V�Gh1���m�8�9T�����v���_q���Ϋ��"��tpD/�+=�'� wYz��nr��l���A�(�K��sT��;�Y���D�r��~���+N�J4��T�C��dȡ�_+���\�Z�{�)���{dݾ���5s)���U�8�}(�ks���{�M�1���X2�>4��$�q7:����E�ߖ���;��K����
���?��×�2o�r������p�� ޮh���Z�l�|E+/��RB7��>������q���p��3,[q��S�R��*Y��k8HQ�.ʫ�SU���Ɲd�l �nٍ��鹇��{��ۊ�|-��E$֮�����֣˝��3-�X��������P���%����\*���`̛���g����u9��vc�\�[�,���߲��a�H軗����WT�]�*�֠+[��}��^��p�/�+����f�����W�H-��!g>ų���1=�Oi�k% �]Kq�"@�b܍`��},�Sd�p��{]q
k�'�����+M���뭥?��ol\�{�Q�gb^��-,�:���꽎���ژ�\��ۙ?q#���ϣGo����x��=._}��c�1�ϼ�t�˾�QZ��R9�jr\��i�/:'V\v�qU �s��s��/�M�pr咜㤏��=�5~�ǰ��A^gZ3-�a�DT���sN*��ɹV���n�L��db� Nm$��tliHff��Z_�>�����m�t�<L �&^���,��)R����
t�#B��	pw%�D��& L��@���d&C@(�NnT��MW%�И�����O�-7�^�v�5�%-�ޙ�t�'0�8��E	�(��D��Y
��cgxyc��2�[6�sb�A[Z�l��oNm�	��N֮Ր�F}A&չ��g&S�OV|�&9)	�eg���HVb�&���$D�a!\�EA��M-�c2wB^Lt8fy� ?|�}��`�����F���-=��g��>D�;L�u�2�J��L� R����X���`���bLf"9��-1w�ܵİT��2D�^]ZȒ#f�J9zN��K�NX�+
W�uR �Z���e����>����D^L,d��E�JqE��u��&?
��O	e��:��{�Ӯ�R������橵�uq��B _�\�~;{���C?� ���1�#��R��qSKjx��efW�ʽ��f0�R]ƚu��d�Ong��޿����p��>��u���2i�`2BC�Jٹf;���Nև�^]�#������_�������,@�-_�5��>'f��q��3b�8֭؀�C �Å��B/Yȋ����K��ڽ�<z�%>��-~�����o��s����W���s�=�����w��$ ?sD+_�w�?���������>�/x������O�� �߼ŧ��0eHo�}'ҽ�J�����Z���W/�߽ŷ߾��~�Ͼ�����X����_>��^�߼��#����-�1n>��X�ЛS&�z�R�9ĉGٴu뷮aӶUlڱ�u{v2q�ƎE��7������6���u���0�/߹ɗ�
���/�v������מ��[x�׸��:��ޅ��d[b�&5>��i0��?|���o~��<�C���#>�����M~������X:w:%�y�=r�i�f����~�x�?|�>��;��w���o�㷿��o���������f���DX,Td�o�f�|MN�H�~��S�u~��� ���_����|ˏ��W���/�������� )� OcX�n⍰>M��{/�<0Gi��n`�6����j`�y*v�#�p�yY��T*������k��7�s_* �����j�՝�pmV�]m�E$7�]�qS 񪼏+�]�r! D˵��T�2��C�&�@��Hk��P��qZTH��	�>	Cd�@.b�Bj5q���9�/K6A�x"CD��R�=�~�c�)e��QήZ�-T��J�A���N�d����iβT�"e�՛t���)QYw���,w-�OO=5�X6�~�8o3+�Yiˤ]�7�ŗ07�6�2�!�Q���1���#R�=�����᤟�ˁ�<mGҚ��èb�M(���2>��cs�6�A��mr>�Bⴀ�7�c8��í�;!�?���V򿄼(�S;�y?��{m��Ź�9ԥ�O�5~�5�^����0�;߭�/}ėsVs���+��<远����kO�Ή��Y�u3J�0 s��C�1��6z���1��ڈ&�B�ɏh�ړ�VR�Ą7b��b� 1����b"�1���[B�X0X�	�߁��x[����Bj�)��@K>�J����Y�1�/n��q0U�i�!^A#��m�&��7�s��oT3��^xƴi�J�]q���O��'�x�=������B��?�n��,���u](^G�HW�is��3��axf��>�q���5j"�ѓ	�[�O�\����<L�u��!n,	qȟ�C�t\S'��4��^8���Ќ9o Q�1��"�~1��Hhۄ�l�����q}�[5�=����3�q��C�y����"S[�33��3S�=w{k��˗}.n��g:��M�PA������UYw]�)� �U��Z*9+��@@'�ؙ���	[���wT�sB��q�.�!=���FQ,[�0�$�%��Y���B/v6���4�v��
�S�s�ݜI	�#+З$O��0H�QL����ĘPc#		�o�J��_k�
�&�g��҈M"5%�ĄTBC"�����FaN��ŔdP��C^bYq)���MH'?)S(���*�� œE��B|Hi�
�(LK�<7Oe�sc�ئ*�r�-,����ny��,���,�2r���&3-S�+�x9����L����+.&CΕ��MzN���!%S�KI"&!��ؤ8��	�L��L���u~>�،z����w*F\�M���!ѣ�5L��tȳ�)�`Eysҋ����,v�Vs:���&;W|-�v��%_wl1,����1hql�v'īN���EI?g��5�>�]�'�����5�9�^'�uO��Ѹ����;���Y��n����1ξ<!��5}4�h~[���*e?ե�2c��h�1�e��ݏ� ����)5X�b��EL��^�}�VP��u;P� �ؕPOoCm�&F`��c`���,Y8���j�b"I�����������u=Ƕ�GQ�yU%錟<���2j�d:�g��	��8����ӿ�@��{�&ecB��4�veδ�l^��hoo��"aa��ePR\FQ~�	��R[SE��F̰A���Sth5�x�γk�E`6�Ǖ���8�oO]�,�x��_��{o\�7o��[7�@~��g��aPc!�N��&��,�*/�C��r��.�[�Ջ���v^�{�w޼�kNq��n��!=ȗrwa�Jv�G��yי�@E'D��k'.9�0qB�fBc��Z	�'PY�U�9���2��ZÀ�R-��J�7����O����-\���#Ƿ�w�:��$`�����1az����(#�8�R,�YA@�5���'p��N�]+ ���Ƿr��.N��ȉ��9�o9����GaF�Ϧy/Ũ'����%�7��|�DV-��d�I�G1l��.���͛Y�z5={����Q�����ө�z�Z��$p�8�7�}�G�<�ÇW�R �����W���g�ql�:�Bqt�RF�8Ԙ<UV	X�*��#[�u�X��Uj�仾y�:�eo+���z�&������+z�.u�E������i�0��Zv��?�y�	���H.��p���5o����

�	c��W�b8��A�oWl�Z� f:�1L���_5n����L�.{H)!�u�T`(��X����&��|�T���ĉ~��T$v�P$�ɓl9��3�[9]�ʯ�+NM��\�U�8s]��EW�˺
Y�X*����
��G�)��I���k������ o#�D7��b���.&VF1P`��݅��q�;82] �>����8%Ω
}�;X�3�@ �]���D|"��7�σ���Y��^�?���mB>7,˦py�Q����&5&�m?��C��������qq�<����ք�|�����$6󡵚��n�'��y�Uv��LX/����S���S��`+ᠬ_��\K<3Eϕ�����p�I! ��]��U���R8�<�tu�R�f���DWG?Y���I��s �.F�q)NB͊�ݽ����.��&<R�M>�Q
�^Ρ����O���at����M�w�B�'M'��N(=@�����LO�<n;>r� 'f� ,R8չC�3�p��kx��N|�0"�	`5�T�.�������;k�SpJ�����c�T��8�����O��˗�_��^��x��px��]8���1kQ8�7�%�g��O@b+�̡���&�z	q=��������=��������3�}�6^|�~č�O2$���M�y��8����֬f��qA��Ug#ץp�n�3�:Yp^���T�+"W�^�o�?���M�4�;)FO�]+�Q��;!���x�b��|g�R�op��9�i�ލ�YV�ϖ:;���c���Q��3���<o'g�6�^\�(�`�[�� /!F��j����Λ81��q�$��I���ʤP�)S`,""�p{�i�dd�] pW�O���<��s�-P�Ov^.Y�Yں[i��'��C�x��)�>���,���|9_Zj"Iqv��S�X�SQ^BYY�l/$S�MNI$=!���8�XR��H��'51���t��<����������2��I�H!A��,�-E�E��)�3u�y�����E�ͪ�fy�i�jc��5+�O-5��4���f�`KYw�(k�-�{I]�iM�fH�La\�
�)/��?�!���T_��mjpp���E� �I��Ϻ��B��4���5���(�;�><-�W�R�`Oe�@��M�s�ʱER~�J�ަ���%N˳��\���f����c��R,�V�t�
h�Hy/T&J�J����\*J:_~(��KH��u��zL� t�^$�ƒ]�����|����eܨ�D�Z�	�Yuz�k�{��p�PJl	�:��d5t:ݖ������d&�h!�N�)��]kXRŠnM��]�3�_GTh������&P׽V��ګg+]�*�\)ci'5\ ?�LuJ6��*:W ڏL)�zua��l]ޟ=�Fp`�X�m�ʡ͓9�y�����q�]?�^e��]\(���?B�<�K�W�����X9�����w� M����q|�`.n���!M��x1P���Tq�t�&J��spH(��plaR����I�P�P�H�2Rl�J�ɀ�R�����ˬ�)��?�ms�ع`[�`��A��5�-"+'�d��^���A��L��I�
 y/�W���=�;��u���0c��d���,��O����ܳt<�5�#%�H��Y�LC�)NKx�M�KJ��F��~�
�76�����Y,B,ia��<v�L���D����c���l�0�����e�26mY���;׳w�\�k��L�P��Q>�D�wP�z�G0φg�08^��=mZ��7�Cx�5�W=�y�+��JBy�-�&vTe�xh��fվd��R�='x���m37Hn�rG �<�-�~K K�S?��r���Th*#��w# ���.
ĜQ-X>� ��g�C �DL��_v���ؗ:W#ݼ�(�Og"�T�_�v�}����k�M���dO=�S*Xw�؏|Gq�~!���9x�+�I-* ,�PI���[�]O%u*d���z� Mz��_xb�H�<��n&&��9�5�Y�7�8�X!<�ߗog����w��$�x��qW�\M��wz^�粼��>a�ͣ�X�yK���z;�c��+�$�8�?��j���)�S����G�ʆ��q��o �����o�쵗�0c.G���s�N�ᩩk��������{>����Ͼ�s���LE;7Sj��6����器j��%pZ>�~!�bt��_)еP��$!�ᢔ���Q��ZD���1;��O�|�'W���8��G>�TВ ��z
�#J�mY�$A'y�/���A���x�XD1)18:jL/b	s��Κ(�,-����[D��wx��{8��/bQ� B��#��q������^8���98���A��|�3�1
���8�L�%E��g
�)ȋ��K��r��V��ڍ��;���'p�$ޓn��q��M8d��)~���N��Ƶ�f�ǚ1{�<��8J�@�CLo-�J|�r"h��٣7x���9~�^~�S.���p[�S�9]ޟy�܌Y��/L*�E�'=B������\r��T��R1/;zi�?��;��? O�5S�w�;PK�vH��1���M΋a�(�z[I9��9:������ʪ.r��椙��
>T�0/��nR��x���`�^�,�@��D��ـ�%/��C���(2�X�RV�C�@R��"
��R�	�
#*!�5{r��id�g�_ZH�@YNa�ϭg
�ӓI(|,
�� �e��C��/)�ȨP�u)/���@�,չ���D�EE�NBD$i��))d&'k�WT�Gn�\?+���,�;�[�Dulbr�)	rOzi�Z�mx��g���p�@/B@#*Ă�������Y�ڨ1������M�(.���57�Ɂ�΋�}K<��/��Tc-ϊ\�.�0&�BV]�!R�dY/��X��[��5�3E	�%���@޳�8^�����<��s?�k�~h7��)�V�������	�t�qB��y^�Ǐ�q|+�v8:I��)�#Iʫr�]��Z+B�{�_�K@0��1W�(����I�P�D�x��z6�{�����,_��5;7�e�v����Y�4��b6j?Bg"1�B��T�K1j,h������b4��7P�Aiq�ą�l"�q[��
\TA� BJ@���@�6AC���Ȕ��X�r�FO`Đ1�Z������"׷�*�`"[�'��F���t�7S�t���)��>�S�G���Ԧ�^=�#kFrb�hNo������-S�.�!K��V��
��u�w�����-�9�~�����!�ZݏKZ9��K�7j��ĉNwӑk��f �$%`�3�B�)(����c�2k��/�Kk[3�R���QT��&�P�f�T�nR.�����5�ط�G渀���#E�sre�-�ͱe��ۗ��(-D��׋hq`���K�f�:N-���y}�+��9�?�fߊal�ًˆqu�,���4���g���g��ia��c*����kX��KV�e�],^����z`�7u~1�9��7�nR��](��޻�9�Z�6��Û=��c0�Of��gBc1#kr�g&%8�8����Vgf{X���k����W$o��s�7���kH�%S�����Ѻg��4�@�
����L`��Z�=C���y����2V\������"O*�{R�Ӿr���0p^ �_${d���(�9��`��&�`�j���(v~���!]}�.�t6P�h� @���D���B���*8y�l�D�K�KT-��R&]D�;[�2����X%���z�ā����I����\/]���&��K)PI� n�Pz:�C ])�#�Lv�e���J�u����)�r�z�Ӿ�N2�W�!�6y�]Ի�qQ ���ۧ}ô�b�[��oDL1��m鄼/�2�Kb	��R�S�ќ6�j��RG��Y �ޒ';�����?������޺���_���A|z�"/O]�;�4>ҧ�J�d�?ǋ�o�����<a�۸޶��&�Bd7N�GjӨ�	��rճ���e�!���%W�{ ���z1Ѝ��V
@��Y��y�I�ʭ��PK0qq1bH�ILK'>9�؄,������HB�x����$�a���\Ajv6s
�H|ܭZ���܇
j���us�Y`�E�A�y��?�7W1t�.�8:;�$@�)���,����I��,�����5{L5�S��eN�e8��p���%~$�	pN�.�6K�n�v��8�N��k�T�g�T���{���~'��8�C�Z��8���x�M�3v�6F�?�/�ԑd5��e�b�/�!��6#�l�6��!��'.�7z�Kn��9���:Ʋ8H*�1��Rh�I�?�a�T���\t5���q^��y�s�>s�\czQ ��|�����{yj\�y1��]��
bGZ��ݵ+�q�zy*��u7_�(0��]v��	w?-�V�7���$���K����3���XcdW�(�V�04̓R_g"�[
���Wx]�8==�za�'2D<� /��.�K��8{y�	T��Rӭ�n�E{��ek e�� 6�.�(�CB��R�-222��ʢD�օb1P9�9��f���NvZE��yr��R��� ;���8��	��&i�@�)�Σ$7���9&_kM�J�=;�d1I���)�I�
䥥��=��C��_HAA�,�5��OJ�K�z��u�j]�!V@T�� �^�N	���t���(gHuwg�Vժ�ƺ8i�1:��%Eu��o�8�1��W�.ʷ�$�T��Ӣ�f˶d��*�6�60��(oȾw��O-yvG'ٿ��ےy�%��~\�~�E����ī���a�8$J��y���婍�k���_��ݰD��$�UJ%O��.���.a�&+I�M�<��x����%x{��D���6�DMI��ev��3�m�� X� z~e�VWh��	q�zb�-#1f3�n�ڳgz-�/ o!�LQf�yZ9=d�̣��Z@ҌM�ن�lz�1w�(�"�דP_BM<�V׬Z��EK�ݫeŕ�mݸ���*l�f€�
���3��wR�������\�>Z�l(6� ���"�N�Ҧ�<�c8g7�g�d���#\�xWG�����)��2���hrfS��_����X���tT-yF-��j�4��i�Ku�ZB#HHɤ��`��^���I�) $�����P��L�����%�NV3���sp� n�'����U�8����kzsjc��k���F��i�5W O�q���6A���P�)`��:���!���ڡ�Z܇}+�r��K�qa�hV��Y���4������:���R%�(�,��f�m� �r���XFRB�k���i�O�Yꟗ/iR�SD?&I9[T���X)�7{@7f�a�:f��`^��涕2�{]�M����
4jvKu��=}ǒƯ"r�$(����y���*��E��,w�瀯��*�Rx N�+�8<���*$JwıBl�^�@�Y���jO��T��&
��=$��u_+7=-\8<��b9�]k�q`�8��Ll�r�S��V�u�,=1�ş�b;�
��r�g��?����� u����w�N���ًn�_��_(�U���=Z>l�I)� 2�����&'4���r"Ɋ�'��LfR����DR�RIOL��=�(!2V5�8&QTi���B/sU��RG	��Ų18��j�TD����Oׅh�w�+T�K�*+��ջ~ѷ3��;Aw�'�<
��Z�~eI���d����i�<#�rA��+rNՒ�p��� �?!�1��o!O���گ�̵E٘$�Z}�<~�ק��c1������1��V�l�<L=̇;�py�z�����n�PD�B�9��QK�	,���/��~Q���-p�����P�c��M]T:ձ�t�-$ݞKh\&ƤL9�
K.,ƔWHPz.��%U(�zDD�&��cH� $5K|2�1	��l�DǕ��ZM���@��}}�����ჳT4'Q\���ȝ��spU⤁��53G�5��������(\�	R]�1�D��ҙy�+�Jp�l�1z�sN�y�3;/J���q�C�H�$R��1���`W�
��w3e�<����7O�d�����ށ1yi5�H�[���	HDl���#K�K��Vn^��������}+
����&��	��j��)�"'��#睃48?�b�Z�.JE?/�AA���Y�dg䝩��{��Ʃ�q�Uq�d��<7��-
�['H8��k`_�f�N�ˢ�y��{���;��9>8���S8ޞ̬� j� |G��y�4w�_`\��5țP�7!f?�5/6�&�� �,�e!)1���d��r))�!?/���4��R����*�L��рO�zyy9�sJĩ1t��m9�t),'?�@@�D �T�)&1J�-Z@-6E��tQ<�ؾ�tr��R�4Q�Q�SИ�(�'.Q�4�xY*�KHpK&#=�S���0��l����99I[�%����BmX���yzh���A�
�����f4�E|��ٲI�Ndy����������M����Uʾ�A|T���=�կʁ�ο�B'�M�L�謺m�D낹%����m1�Lq�Jy҂!�<��(����$���x�O��i9�m9�Kn���tH*��cW�+�Xj�"#�=x*2���X�����r�E�1��P�5���Y��g� �Ty�F}���NNdJNB�db|��Az+��qb`���&d�s�^��>���ٸn=��'[7q.T�q��gWg7*�\�\�&7/�h<+z*cEGk+͵���ja@G_�v�	 E���)���v��C���j���n�f�R)�:i2˗�`��iL;�a�Fhe-�N�@Y���<9N��j%�h�շ�'�����!\�8��ri��N���i(�v�,;�c��;h����U��=J��c��]N�oӀ�얾�R�ɍ�W=8��/s[���l�����z/r�=Ix����3X��ka�2��sih�EbV:I��#H'�,��@s$3#��d�b�%��Qv�t�s|�`����m#8����6�ouO��!RǑ���Z�He��v��Z�� N����'�yQ9[ײoU���e�JY��ˁU�س���fǸ&��>4��Id!�ȯ��4�=݉I��.`�OTt��R�b�HI�����Iʕ��,����Hz����Z��"B��ޝY�e,Xɚ�,R����X3��5#�Y;���-](�w�/��1��H��k��ZK�{����ѵ�V�YU}�)2Y��
���9^����>�3 ����9��w窀�j'?&�~�+ev����R�ODq�?�'�v?�g�z@O��n\��V�N���0��j��FwO�y�����V�u��v��&c�q�f���Z��d� ��r��b��Ŏ(P�[�U�Q�،<ٮr$�Sh�&9�r��%��1!ȥť��NJBI��$�ĥ���G���Hq��	+(�*���*�rpV�&Q��t��������|:�ӽ�����d���qY̱g�K���C�|�g��w?��;&w�'��uO��r����~��q����ԫ.[;o����9�w�q| ��W�$�4'�}��xQ���X�¸h� ��-�:3^��@�
���m������{~���/]��9��4�O�\���xMn�cK:���Gx.���L�����%��r���s4����yc�&��X����lm���.������,�&:�n��ڴ���j*�[���޵��J�2J��*�W<#��
%5XJ��`��=�È����_(-�>+���mKs[)�X|���nL��UF��%J����-$�Ps����[��2w'g�%�A��
�&FCA^�� )�JԬ�)��B�:�`��URP����
\���`i�������D�4\#��>	�Љ8DM���9%.�9e���ӗ����<��9I�)�p�X�K�t9�p������6���I�v_��
���&�`$�5c��bc&�[�r��sZ7�3�_eq��He;�7s@�� m�JEs���q�`-��5Y^r	�O�sr��1���J�
yj�������wR@����v��ξ��cʻqz�J�Z�����1z{�@������yܞ���!��#�a�ޔ���Ƙ�5O�W�SЃ���:��q�Z��)����f5�2!&.���h�S��s��*��L�$7'C�>�ͪ�[U�gZ���P��7%��-G�O��zWT���e��](�I�("mʓ�LI#A�TrT��x��&�i�efi�|x��bd#�DG	�EŊ�	��&A`/)��$h�|�)�����ň�!ǈ�cc�.`��%�U�'��$�����Yʺ�;g)�ʩ�st��$�$�?IʿR���d�h�d�O0{�k�x�ݪ�
��Z��)O��F�{g�Y��+���T~�1p�9����)H{�];G�
�p�A���к�/	L^�s���j���R��!��� m|R��k�5^O���޶d�)�����Ie+�����孂��U�'%�|[7��[x����{��������sj�(��;iUZ��hy7^d�q��e֬�Ė5��v����� O�N4�Y��q���&���^�O9�&��ؐ��K�ߧ���Z*+����@�8�� bLzD�0C�橢b�o�Mr��j���K�8)!a�TWW3o�<Z�Z48Tc/������L��t朽���ռY���RF�ӳ�=�[;�pu�`��c����M���l Z*8\ڕ����dv5�������#9���&g7����A��4@�}v}o,����&�ԥ�99��<*����zvd�h B��!8���*&L�����p	������{R��1�f�t�7�G�ۺ��G���6�����=9�f ��sxYo�L���\/�����{�`t���������ae;�����%��^R��]k:�Ъ>\ї˚���x%���2��?��r!)���X�^ƅ	������6v<3��g�9T4����A� 3��y��X>�9��彘.0^m�fRc>3z0������1���S��{J;맵�zJ��=M�,�a\.ײ+����=C�6��M���	��Mb���^�ԉ#Ъb��/g���s_=`�Қ	��/�'pw�+�K>�L�������fW_�����E�����g����	�t7񤳉sn6�9�h�����IIT�<����jo#;�l���#�ut��T0�Mr�1�M��C�+6�M�z������S��M���J��<wyr5��t���#�ȰŐ`�a�!$$sXƈ4�t�t�2�M��'5��B�J�),�'�?q����~�rM
�b(ȧ�O�3�CF��da֯̒�}��#�>���ݭ�]�(L�Ҳ�$����`c�.�3b�
�=!pw���3�3�@�`�d�K���h����b}�A�u](�B���xj�	�~	x���)Z8���o�{�K��#��'����+<�`1o��󥽈׆/䳥�x��w�8�&?�o?���E싓�WՇ;�9�s*��F��a�j���X�����9|8DzA����J|����q�R�_yQ���Ft~��}��GdM/�+���ƺc�y
_��k=8p���'�s��eʪ��츚��
��#,)�^6t�H)q�Z�1�xH}ܚ�,� �QD�rx������R/�O��M
c���W(�R魹�q��[L9�	u8��`荣m��#q��{�h�����9���1q9.��:�I��L]�O�r�Sk� �!yA��-�Ko��b�Md�R�|��x���?�%�HL��>��#�vq��8s�<g�e�5��b���Gt�ì
=���8&�Q������.��yI P���l���@�	1ڝ��)F�syJ��ϐ�c{F�B��x!����FN�w��G�R��*��;Ti[n����[8�j7�����fAm2�����u<�T���hC-7'�$WO?�9��Dե��N����r��M}?LA>D���W�Od�{\81	��'D��-K���x��3S5���ːe��Od����
f��&Z�I�p%���|5sV<E5뱳��PkeKo3::Fd'���ݰ��I�'%j����kU�ldx���O%`CX�]�n��j�H����$^`NM ����mф��i�� �����<]]��
??��)�S�"e\uݚVTN����!&�4-Џ&�7#����Y~�u�S]��,�r��̙�D���%C�zG��i-y*�~7?m������ƾ��7j��low�Q<�����:��!��B�s��\�)Y�f��Zh�g�����<�ֽ�b���$�vd.����zto��H��'1�|%��">��?�+��"�I(�AX:�Gf�0(�w�9��X� q�\�1
$�T�Ы�7#u��9�� g��޻�I�|��Ɩ~Y����,/��'�ŝ(��~~����`�{T�E�84�T�����t���,�غ��l�:�o�D]4�nlfm�ƌ3غu+7���;���,[�@�.uqDp������l8Wv0ͦgic�7���\���E�K�����c(W���2^�*�%-��҅9K�Ӹ�f0�����~��o̅���V����pdIG����*���|�2������=�?�D�g*�j'%5��-,Y����jK��m�	<��X�R��m#��{��˯��fZ.���8�Z~oh�����Y՟�+0�����^���yS��#�-,�?���?2�i�e{L0k��qi9����X�ĞU��_�ʱ�}��Y������/coZ<_��ش�Afm���l�]ʺ�e{n�Q�L�IUsO[��z�FM�����81NLM��@�[�#9U؃�/�O��d�f֌�g��V6Ohe��>����Y��4{ �z�3�����8n��y-4����x�7�7Eg�I�K]zE��G���'��9oe�j#��U9N�U1�4����^���؁�N��֮��[��/��_.5�Y��uq�T˔��nV.x��E�wH�T��e:ڽ�����<� �y���cd����A�u�g�s �]��g�� �@���t7P�W�K�蝙���Jzt�Kr�R7���Ќ��Y���m���&���OD
^y�y��8'd�Y�[~�-�*j1to�T�TՄ��MsU�cZ��Cxe}�VJ�82�k7gs���M������!#4c'Τ�u0eI��4ư,*��a�Ӈr5 T�h_���ߗu�a<���Hꨊ���1���|fN��{����R�M���-����Sy���Ғ�?�<w��_��O�����O��ōk8�ԕ��Cx��i�����\>�,������$w���V�Sy��j�.޼�g�gGHC9��	Sk� .I*ajN7����q��1v����j'�w��S�h���֏��l��15$��0�}!���������2���p��^��/s�~a=ƕP30��E�5�Rۿ�7����c9�d;e�"#1����KA�O�3"gc8��(B�	�U
��x�⭺{z��꡵�=�Z�T�E|�&FP�t5���[N+��-;���^���V �N�6��"*�^h�H����)j"�8�/�)q.i�5qK]�[�
\�d[�\��r6���0|�b-�Lh������k4�di���Fl�0�k��\Equ;7n���_e���l�MՒʫ	�R�Q�i�ߝ�~k�t4�"NA�w�q��_���1x�ҙ�V��=yj̝����R�sj�1i�@�H���̓btψ�y\�	O��xq�Y��$����>�dz�H�rc|e/ol෧[��@5���7����f�Hd~�ݼ���'\�"@�!P ��銿����Q��S`/0�� �z�7�� B"�DDZ�G��IRL4�	qZ��t�71�jfnRl8)q�'�5Q�62U�nr�6+��$W�A���2�{7>6N����0m|�<5�/5=�$�G��S�oJ�ڪ��uɅ�1�!��"�������kK58>>^�[�ΫD�V�D�S�������b婼�
��xWy��cTդ5F-�C�j�s��b���(���v�o��e)�:�xF�vQ�ŉ�8S3�C\=�:��b��@}�Q�v}Z�̳�VE�q�ҺkUwd��S��U��j�;'��7_)cZ��y1Xj���.׽*��c�lKb�Kg>�Lo-5[��,uw��sqI\X~24��"��#���-���h<��S�Y܎���n	4>����TΚ��aK�����,�=܈A��w�Ap`1�jʫ�L�"(�D��;[ M��cdgkK�܇��h�ذ�74��^-=��֨�ި�C��Q%� 0f��`��hcUr&��`��-�D�
�ɬ���fmNbb"+V,����6X�b=V.�=79�M����΢�$��<X�Q�ͭ#�������ry��r�}Y���VYnP�%����'r�]�kC,/�^���Ʋ�l����-m[�ę�휓cU���Z��.����Z��d3�nfL��i�,������&) �H9[P0�	iLC9}�<J���(zB����a�~T�#��Ɛ�H�ڤ|�q�V+ۆ���8��G��	��_Vώ���Wͮ�5���,�ٍ��I�|ߕw*��ƘP3��oiw�ϭ�������\��ٹ���k�8( ��+�s8X������}������h��Ö"�?��{��p�Ff,X�ęK(�V�ILRp�:�*D���J�) ^��b�`���<�'[&�fۄ>l��Ω�1s['df�"�����h���������ڬY5S��9�W��<��N`ǃc�%�.D�s-$��/�<��2Z���)�{���U��go@K�L�|CL�C���b����G�%�`.9s���i'3��l�}�Y��kd���n� ����;��X�cf���y�����P�o�8O���� C�3�ѝɍR�BG~W*�b��2'Htu����hc����#��KN�->W���Z�F!��e�K��V�b��! ׀������k8!}	o��G,M0�j������y�Չ��` ��n��WGq��4f��"������ͧy�r�L��y#�3�'Z٘���������*�v��x���aܩ!'��ɼkL�S
��J �7u�����2�S�$	��U�
�h���߅�T���=��C~��7~��[<�n%�rjyg�"�z�>w�o�QI��m�I[�r�S��O$�iӷ_-k�<5q1�sx��Q1(o`G�a,9���'R>t8q�:mj��g(�m�jl���G���uXe��:��7a=���= K�PRGL�f�Pf��'�7���5�2*��^�LYޗ�;'2r�0��VQ�ʼ�I|��x���FyC2��b,���蝥Px�d�,��[D~"ޖp�-a���hԲx;{i]��y�Nub�t��C�����J�)�	�Ȯ8�w�5�w[n��8zj �hj���,��$��O���Ǹ�8$����[)��Pd�֝�4��yx�L' }���8��!j ������'������V���RK]�qܿ�&�caV[�P�w��T�#&λ�pQ�0%\-?�Ew���_v1
����9�v�O�wQ ��yy*��q�@��w�)�8�8���$.{�קf�p�ٟ�r���A��p"2�K}�2%��|��bI���o^$�f��ў��d����=���f>[]ə�P����f�ܴۜ�u:�tWWm2���~^.����ӹ`���^t����`bB�I!] +;1V3��>>�J�=��HQ�L�	'�NBL�&�Q��D�iK��
���I�=���(Mb�"e?���pm�|����Tݩ1�"��]@S����*��z?�ȩ.�`�[��6�?F�Q�ةV¸Xy���j��>��Iy�2��Y���U�E��)�%䩙�j�~����
� '�ەR�}�����N8xrM����8���)Pf��
�TZ�q>l��q�[�)'O	�=Ke�5^>����U&�T1�j�J�S���N9�<:˙�Oy�	�:xky:
H]4%2��_k��vrq��Y��d��7��]� ۦ���T��&��XT�T��lqj�ɽ�����7�͟�^:�]ܴY��@�
ҙ1s
���0W���e�%Tu��_�+�`�R��1D_[�x��H�^�_ :� <z��W3u�X�z5PV�ϸ1ô���fԑn����o.��(���}c!"TS� �WU�X�C����{�l!/'�${��� ��� eʽt�\+��J���U��6Z뒽�a ׶� ��F|\�2���pc� .�F�_�ߐo3�ˁ�n�v�����mh��65�������!Z��eM�^����\��TM�I���b6��᪍�K��!6,���\�f�ZLG��6�I�f��S�� �>��yjq�tĈ�&ˬبA��cKk9��'W4�w~-�'ua�26
�m�ǝ�Lވ��OgWp"}<�h
1�nd9��`��Zv/l�В6�XГC+�پ�Y r�'����G�1�d_��v�6>R�j�����5��d�3��O/"3���8U�� q.�XL�&!�#�ɛ(����#Dg۔��ڗm���c� �~l�8�]S3���If����Q�ϊC���Fq��cy������6qۯs�����U���^͈}1��+A��?�B��xO���o��q[���W��$<��yM�;�űW��9�g����N�l��E��.Y�@Oe�X+P�V��� �z	�I]��g�gӣ3XPPǊ��,i'�����t�<�ڤ�T� mbE�]�[��5����pHL�!5��<�U�a�6���h���{��*��o4���ؚ��<\�-k��T�*�с�e��}��Y�ƃS�������x�6>�l�~5�9��Ih���}����0���q��R��7�'.�ԯk��p����9<��k�L^1Es?ЪuϾgP9��4�{_l�c����	y?(��$	��y2 ���|��� �����������������ĺ����k�g��k7y��h>�1�ϗ���ժ�\�+�fȽ���%�y�H�@K����W�y��O�H۔�A� ]X�@B��j4mj�����CZ:�j�C���TM���5+��9�����<%=�c�ѽ�|�����y��-.�Z�����qo%������|��N�|����֭��>��Nf͞�&zXT��{;]j�u��]��T�j��H@��N<� Q��~-ƞ���O�y
�{P��ֵ�!� ߌ8�t��^#�׈gX?�-p���!�}�q��)d��sp�Z"��Z
�&��-���~o�)~5.�+�V���#}~Y�M��W� ^p����=���V��걤u_9���fZ���^��cuu�Ar�ըy^���;
�Y����rV��g���m�l)嵩,�w��ז�KΏŧS\���i!TN�1�]P�3S�p�i,[L�\�{Z*�:�J���@�h9*yL �D�d�Sˉ�sE�qUM	�����j��b�<R�g+���=���F��cC���@��qT@bv�pA/�+����9fO���m�>�D����lÃ��f
 "X��� �F�m&��n��^L:m}�^%����_�� �f%6����E�/`�$A`-Y +M@+E@M8W���Dq*�J� dt��&瓥�H�KMd{DD���f�hK���Uk�Q �D��)Q��ZU���E��X_WM�.��8S5�L�;S�/��������H��(Y /A 9��C��R/ ]/�	][����b�Y��LtY�ٯüŹ��rS��fUe�~@�B2��eҠ� ׶���I�E�_�pY�=-���ϐ���e)gjϓb,_�u���=���G"W֥�E���J5�Ou%e���\)��Ų̖m��7K���w��Se�P�f��ܴ�~j�q�@���W���ٌ�0����h�B֬_����'�Q�'8Ȉ��Y@ϙS��d+`[P
Mb Ux�g⤱�=\�����$ƏI�~��07	��'kY
� �:�w�+t�%20�P�8b܆��=�=m��%E��1H�<�[e�H���8(X��E[nrcͰ
�m�ٕ�8��M`�/G����ޜY!��zw����!lO�8�ek�l�x;��O)Oo��M9��W�oʕ��yb�.���%=9������7�uU�G����L�E�7H=3SYS��˨�o!��k7�`��}��m�	�<���Y\Lat��u%O��U��9���m���fR)[f	�M���y�^��a]X?�;k{s$;�C	����)t��Ɗv�гz|5;��`��l��ఎm���?���3�4�[1�;I���	X���94�b	0j�͢�b�).�x�EךF�+�>c!}�Һ��d�� ���dEF+�Ueh��a��Z�Oie�j�c��zV���V��<��}�o�(�'��ᚇ��o"��k�*��o�YqV�{Z��a�w(/y�k�M�Y��W��`$���ZW��t�!��n�={B`�I����t��3��/�'6��%W�;.��8+6儣�#���w��u���>g�@��O�6&o���]���י�. 8��Ĥ�Df�wey�@�̐�Z-7oW��\�dJ�N�1�ML\aI�&$���sZ6���8g��SZK@e��͘Z��kjG�܇`w�:�ků���f��#�4��2��aS������a��Nh��U-$�W�y�~����������_������@	�m=	k�AH��j�Y�go6���kṻ%<y W����>l��ٮU<�T����������jL�Z~h��K���Ȳ�Jx���<5�EE"xk�N�� ��?�����qm�6f�q�����s�c4�vk���z��ɋ��x��?W��i�AEo~՜�S]9�ٝ�#��e�|FL�Fڠ~���1��>vCn��G_�Z�;p�gP<y=���:~���n���u�o�H�EkhX���+�q)g��ʟ9���1c�(������ǿ,���=����ӝ����)O}���0�=���̤��NPI!�)]��/銵�a�z��Q�wR6��T<"�
��O<���u�b���(�S���08�����[�Cx9NQU8���ek��܆����>8�� �g��e��q���[�R\������u����5i�&
𜒗i]�i�p�%��g[�@d<���e�  ��Ќ�����ӛ�b&���q��� �J"}�3�R��Y��bD]�SΊG��ޯ�ٸ��S^'�i�~y��-T��NQ!UT�2�*�ݹ {����5\l센k^������ټOz˵�}N%qj�,��J�8wa^^�W�+&���"xzzߜ��w����J�9^�.4����ܞ�ɚ#u����`���w��Z`U�#��M���ݠ#ʬ'ܬ��U���[�����;�=j�ﭭts����<�t~�<�,���i�a�Ą�~�HSv������P2�Q�������	�)���c��k�A?�=5YD��}�d�.�A��f!K5�^�=F���D�V�@OA��FV��w��$O�����$Xރ�|��!O�/��1�ّx��xly1>Nd�i��k�1G܌<-�v@<�>N�J�D���!�P��`O6郹��~\���´n�%b(��O������D�
��e沏
�㎚�s��I?�|]q�P�ຜ���G�^��󢔧GI�\��a��Q��&JA^��@��GAR��?��������'�Փ8qT>�TR\݉qt%W i��QDر�{a��#@ޕ��!?/�}������L��sYY�#�r~�����<���u���؜B�8M�d�gҳg�|�8�z51q�֭]���H�ED��H��Ȱ��Lnn���"�*�Gʶ��3l�`FΔ��3}&+/e��9�e��O��m�e�[���yĻy��wc���Y1P�'����\�6�s��qb�(�ʑ�c�?�sBx��+;��I����>���s`~;gt���C8�t �V�����[���U̯ͤ_r4���b@C;q~A$ŉ��hcK��%�PRV�98g7�iY�a��c���*�hK������m�uE���j�@���5}9�y4���#� ̧V�c��?����I�`{m��%Y �Qcb���άgɘ��V�ܡ�Zؗu�[Y6Z�۸
��;�#���`O�Mc�F-ؾ�3P3��C���=���Q"���������!X���rT��Ū�s�HH���K�ޅ�]X3���S[ٹl<G7�e����0��+��u�P&wt����r��F>�;A໔W�9���k�$������-q�5���q�_��%����y��&�U�o8/
�VY,t�ZH�<��t�k10o
�]'����U�2w�@^0O�y�e�3.AZ~�S�)0�9�s�я=b����i��C��^yW[�=�"ul�%���6״���XV�eXA]C�5]��Vt��-0���D���1E��i�567)�y��UX�}������k�������k��Л�^}������H�?��!�)����~c��<�Wos��W��m?�6���-��^Ƹ�˹��q~���	a�ΐ�l���)�>[O΀V��$�[Q]K2�Ͽ1�O>��W�ܟ�d���ya&����ª�\��KR���($��̉|(���$>0E�8�_�:���%��B�
as88�77o�{�vתA{��_@ޏ�_��2O.�͑�t���p((�����.|d/��5�[��<�ǻ�4>5�ow�ւw����#'0z�jGͯ�)  ��IDAT$�m$�����J@Mޕ��U�ѿ?����8gˮ�d��4,���~�˶P�xESƓ4l(���k���q4��rz�J�o�p���z8�pK1���4���e�3A�� _��7���'�-�/�����_��3��h�����S�Ea9���*j����xn��'g�b�M���K`�]�fæf��h,�X�|1IA�w��#��גG��ߠ"L��+�5��TG��7>�v��O}�������>��Y�%-�G�/i�)��L[�{�B���8���!q��qk�!�
��R��r����D����e$�%�I��`�1���:�\������r�[0G�T��j�{y귒+�,����qxj�c���8(����$�T�wA�	��
~	y�\�sK�EQg�x�7X�~��p>�+���"+$^��H1���ьL�fq���b�WT�݅A��R3�=W�'��Չz>�V�3�Y��A_�%A$��`pv�Z�T��o���"F�S�Zn1$��KQ���G@N�d�vQ�����-bD9���#^���	Ab���W�'fĐ ��>%��F"-F-���B*��f�*X�$ڦH4���>�@�I#a6�p+���d���� ���;A1Ҧu�F�Y��kX�~Ѻ�c"��J�kY�iq�{��/����S�JͮU�"�ޗzV5�Q�R�Ѝ�v'\��u"-ȓj��զp��l�5^���E88.
Z� �Y�#�NY�y�?D�ߋ�bT5Fh�w�.E.�T�.T��,5�N�[��c'ܩ��j��[�V|J�ܛ�Ѽ����D��h��00�q!4J-�s9��9gJ�J�J�!�tu%�MTu$��I�;U�Eu��/���3tw`�Բ^�}��b��	���;�fu˻24�"gp��R����Ğ��虑O��7������>�wSP�Z��ge�����3�Cc��ͦ�+X�d�6k\��4���k�X����S�WS=�ƍ"Q�rh�� @�⌎<���zĐ��=�`�����7���'��k�ǯ��/���o^��O��֫g���~�Zƨ�855�-�Y��Dwo���{��gq��ݼ��QM^������߇y��:.����B�c9�[ ��xy�>$��#c�Hy�����Uޡ��)� r��N򷪳*�c��J���~ݛy���o��ŅX�K'�ѫ'�招|��=�W�ệ���������;ܿw��˧�M��|�C�&��M������𵳼s�?|��T:�G������˼��i>z�sƵR_���uۘ�0Hv����.�J�U��R��%uL-�=]����-�H=cSe���<!�7R��X=k��wn��g���߼��~�_���>��/]b媉dE��l�9K�`�6v��5�7�����+�"��vP�nb��Z���h����g��\��ϺEȺh-E��n�@�OUA�q�U��s�+Ѻj �s:败����͏�=Qr�%��AZ��c~�p1�Q��no�=��):`�ԃ]�����������$F��S�Dw���;āmG%;>�{���8"��&㚕�����z��c�;�����I�n=�6�KW�6q�.`��l<~���^a��s,��-�/��kx��Ϲr��|�U�>x��������x�9ƿ����\d���V^|c!���4k.E'ڥ��d&��+_lf�ɁTm�u��_\�sog�vFO+fÈ�����9��������ol�p��賯C�4��cj1���h��!�c�7�پCh����C��eGՒ��w_��Y�ň�䂧�;�v~-���9���y��G1����Y���D�(��\L��i���q���Xz�@W�JpeE���}�":vlbҾ]�ٴ�����{�V�;�`o�����Z|����&�^�N@�A��G�]VDvG0/|6�O����!L]���~<������O\#f|����y��`���s|��K����N����>��l&G����]A���
1u�E�]�r.�	8
�����^&/��D�z�]0��+�4�[���� �X��q�DR���_H�O��.���`�+��_����`]-!�"���5���Exx;QDF�#$��0k�x�ݰc� .(�D}2)�4r,���v��^I�.�ź(�L����Su6i1�W����=��z?��Q���f`���%�)�{,��；���L�������L^͹�1l6�i���E�&r�l(�]���jGݍ\/�cv�FB��������1,�jgcMk���?0��v6�k}���u|r��O�V�냕����g����ȓ��
�$���zz�#F���p0�h	�����u��&*v��u�@G�Z��?E�/�M�/D(�����	TSJ�l�h���T.Y��'�z�E1$��gQ�Ȫ�QuG[M��@5$-!Jk����<�iA�#B��#B#�h�Ժ�T�qZ���d;�pz����e�pu�l��sr�(�H�Ù(ogb}]<���� ��RK$�ژ;-�������r1�ݝ�^~���2\�o��)������k]����ڻW]ê[t�W ��aZ9z�籨�<yj��U��9b���d���#5n�X�Bg_-_���g-h�vbd�\5�uv%ӭ�r��;)ɑ�O�	��s�yb�ImV�E�Re��*�e%K&�d��q����i�Y<yk�Lb�ҹ�1���"�.:���dͺ-$�gh�@�ɇ[�@�� ��&=q�C�$2<Lk�+HJ�KJ;.g��YZZ����k�0q�H�,���E�Y�t&Ӧ�b영�=�~���V�O�I�*ߛo��P�Ͼ�iR��\�H��Gb	>��y������C��s�/��Ϗx��-�Ų�J>]��9q�4�ݸ�a:��c���/��?������?��C���_�������-�|��G��+�{�>��-��D�9�[���ɉ���Pץ��ne��QC{S-�Ft0tX���E�Ψ���u�
{i0��̬[4��~����-�y�o>z�Go<χ�^�����W_��7�j�J�-V&��ߺn7��0m2]��\��>%VR����i� ���?��������W�����s�b�VUrt������^4�%j�aLz5�]hl�Fjjݪ���)��"����ߧ݊K0x�R����s�U,�˅��w��w_<��^�ݷ�����p��s�}�&o��,�>�|����
	���y��z���Z��bs^�s�W���W������&���O��4�{I��|�+�{~1�� �W��]��O�6�N��[.�H͂=  �Bk)`T]�����:m��Z*9�f��L�6s��ʑ�(vy���ꭵ����=�uM\�2}|���w�'<�/q���7�2H�U�$;��̚�b��)!I���b��+�cP��zD_݄[Yw�J�	�ћ�	3�zӶ��ʃ7�����x�:;��ԵKܺ�<�~�ur���<����8w��_�KR^n��*��͝�������׿}��~�?����k���f)��՗;�wy'����c���0��'S7v �V��y|9�=j5�7��Cw���8&�θ��:e.O���K�=y#9�mq|��Z���T��J燔"�M���S���5���l�����S�{,��?��u��Z:�m���w�h@Oȅ?���!��Qz�|�m�5K�Ę6�q�Ƒݯ��V��ȇhGW�Dx��X�7�{���{�K�ü���pI���ԇ��>��Z�V�c��@�иY>���;!b��]Z	�1�����6E��r���:ˊ����~��5���K�)���?��J���?��_L��d;�D��Q>a"c�dť�l�|�EG�0m�.��N"�����l�d镚�Kl*�av�-�BEIkJî�i�(j���V����U��DW_Rݼ�p�#�U�c	���$�B�[0�R�z��S�i��T��RQ��F2�?�A����e�_2C�S��H���>q"1���ߑ��d�xg��.�gA`+䛩ʵ]��.�t�a�R,�Z�i]5����'^����ª@�g�`?��y��M��&~b��8�!�U�u`��?;�����5�i�Fs�6k���Sr�Qg?Έ7H�?�-@�^���,t�!r��	a,���V;':�RkfY�������p_�m�����K�|~B��b>�SƭIq�-�e�ف�F/�F"|ē�� �A �Q����������E���n��_;�h"�j"����+Q�4Z��\�����.�U�z�\\5�T�"�Kʑ��&�k���u�	���V@�n����t��ˉ om�@��R��
�0���ĆY�.d{H�F_n��1��ދ��_@��htQ�]IM��"�߃x2uy�z
��zzkݢ��5�ݑp9�j=���qk(����w䢼�[Έ2$���Ʃ��*x�MΡ����eQh��e?������<Ւ����r�㚏�MbDT~�1��nbh������u$B�.J�q�c�cc�=�u��$^�%��Q�䈔����ݟR�+jL^����m�+����t���O�+�Ȥ�=9�a�o��gOp��]ܽu���]������KWx텫�Z8����d��z�*�+�{
�F��T��i#ٵsW/��gnq��)�_����8t`Sƍa���L��ɳs7���%,H/��ĩڶ���]����Zt����_���N[~��O5�u�<G'$�@cm=���2}[ �)Ψg֨~�t���4_~v_[>{�8^���>�G���nr��VFf沾����>Ť����Y�y��->|�_|�6���'�������o��7�����y���<�,#�k�2�y�^ښ�#Eg�E`nޢY:����x����W���^���_�߾�W�}č+��&ߠQ��yC���ڔ`+#�{�}�|vlYƪeKY<o��f��L;���g0s�lm��<a�x�,_�54'/ң�Y42{nb���lܲ�-�w�m�^6�9}"�v�n���h�/�ɹ�1r>OuLcnvm��lؿ�o>���R6�q�o?������G��٧�r��J����j�B���@qX��es&r��!��%�� GϞ`͞M�پ��{6st�F��&Rb����<�l�Rry��Ǟv��u�T�:��t'j���j�vYl�u�Hn����r�'��~�<r�3�{zq�2&H}���Aw���D/�p@�=�&�y)����#�G��~��^VK����n�`<;\�H�Z���6��;S�s~�v��ɜ�����C�`C�!�4�%Q��B\r<~1����HI�7�S�zL��-���b�ш^�h�=�cg2|���;ʙ�/������b���l��z�$;��t�;����=ϼ����'� P������S7Xu�W�y�w?}�?s�Xď��X-um��;/���[�p��Wx��OyR�p؂Y����̍����^��T�f�n��h:��e��J��i`�|��#Gp���ג2��)�_���|����
�
x>,^ /J /B /���T��eݿ������\����1�|\.�tX����'�LޔB�P<����x��$��Z���������U��ZZ�����~Ch_��QRy�m�ρ�w��u���Z�@���R������>�U��R�Dtu/«�����h�^ы��!Du��[���9�|��p����SW{��`��(��jn<?��L��OT�V�����:�{�c)�!�c)�0��c��w�Rv�~�CO?ϖ�W9p��#&a��\T�����.ո%�h�p=-���T(�� Q����`�T��V9nUL$D6CD��tqqѢwW�65��M��l�/`1�Ս�b��ɱ#�0�������s�b���,o9�Y�����X@i���ŎF�;�V�mud���.���u��������9&�_�q�%Hkz��i�YT+���sn?Ͱ��8+����OF�1�9w�-S]��UN�	'N�Q���Aޭ�+9�<����$��'���~�%��=��mS�i6�`��Vy:{'���7��"�9%�S#R�Y�Ǻ�ἰ��>��w��|s�_���7'���@w�]ԕ�="ls�)ؙR�3����qfj������*�sq��� �v�u��T�`�qj;%?C�c���Rwyj��18::����	g��NR^Ե;�dɶǢ�S������TK���6&P���.e5��K��[ ���Y���D����c��~j��
b�D�Q`�$�����ʹԽ*�U�Ѫ5�,�wu$G���j$I�S��%�	�DH�ܟ�,aq霍�&(��o����Q�gTNۧ�a\��1�ߦ��R]��~xȳ۽uZ�����1�r�ӟK>�I�*S������P��N)�ٲ>\�Q�<����7Zί��hKGK�ǋC�.u)K�j��+FLM)��+#��B9��#�e���K�o�)����ffj�3�<X8q�O��օ�=��g�8����s� �n���ͼ��Y���Lrhe��l[����\mF~��$�,�%���~��}�k>}�}~��W�������~���;6�N�0ysE/�4����b_r��d��)�Y<�g�������^�����'��կ��/���S�ټx	aR�:z����wi��N�s��HiJ�j�<| �fOf��1�ӟ�3ǰf�X�O����Rׅ��8N���9�ٜ�G� WZ�Lj�ɼq�Y={[�/YĆe�X�|f�׌ؼi(��#.(�#{Oӿ�P-�|��73&�׀�򕳼|�6o��wo_�Ƶ���8|t'[��c�ԩ���˹u��EG�z�j&�f##&���H�RI�N%-2���Lb#R��gb
G/e�*���I��5{16k$!�F��$'�	�V�ZSHM*$'����R2��ZLLL�!�w�HkF	���b��Ĕ2���UK����x�է��@��7y��gx楧�+˗�į���7�FϊzҬ��4�n�e�̙D�$�XUIc]-�mm���FUMw�UTRWRBQR"y�Z����L��X˝��ٖ��;�|�-z�5�ہ�����R�U+����"��9�9�-�����'D��y���+6^t�%q�z�O�E���n�?�H=�)�A�H�5��^�q���/Hyj�AO�w���Z�C0}w����a�F��y���h�	c�1�)�&X�[��.�t��&$>���cpNOſ��U�#�eX�pAC�ʮ����wx���t�uV�;��-;�w�0S�c��=�̘��]{��{/×,f�����w��Ek�����ΰ��e&l����'���0��oc�����K����ÿ�	#-��,Y�������#l�c��9����p�X�o;�-��?����W��;c9*v���~<|��Ͼƙ��LO��&̙�E�����QN9_��kc򾵤�<��V�3�vΛl�4�q8$�G;�	���y�F�c�����ǿ;!���Y쎈f���	�`�-��cy]'�#��3�F�j�b*���؂�����*���f�4ZW�`ι�Lj�6~>��c�v�MhU;�r���X�։��k�Cxea}�﫲�𮵄��+��r���'�U��ѕ��{_~;��k�:2�Q�뙱�;s�p�t)�~?�?����1�`��OZ�@�j�1�b�i#�����X��#w����`�����>�����/(A_T"�QE@j&n��]�!����C�E�K����/�&��B5�\uc�`�Νc�*ī���@�N�A@�I�]/18*�K�H�T��b�ƈLoj���HsD���y
�5Y*�B�i�C ��$��U�~�:r���!G5��Wkr���U�`��Y]$W��b@�A�
��ع'�E9��;'�I�d</��,���.>�rR9hݵ�ڸ1�j����+��'���e�h�:Ql'=�����N���2q�S<A/=�|�9���n���\�?�b�<��;�2yae1g&������<1�C켿���^̗�Z��x_�n���Z��B/~{���הp���]%��N�p�639~��]5�Q���;�;w�{w�gv�� �X��S�*ϩ��g@{y�E�����*�)����S�<�����r����_��-~?�\�q���buuu���M�����쉧8�����	�ރ�'?�Ew���D��T*?'Gyf/m�{� `�l+
�Sb$��G�J�d��{d9AF�+_�_�¤�[��c溣��o�8f�b��Bc[;�2q
#G�����Z����Yk�;`a���Iq��d��^�n�<�	�F*��]}ǭq�B��S�'b<;� V	8�J��fu�̪`ql:��Z��ؗ�u�N��PR��Ws�{��ZX���T3i��Z�x
:38��+��Q����ݝPo������*2����m������u���W�25��XXL� 搪�잷���"��;=�F_1P
���}5�lP}+cz�gɔ��7���rFf3=*���,�!��k+baX.�V�0�����T3����}z1c�@f�����6l8%݈��ԯ��G��ŀ����$����j�(�"��Aτz%d�3>���,z�dИ�AmT-�ɜ���-�Bn���w7PAs\����L̢95���,��)KI�Kf����lԤ�{�x���F�'7$�܄L��S]�U�6����ݺ�T^EQZI�L��d�a���ӵ��'�1�R_m�nN������'�ONl���4-"���$2��Bt��A�~^1m�@�r�a$���g��c��6F���bM&F�0]�8BV̺̾B����<\��g�LaGb9��I�R1��ʖ��Ȼ���B�������G_��;��i���K�,��]X1u	ݒ��1�����ԓ��Vё�>&M�$�3%��-� ���~�b衋�y�xA�{gJϋn} P���2*���|ڄ&5�i�ؤM��zP4�]L\u6�O��b��;�{b�d���Έ>)�(�T��J/V�� TжAt�q�/�}[s\Ρ򜫙�������r/G���6��K O y_�Q\]����&1V��l��;0Bƨ�:�J�q�f�u��\b����$�[%��^褎�+�	[��֟��㙰n5�.��ڛ����&m�π�)=��~�(��.�m�bz�ZN���6�ƙsi�5����fȺmY��A+7�k�r�d���0p�V��̗��ȏ��_z?�k��|����e3h����9�hY�F����58��L~��&����r�B��2��|�J~���|�M;���;��A�8o,���ټ+��w�Z?��Et�i�<�1���#��#xs��]+�'���=���򿅼����|���<�z	{��ة�T�W�S�C\	_G�񨬜�fNc��y�(*��ܥp;W�ZЅ:Q���e����͟GƐQD6 ��/&<ceƮt��
���`�ZY�������"�;З֢/����)�um"��7������O ���!d��o��˝�Wq��z�<������G_���7r��ʬrj��Kl�vlE�H���%H��R�Nb�@r[G�]
ǈ��8��C��8C��3��]�Tʢr�œt���5"���vR-1�H%�q�<e�Tw�E���=� ��zR&ƴL��j�S���\���J�l�)F��Ho12�Xzce�)��gj������_K�T�2���~�� 
c��>�D8, ���YE*�c�S�wN*�{y�Y���(���T`�={R��']�(@q;0�ˮ���9+�zH��"+���u�=!�r�������!o�%���&m����iQ*�T���mT&�VYD�X�XP����xyi�l-�ʼ,1!֓u6�]ҕϏ���پ|w���ԇ?]��O��������|��ۍ�f�q�O�
�a�b�Ń_�"E�����?���ߝ��L�	TuB��]�
��~�_ ���1�=n��`�y�s����S4��o��ꊛ�j�e롺wW��q�j����f"̠Ə
��:�FXD0!!V���N�Z�Uq��u.T��
3RD�ٗ2c u+j"�J��Q-xc�
�I1����W�x2(�s�&{���sE�ٶ�ic&1��P��[�;G�����2r��ȩ��`�!�u��f���^R~����C+t4����M���
CuM�K����>�RӇ[���Rϋ�}�٣Ovi�aQ/6s�{O��n�݆���k$������{'�9S���I��Qƅ5�hN�'��G ��8i�^bt]}�ɺ��Ҥ4rc�T�G�բ��`xu���26���릕3N��k؈x��D�(p�a	�\`��(�� +K�����|=g��*�J���/� >���|ڋ�޽������g��D�9��c��� oHCo
y>����!�莫�`���м*Ɣ�2�����hIʦ:2�R����\.��Ο�X���d�=��r�ڰHz�e3Xt~GN�E7�H\Uà�&�s�ȵRT;��.�8�f��۵���T�b�c(Lɥ������
+(J�&Q�.D��M�LqZ�@[j�r��-����&��F�Яk9�%�t�j���{a�IYd��')� 4�FQR��v��]���H1�k�ܯ�Z���+�����m��B���pq("�QROl�=D_��)v��E;8�:�=EM�����3� :�At��82zхA�fq�l�q��t4��'��@���,�����y�'���m���5�L���B�@��`q���h�3y%/L���Hq�ͱ�-������ġWc��D͖�T������eѳ�n;p�5X�����TmB�UY��@�s���:<]�5�ӏ�AV��Zŉ7q��	�~F�MK����N<�']�4{s�U�w�c�pNew��śx~�Y����5�	r�1b&�$0���]*��?�V3��H\b���^�&��c�,�}�X�?�m���_������Y�/XJٰ	��L�����}<��&�:h2�æ�7r)F�>`��G�3d$����Lì���_J�����1��qS(1��3�>p0Ͼ���k���"���Y|��tV��ː6��"}�-~ob���=�����Ϸ�1�Ͽ��7ZȟY,�2L`��������
'u�Խs{���ꦝ<=��*���_���}B)7â9��)���Q<T��/���	�=n��@O����_� �����
��Y
�[�}�ݰ,>��ɥ�#Y>g:}�Wو[��5���c�&�e��c�������NPyl�E�Դa��V#��A�SMo-౭����؄֭���������K���S3i��ѕ�c�"
�;%�#+8xa_�i?��?�F�c#��q�|��5�il�V�!����TV+�i!��@B�;�m'�y �������hR̦��e,:p��'N3n�6�[�y��`��aW<�3q�E�n�`�a�PG���Pn� O��lы��@*tq��-�� ���7�ѝ]
���"1z�}5�[��A�Y�Q�m�J�[@O�\U!J��
yZ���w�+��^q&N;�uj���R�,�W]dg����Ӧ��	��\�pF<�,��Z��8��m����9O�ų3�^SF����Z���<�w�1�xJ
�Tw�R1������D���_�nm�цr��Ս�����@���<����K��`-�=��w�{𧫽����S��������OV���r^��Ʃf��z�$����������K^�+v/1�nNx@��"N*w�O��U>Rg+%?A�ֽ��j	�lY{,������S�d��*'�=���O���.�]��)� �䗿5Q�>*��8jr����&k�ٜ�r��l�zw����IK��M� c���6ή�э�(:�ʹD��LW[ UyMV=#m��yk-�c��t��X:U.NJ��o�e��������"Y���@��]��@!	!N��wwwwwwww���qW\����3{��>��};�oZ-��UW�}�k5
�uc��d5�e��z��ڌ�8�v������a�[K:����l X"���X\V6�}�o�5����<i�Z��v�\	��}0%�bh�G?HxX2ғ�i��1�}f���{Zof���q|ӈ	f�Z�^cs�Q�6/�^#VO�Ofx�v�;k�m�� �A8M%��K�nDQ��f%Qټ�f9y��.e����Fjq+:,@3�����:�Ԏ��om�}C5�	�B��h[X���:c
���aw��,J̥{h�����q�"ئ=��Laۂyl�5�I�usH���eE��3�s�nܼ�	-rJ�/@ۼ�P�]�Ó��h*g�9���y��ʤkI��O����R^�|��˫�9�0��Yy�� )"��T9U9=[7�mQ=�;6-�}y����
�pv�yzTvg����J+ T��JHb���toݞ��8r���ܲ��5�a�(<��p��E��8���K;�'�̩�i�[������C8�{?s�O�yAM��H��H���u����{Uem�k8�0Q��ʙ���$���-�V�d��7N���SSg�V-0�r�o��;7��d&��<�����e�JF䵢}�zt�l�ݯ����^6�r^|�����ji��(�T@�G(�����@Nn�D��@���NSt�M���̤�ca�"�!�%-7��51�!}3�qy�n��J�8�	�1��Q-n�pDߟ��\�����\u���������ӧD?2��q ��Z�C�{��},��˷�\\nu�l��u���+G6�=mxU���[��Eγ�ؓ���ȷ��jsO�x�1��6�vc��Lnߛ�!t����o��|=��(i�LX@�vN�zI^Z�&11ئg�UR�{~��A	�r�NS0�QN�5���댥d�CDE7�T�&��A�	,�C@Y7|K��_R%�W9�J3�&�^ي�v]4Vi2P �G_mph��n%}J�f��BK�E���=�>�qU�Dw@H���R+����f
P-���ޜ�ւ�{Z�h�0v��Ƀ�����|�cgN_�FA�B�r
p)m��V�c�&M�l�A\�j��l�$��͇��Μq�b����r/��=�/ �@�_O�����8/%���q���)��o!�����7��<�M0J�K-�~�~45�n�VR2b���9$g�$�D�����Ze��#;wI������JJ�&�اhR�qj\$/�D�Q�q|F��6H�P �0"A"C.��I��B�!���6�u2ٰ���Sh���8�cr�����&�f�b�8���MJ$�s+����|@g�:� �I+�Һ`֨�yʹ����G1�i�@\���$j�L�k���?Ʈ�{HiБZ&6ԖD�]�B��^GO��R���L8Q2GyY{9z������5�kȫ��3� o���V�'��<I���<��!O����u�@�z]�j�fzڀy{u��gl�jS[V{�bi��oИ����s��{,L�ji�:��w��ќ1�R�q�7�z��Dfq��d��t`����!O2�R�S#k�Z�0B R5���Ql�Ҏ�<ZYΝy)�Zܘ3c1)љ2s�mt�m��Aܘ����iC6�m����2^����ּ:]	��d[^oo���;,���٘���4G�':12ڞ��4�!�ݔHKyW�:8		�
�����OI��S����t�=�f���{���}��	y��w��{m����S�vj?����D
�TM���>�&�h^ռ�~k�����ps ��F�mV�C��h�fB�0;��z�7ڛ6!�4��B/kr�-�P�[����̴sc���V����[r�΃%��;�h��*�T^֊q��#��!��ۺ��%�Ql
�ך��
�J�b�)�J�b���z#3vI�H��#�3]j�syW7�bh����t��,YW}]sE�E�$��/��)�����&ۊD�^���|ѐ�Y�e=\�5�P�Wπ��1���Hb�������޶v����f��׊�� ��2k�\N�>A��b�ãت'�~�Z���;3�_�X���j���J�O0)!u��k%ɩ��5�[ׯҾY�$�]�{ ���T
�	PFE���J_��u3gs��!�>�ԡ��ز��c�q���K��(��ś�%7�F��A��l��yJr�J7`��N�ʅ�ٴn{�������<{����p���c�pn�$~�q�e��3a�d�\���sY<wk�c��L6���g�uo��1�-�����i)���)M ?=q�����&�pVZ
����K�6�%��Վ�AD2cG�`��$�4&O
��w�y�bl$-�T^��mX�h5=��$=!�Ƞz$�M�� �!��n�5�~]�%�kT��,��#�ϒQCG2v�|�3>�z��qq�R@G��st�ө.UŽH��OBd6��n�4�7���{Q7({�1g3tm�ҵ�Z`���Q��K]+j	�d�ej5r	u��R���i�=}�������K-ܜ��2q�B��2�1�rt�}U_�.���^�9p&��Neu�N7�G���U�)�b�r)��/�Zr�:Z�;G؎ĥs�Qc���嘀�)�H����p�.�Wp�#�s�Wdr9��sQ��NȨ�&{/�w�8�Rqn����n\,�ȹ�6��h����l��vS�<��ac�~l8�a�U�ע��������O�aVt����x�a��qX6���(d�X�'�/�������8K�e���t����]��\3f\����[|�:iR��Lmk�i%�J*	(nV���^^h�6�T��'�߂f�7�@�6]�hՙz��ݮ?A��6Q�����t޽�͛7}��eO���NiB+��۴
��\|�?w4O��������3�S5����{�sZG�������9���h��oE;̲˱*iF���l����}��kZ%����O�n���9�@���
�-��_@��j�}��1>���;��{<��+�����.�ّ3L?�6�����gS��3��mb��Ķ���mF�`%��ʹ��Y�C��l��3�����=3O�]sI/ŭIs�7�"�s�dv�qɹZ͛��b�f�S++����J�������cr�(l�MY�2*2	l�݈H�
��@�y� �$P&ɍ�Gu�2zN	�o���͑l9ԛ�˺S�V�<��̎8ȽX���XBn�q_����R8��9��թ��DL��0t�=0tv���)%Y�[S���� O�\���j��5SՐ�&�y�������[�Hs��4H4Z׌qv�E��T-�l�6W m�HՔ���C����AG@Oω��.�#�̽4�S����ڄ�fL��nO��3��#�sq�\v�d��VwH�:�V66egyf{ՖLڇ������$�+dqq�,vH��.������!�N����ʗ���0�34���%�\��h+�J�%)ܞ�Ų<�-�]d��Iw���D>�ׄG�3�mc>?�����Vp�o���u)�]���p[8Ԛ������dn��B�P��gC�3�R�k˄psF����Ϛro[�],I�1�������O��V��ib& h���)f��ZZ`ff�������U�r������\lL�A]#L�060��kP-]٦#� ]���C����q5��:zj���݇�*��0��>�Z�>YWPi(��A�����Z&��	�6s�I�ڦLn�ɨ$G&g�2>͗Aq��r��ߖ|3��۱^J��$�R�s���į����`�Wm��4�yj@���9]$��ז���Zs�Q;�iŜ-��l���[���gnB2�c[��X9�F�I��=��#{�.߉�A���O]U ��Z���>Zͷ�|S�p����i$qځ��.̕g� ����OV���;uR9҈�~��.$ �<.�=�W�,1oS{��G7"Hy+��"7%���e4���G�V�Ʀбik.����u;��m�r��Jj`�֍�}a=�����+!nDz�R�3P ��I^R*�d���ugB��,1]
�4r�c�*r����%�AE�t�hN�Vm��m�9L5�U�VR?�-������*m���:�s�$�����Y�h�f�����c�8w�4W/_�ރG�)yȗ?<����l���K��˻)�д�Z��ݓ'���N_���#'ػc��������������[4�w�U�9��Q)�O���!�)�4+l!P8���3�Nf��y�6���|�2��� ,���G���я��d��I���c��th�Y@��iŔ�Ӯ�5��j[��])Ϯ�0��U׳n��6iAz��c�HkAi�^�5���fӿ��t��᳨*������Q�\�ue�֣�0�TyO���$�f���Mq�2�$O��."!�1�YET7������l⢒(/l�̩�5y!��uȈ�e�������Ǵ��C���Ɣ��NF�<:�dr�y�t���Ɯ��9a5��c~�|�f6��I��1~)ק����5|2s_��ϱ#Y��٬V|u�?���u_X'ල~c>�;��?f[ߙ,JmùN�d�Z>������ٸE�k߇�u��ܥ�Wla߲X��kr�V����M����3ײf�,����k81S:0�'��V.t��`Px}�2�
���ݍ�NN�����h�����]� wn�e�֭l�p��3��+����ϒ��ĭ�7Ƀ\��4�eʒ�OIK<+��P��|<���N`Y���'qǧ��?�&`�U���.ZS����&�,X[ų��5�Y/�����4�׀�B��ঝ*i���Bm����כy�d�ot`ʊ!4�ؙ��VZ�p�#h?v$ݦO$��R�O[y'Υ��*kK����������s;�	�\�����>'?��pc�Bx�L���1�B�(T;�Ju�<�&����7.p���_��O���Ͼ�;_0g�6;�КY��phR�pِ�Z�Xa���aRfu�P�[�|�$�GF��O�$Bn��4N�5-]]딒����&� �F������*�y4�s/:M����k��q��a�~)�>Ɔ}'Y��0��neΆ���y�ev1b�R*$��d��"�ӘTjF4 a!:u��E�	�����y3y�z?�0���;Ф�	�э����1]"CnGͪu��m~���[<����_��Om<tj��')��9�:��" @�R�kTF�#����� B2�x٦ /S2�l��y��7����Yx��ͬi��6_��?A�ꓷN�Z���R�@��g!%���ڠ�P�:T����=Y�ӂ]�'���7��K��q ��cwRS&:�f�|���eOߑuf��'gkZrJ2�#���4C���W�S��Y�]kXa�N3b͉����Ϝ�]c�f{֦���4��bG�0�{�R�H�C�t��ǞA���0�W�i�k��\��}�yq�o�VC޻3��RW���v�m�ys��vW򛔶MO��!1\�Z�S�8\�J���ɾL�ucx�#��mh�kJSw#�\Mh�dA��)1�FԷ3���%��M�4�G �����E�vV�)���6x�[�" �l�YY�ha���A�L� 
}�u�3ԓ���6 Bպ} ���������5Ws�&r�x�%�`�Om��Xsr]Li�i�����Hwf]�Z��P��-��خkZF2��.�.҃�~N�std����I�S�d;�l�a. '�y[��C�O��Q���ϒ��̑w�\�)��$/��f�w]��;��̔YQ1\1�c��r�`���6�礩�U����Nv�=�~zr}�P�Y�Q�64�v�|���׾54s=���R#[��ۑnnK����̫-}�א���9Bkfh�A^Q�z�X��=K׳f�R\�m�˦isY;r";'�d��i��7�]#�qj�d�Kwpe�6O_��)�8��$��Ɋ	��WՖ^-� i���đS�<j#{�d��)L4���M=����2��X��.��u�63n�捘ˬ�3�u,&-bƘ�L5����2�g����ܙK?z}:�et�ќ�w�G��a��]�[��c��pw�I~�r����rk�)�=~C�'��� Ww�ç���G|t�2W���}W��mN[�GK�s�����������>��e[9�p�m����|}�\�8�6�a����O������'|r��n����\?|�G�?�����v�i��k~s���4��w����{��n=��Op��>��z�
g��eߦC��r��N~ą�g9�a</�?����ػa/'v����S\;{�+�?������q��sv�a�Q��͵7���w7_�����,�ocϲ}l]��K��k�i���}���4[$N�[��M�v����>�ޝr�k��o�A����~��+��x�v�<���c�1fMZ.�}.��m��������SrO'fmg�����3vpo�Y��?ȶ�k90k+_m>ϵ�SYX;�U��@�IN^���ά��Ʋ�m�<c	�w��TAW�Ǘpv��^����J��a~h�OZ��u�Vڏ�m����l�0�i��3?�9��p8Ȋ��Y/��k��,���%�X�`���e��U,�����70s�2fN[��E�Y�}]<���.~i@Չ���_w���1���*.Mk�sL(K�#�CW����΋'��E�|�(����DM�c'y�c��]A	�
�*4�ueb�C@��D���+e���]�_~9����%���Z��k��a9��3����.x'�3in%/^/L�3F��x{R[G���V�UG�SLf�fd�N`�T���!45��bǉ1�ҍ��n���n��d�Ð%��h&�];b���[Y;,%�{�{���d������1���a�C ��>V��� �����dz��w�_?�Ճ{��������e��=�	�z���_�]JA�%��H��QD�j������K*j��D�)J�ҼI�7Ε� ]B:�Y�x�i�l�,����N*&NJ����b����>�s�$a��1�=�%z"z.�y�P����w������x�����=��-{1t���J|�20�(¨n˝8v�=����_���C��0�_w�铡��ԝ��⚷�HW�m�R�s��Z���I�э���l�je�bT�>�a���Q��cg'Ћ0�!��T�}�2X��D�k� N2��y���P�l�3�u�̧�d�
���	y&�M��j�3� oqMs�I�\�||�j�T�X5�B���o&���9;�تgSmJ�܋�Nl���੬����%�=��,��!)1�4���YWى������p9�b��gTg{U�#riL��\�^|��ݺj��?!o��;,]�-�o��5�M�)��`c�F<�\�Í)��!�o�fs�{}ֳ$�A/�j�l��,������<\؄�g��b~Z]̟��x}�%�kg����=yu�|9~�ƫo'����<�ڟ�'��o��yy1?/�������/\&��`�;�s�ِnŚT;D�1��Ã-dM�`g��8P�fK��=%�Nz;���D�������=�>v$x���Ӂ(7{�8YboN��1~Fx٩Q���X[�,q���J��|�~��=t44��HG���K�Rr8t31���W�ͤP!�f�$Z���`E/G��ӫ�#��Y��ȖJN�����u9?,��C�872^�I���ڶ��	�]}Z���A
��if�akeZa���hnP]��⼇ܣ��pz�v����3S��Y��b�$����QS9���\7�o���9�W�:;9V�K��f���dH\��3�[ ���>���ٸr�Λ-�G88��ܔ��=��7f�|�����^+PLt���/�oD�#���{_R�;�ѣ�|ga:4v`r�~,�5��KV�y�z�.���	K�9|67��L�q3�7|_
������sz��0-��pɼ���r�]�v2{�fΘ���+�;{%��o`�����r�ͫ��t�
֭��9���8���<�j~֭��έX%��a���?���ضj[�[��m{ٲ�0˖ne�ʭ��v�{��x�F�o�ű���1c_�_��3��͘e�9m����ɜ��:k��^�����ըE�:aO8^���c��t�"�-��W3�r�>�����ϙy:{3Ofn�Y��i�
~���o�,�d��7�g�g�m��|��;O�C�}��\\�������ռ��'����ą�Y����k��,Z͒�s�:l� �rv4����-7�Eαd�B��ɒ	�Y2r
;��M2�Y#�2o�F�J�v=�ڪ�؃z�bP�ь2��}'����u�'m��Y���h7����h^��+=�.��h�h���C��ں?ݪ��]ԡ��[�c@�����K�J�'���o��toݗ^Ӳ�3U���}4��-e夅l�7��}&�ِ���6^ʢ�6p*W�M�ʀ1��5�fs��d�˽]��u��p�F��d`.+#3x4y�z�`n�\t�͹Z�LJ+�mǹ(P�Я��zpU�roN3V���&�����@�a���`ۑ�)���V<;�"X�Q�E�9\[���k�q�Z�L�Ʈi�6u�%ެ���u�V�a�j6LZÚ��X.з}�J槵��y0��ސ���(��Q���	}I��ᘜ�kz!����9�U�aþӜ��6l �� <���,hA���&V�&E|��6���~{��5�\��\�Zd�iR�2�
[P��){S�g($�?��2T┚����W1`�*��_M�>���t�}/q��I��b.+��I�R�ZvԬ��eжwkvOzs���ܻ�Lx�'/^������IT۶����j���ܮLdВ�O��nj�+y��bf/%��p���d�@����)�ۋ�
	�����D2����|t���p{�Q���ޣ�i?z<����y
����ѰM;�4�����)+;!h���x�K`K຦d�Lg�b��X )��\��*��y6��B��ˇ��$w����޽�{�
k����ChM�o�jF�߽T��j�C��/~������0�S~��[.�>ς][h7nB��U^<�q� �<������Q�>�˟O[��UW�x4�A�
�)8M���-�{o�5'�
�ڤ�.%�JITz�]EV��87l�qX8:~�k��$�v���=a�ZS���� zA��d�X��uʌJ5�)S*5���UrL���<��I&4N2��|�%�S�7��1�d������f5�))�FjT�2��]�V�D�Sό�z��1eVe��K�8^؞��'2Qѷ���P�9�).���1Q£�_ۚ�cg�ALn���ױG�<[g����\������*���V���Y��@�E���ȓ%��nt�t"VA�d�.�l�����|������������FV�{��cl��dܞF�v:i�����|23�/��p^
_/I揍ټ�SC��:ٖg��ו��~4YJ�D�X�|4��#�|>n��}����f��T��Y�:7����hT4���p�W$W��3W��,��e��	da�3����(���4p������H�H���cO�[��S�k$	�)�lS�����%�ב��^v$�[�lHv�#�՚TKR]�Ir6&��@�Z��XSbG��y��TԲ�u�%"��Ί�@�6�`�P��<��ȯ˲�aa*?,�^�ͣe9ܛ�ͥ�i����N���i�>����f��'S,��i��LO�	@�3���ɩ��ʘ����)�Q\c�۹2h+kG2�҅E6~,���Ήs8<e.kâ�'%��R0<=m�$�V}�6���l4����݂��3'T���7����Ђ��n�1wଥ=[]��cb�N���n��8�Bǐ�f���f�Ś�7r����T�Z�H����~�G9ohMc�IfT�VuC�w��#����	Iem`+��������Q�=u�*4��!�D9���B�w�5�W�	8&��b�A�k(юA4�R�{���i��K��s�O(�\BIv'�ܝhk<�e{ �^�����;��I�kmҜi�D�g���i�Qr���ɽE�-�m��K�}-6���\D1W�q'���d�rX:W�er)2�s��8��ͨ<nEqS��ф��Q����JB��J�����&\���Rx:W�3��Ý�f\�)�Ӹb�5i���6���ԇ�RbH�%6�1N�4u�be�d�&�V*?6*�D\�6D8yj���G�_(��I��K�k-҂��@�C�Wm�<��e�=�Ň�@홣=����K���pW"<��0����/<�[k���j���DNyEq�A[��o+���	�jS&�3�0Q`�G����u)u#�ԗl_
���~���Xωt���I��H���n4�q$�̛cGZ��bz`��'�XhG������hV������NO)`��?$�M~��8���m�t6�qw�xn��ͮ�e|V�	��
95`
_,�ɩ�"v�7bYrK	�_�؏��7J�[݋���d&iy�4�Gg��saI�ͩ�pew.�X��#�:d%Ǧ����U�����&�f��l#�-��a�
��]���3߰�.�u�]�1��E��⮙3�44�zu����1��Va�D�x�,��s��3k)1m����X�����;���MPA9��ex�>��x�Ľ�J�Kv3�"����O��{$�FOg̚,�w��7�r�럸��O<��g���O���6���+~~���?=��7����_�|�"�?8̣�W���ݬ�6��^�I�2��.C(�Ѕu[&�셪���W�x�v ��V��s���t��@�4���}	�{�)(%� ��v%��2���m��
q)m���u�ͣj|wv�B��ѬK�g� �6�>_�^
�� ��η
�h\U�>��O�����|{���a��%���hYٳ��@R�^�.����!��ƅxU	mW��R3��-�/��Zy���b������b�����1���r��_x*����^�y��뫾�7ɍkRħm��-�^=Ѥ�������ۯ�����X�??����~�B���o��q��h:􉦨���e�����Ql�RA|a*��Y��I�.N 69���p���s85)aҾ���k�i�nH�uc�)�/?l��𶱢���6b��=�)Г�n�4�k,P�D`��j�\�r}�<9���F�;���5 �� ����d]���Л%�7W�g~�B�2��L�B�Z*c۠k�6Cvd�гךhUәt��R����q��8�c�F�("���V���D�XTg��blT��K� ���C���6K/�մ� �U
lT�����]у>��`$ ��h��2�Ě���L��q�$���mH2�%�؄wK�rsnF5���U%�ߐy���;h�\t�4{n��:TDڲ�}N��ǭ�asy�(�o������nǋC=xsf�/��C��h�U����|ʒ���kѓy��L�I����<�ԅ�'���`'^�����<]Wȟ���eQ6?�m�w�Sx(�ywX�����ҥ>:Ep�k	WI��B�V�ņ&�˴cM�-��lY����l7�e�3?ف59ʉV�O��0;ɖqv2w��d|�㢝���&$:03˕����ueQ����#ˋ\��҇c=��<��5��e������v��xo��K^m�I\�sG�/j�x]���"�~��)�#�ޘ\��c��[�Ɯ����+r�x�hh��A���N�6�r�͔�8.���QcX���!�p����=�&��t��I&��,hƉ�˘�ތ�N!,2�a��;e�A^�\K�wu�yy��M��'͏�=S��[�O�8:!��q� v�;i~�'�c�\2�ऎ-�$#���!�"�~�
֓sG�P[OO3��<d�7������\�r��Ss�~�́��w�sYq�1�~c��fzc�W� S:�3!�!����9�!�y�p"���a{�%���Ԑ��"��X�	u1=(�q�!�@��T���=�*�,�o�<��Wfz�c��/�E}(W4HaK��J!�I _�Grע�����"�/�}�m��my��T���3K?>���}	���e�!�{���PT�m�'��<�]��ɶ��4��S�t��}�p~����=�՘Y~�:&$ظ!�X�V�����;�p��O�^jES,iR�SO�}��-1���J�4Q�KIy��4#��E�պ3��NZ�:� G��]�m$�m3'�=�fF��[50.�J@OΡL[�0d���U�p����h>��f�M��=�r��ĵ�݁�,f�s5V 7Z��:�g�8Q;�Sa��g�wgj�q�/�Ӿ1����{$\�W�d�C�k���O�z��G3F|�҇�^7s瘙'�`r��Ks=v�Z����[.Y�s���0w	$��7�{�wsa�NN�X�g��r}�~6�u�[,��jK�*�k�&s{�F	(����mk|�8 �v�ş#��,�#�8����P�q�ߒ5����:�3w���\�����)��9k�6�x��9l���5��`�<��CU\�d�?��~��4�����#:�؅��>*��l"�ޡ�f΢��������A�U�	����u�%�J@���R�iB`q�E�qh\�s~KͿ�Ez)�[~	mz2|�b6:��_|ɽ���g/��@E�zH��~�WHRRX�R�*��	I���W�������:�O�e�t�p9q�^�7���t�ޏ=���A<{�_~7����й�U4Ƴ�-��[������,��exeR�OL��7Ӽ{�.-`ȼ�;������VO �!�(;y2	'�� �lU<���
���wn��橣|q��7�$�gL�h�ܦ�$��=Q]�Ȩ�>�T�{�^�{v�&U�ڻ��������Σ���DmPFD����5W�-�ǳ�%7�\H����#��d�A�:�}���+E����c�ݹ�7�|�+����[޼���|��?����x�~;�/���u�d�u�a�� |�I����)��o���j�Y5�&%����3�%fVَ��2b�*<R���ed:n>�8i�*��;kaC����'O��m�F*����d�|�'�'��5�cUsm��5�\�&�u�XC�a5�#�N�� x�E��Cޢ�5�)қ%�R��\��6vg�dxʟ�!ɌwK��л>�Z�ܠI�A�9�6l�(t����\�v�lIܖHB|<����}��р��^֑LV�e�,�0��ss$���M`r�$�k�H�mh&�t�@g��ML��5��Dژb{&���L���������5������ڏwCB��p���R�C9��s欧#%xz%����/G�Fs~T#nMM���l~XV�o��dW{���=�.w���A��f,o~�g�y�bϟ����E_�����m*o~���/�����?�?
���D�Q_���Ii�5�n	�[�vkK^oj����kMS~^R�7s��rr
_���ᘆ<��Q�|16���6�1�|>��������tp�\�6����<���p�SNu���u8�=���"�14�ۣc�3&��&&rr_�K�וMx�)��;�xw�P�/�5�����zɽ��~�˽y~�-?o)��I�D���6���x%�N�zؒ�鬹�B��d�E|V�Nl%n:I<V͵ٲ_�o�f��#�S82p���HY;�7�f���7����^�Y[މ#�qb�4�7��5�u�U���ɏD���d�����@��5���3��ą��m���^]
���[G��2��,�J<5�@�}n	h)�˖߅�jK��
e������d�2.��В��|�c�Y9�3�״嚀�M��_Xz�[}��h�y� ?����s8��G���ڒ�r�&�2��^WB�$"�O"˶4�T՗)�|�����L>kԄ���� )����"1�R�W'^�ȗ�Y|ߨ�o��Ut_6��ӠX>	�`���<�o��m� � ��ȓ�&?���7���H��Go~4t����d��O�
\�fP����gkO����ƛ�]C��%�?���m0�څ�\��W��7N�<��ǟ39I3+�l�h`dM���N�Ԋ��l�US�W����r�J'_J�(u���Ɲ
�
�n��yM���@*�/2�B�����&�;i�cE����V��:�na-�fJ����O�My�-��9A`��]-��{��؛�<c�>*�Y����a�6�BLs���z|�U���¹�Z�Oخ[�k�;�a^���ϻ�w%��X�i�/���6��d�=Y�X��c#GM׍e.�~�̍�� ~�Б��<�\��rC��ͼ�.�����:���#���!a�q��\��9�F�d�>�y���&2;�	�Gs�*X��Z�k����Y�a {�M�p�>l��P�}�r�2�p:���V��e'����&�M���5�S������\ʶ���5o3;f�g��e,:�����p����B@��|���+i*���十�澵p�<�Z �04�&���5�,YJ��QD��)`���nx�t�B(��)h�oQ�9�ڸ wa��v8sԌI��d��ԭ�9{�+���W?�S�s�>���(&P��_�ݯ~�&��?~��>�ԍ��س�������К�203�5����_����F-,�V�,���'������)�_%e��R�U��b��q�՝زD��"�C��M�����iZ�����^�Eٻ�C^�d�U�S���=��W^����g8q���LЪ��roց�f����xS�%T���9�A���2�5)�x��OU���p5��vQ9]'Oa�������M�^������3޽y3�'Ք�����W���?��e~�=5i�����@�~��W8~x8[6���7$@r�dK�e�`�����,�34���ɢ�lM���㳩]ё+�0|�r�bc���8<�<cK�l��caE�d�
N�����5���'I@/[%ye�6���$sPM�m�	�� �'p7X��n�dT�����W�T �Z+�Tt���յz�(��{$��"�wD 﨔�7�K��Ӗ��{3���]���7c^X6KVr�Y͛�*)A���dIO��pX���gP6�T�ʢ�bN�Ϧ���s�d��'�%q]/�8��B��T�Ԡo=�{B��1��o���Q���E ok������Y�I�pS�,��i�H8�4�X�#	Ke�$�X�"+�d�bme(Gz�pqh#>�؈�s�vy2�l���R�ּ�؝������q
����?�^��[�ۗ��CY-��ռ�c���Z*I��V�d����r�"x<��ɻ����
�^=Û/���������yuy������N<>�A��S]�{zs�5.���b^�lʓC�<=Pγ���}K	l���M���smOd�Ŧ|�n/�}��_���-xwZ��b'�]�(��ۋ�ys������u�[��r\��3=�A��ւNH���U��M��﬍��� �Ǟx;�ukb*�gTCA��%���aA���K��&��6�X�����'Z8��~<����\�nlhЄu��o���m��e}j%�
;���@��4e��+�:��<��D��ǿ�1^���H���l�t吡�0�t�.�����r/�$n`اg���f�߫�����ՐwЯ.Ywkɷ(ߛx�w�S0�<z����)�`��X(�pL ✮��[pI�1����[4�u�"t	5V>rie�̥�~���s�H>1��m_؇����,���Z|�Y���A|��ՠ)=p�B�s-�9��2�y��ڝ._���ok��ƟV�}x$��6�ܵr�K�@����Ks~4q�{#[nHX�4�⾙;��|l�#�ж}aj/Ǻ������o^�����@�P؇q�"����\0��՞��z�,�}f�3���*P����R0K1���)K�|�]������:��a�R�׊a����2���@As�	g�Bv&�><�������NI���$s�ac��.�4�|�&\
��X�F���ބB�&��&.�519����GsأW\�lk8�ɽ����t�����ąH]s��]��D�0�zDHyrC`�/W�����}Om�cS�ypY
��.9hs�K&N�ݙ�r��s�y���梤���Um�+g��8'���^��G��� �j�.	�^1�⒳�:��5��'3?8�e�ׇM��T�O�ě�����`Q�ޱ��v�*�W�����]�6�ny@��^�'�f�(8����\s��}�{sl�l�/�ņqk�6m��'�r�B6N_��!S�Q�U��mו�%����A��//bqLH��A4�={���f�<FRU/B�[�^��[H��Wv#�s?R{�nU;mP�cnS
Z�T�=)$�4&���68��݇յu��W���%�W<��@&�����1����޾���/�r��;��}�)맑ܱ�%}kԱ��MbձٴQ�[N��(m�Nk|���XA@b:�gu�����Y7nVɦ=9��Ixc�;����6L���h���X]&����y�߈^�������׹t�,c.���Y�eں���h��դB3L�̋(�S`g�Z,��I.��Ӌq�.�j�<�k�T"��:{!7�x�K����K^<��7Ok�U?;u//_��@OM_�-7n|��d5��)
W�������k��Y~�q���\��s�b쇎OCk'
�a��E\VI��J�Zn��,G'4��A�9�՗t5L / ��pt��1pr��ޞ`kꘚQW�@I,�D�R��@T�W� �y"�����x����ҷ��$�5&�(���B���;䭫a����"�v];v8ɺ	jXrR>��x�-dS߱욱��SV���h�u��ɑK9�a$��0ۿ.��D����ܣ���r=eHy���2����K�PЉI��m��k���W����X�u�L|���`j���>^�zZmQ�X{6v��ek!�����4�_����L�p&�A���U�LW�}cjH�a.���K���m��ê6u�ӳ������zܝͣ�i�������\�d<+@6��?L��Sx�T��כ�6���:)�����Z��Z-�Z���%o��ۍ�b�,����E��	(�[ �  �J/��9��h\(%��{4V4��$9S�Q��H��qr�ɲ}(|/0���� פ@r�oOU��H�@])�����
�.�.�����ԉ�:��l;����M|s��������<;х_wWqoq�fh�А����\w��9�;џ6Q�Z_�X'3B�	12%��Hs�,��@�Z������ZW��R��b�5��W[83�Ԏi��,�f��sM�����r�����@�p� &��f�w(�-d_MNY���%�T�F��P�ah�y��o�F��&6�/��(���J<�)q�̏�YqT����!�i��v#{͵��ry�&V����f�P��)�r}e����'�C�0c�0R��Μ�<+��uk_θ�0\�]�jhN��]�]9��}� >�q�s���ul����g��wulx��-"�/�yS�}������[nհ�3G���v=�[����[�L�J$�帻�|G�=ҵ�k[>�a�m�%�~-��_YsSߜ��Ts�9�IS�[8p��S�{�����̃/̽�Z���������9a���L�kϖ{�h��R�{h�OA<��y����xf��j�ER����*����Y�o]z31��B9Ӵ9/�����|�P��������*淪p�Q>�'��El�:�����CN9��Tq7�?����܍/�N��D�p�A7"�j'�B����<�g����+�$n�e�Oߑb'�[9H��徧��j�Xn�{p���k�k:'����=j�rYσs5%NԴ�B��;y�GkXqRߞ�F�Н7u���f�G����*�X�pJ���4�ഉ'g��Y���Z�͵]gm.m\8���J��ޓ���8�����JY;�/�����l��o�G�'�볪����-���g���{kس=�_�:��S���gNK���߂��gql�BN��š�ػ� �v�����+Y6|&�`٘t��JۂV�j֎�m�������':��Z��甒NDU%÷nf����-�O)�y�;��kIPyg��+��`�.XDr��7kI`U'��� .�4һ�g��|�TUoUO�eT�����^�P���9}`���_����7���z�����p�w������$�f�����D7/�ny1���UуZ��7jD��
�U��ׄA�����~r�J9g���3�d֢�$�����~��0�Y�*8��=��ϛk�j��T������6��IN��Z�3��2��'�C?�h6�c͎�H��Ss��|Mj]�P}�԰ee#/�uO�n����~�Ջ'r�?%p�z"���Q5z��}lʝ�����a���K	i5��+>���,����/L=��w/y�����%����oN���}�>4�zI�0��04��<,�t�`�R�(�qA��]�Z�����}��cΎ-Ķ�²~4�!�x�a+%S�XYg����RG��Z��+���gJQMc�<C�K�Y%�5���F5���M��t�H��!o�,+)WtJKjk� y�$�SZ#	�:����7װ���Q�޾�Nl�fg�	왽��f0��@VL]����֤R�`1V�cu�,�:�q���]g�$l{$��#��S��m&y��P2'u�Ֆ�t�Z�U�{�̌p�2��Ą`3����#3J�17����pe_�N�yl�
����tpR�wz�n� ����+�S� ����ӌ�XO�0�2��914�+�r{z�6r��f�=U�9&�$��큼|8�7?M�?h��Z_�Wk%���l���Ub��N���U��N���R�Z,E�j�{�no_+��zjY�`�h��K��J��2��_O���S�zrܛU�D�P��4���v|)@�� ��A��ޝ���������N<;ܞ�Ǻ��npJt��H��d����m�|@���]x{���!��b~�X�7˲�11��}�{@2��^ψI�U�+)��؛0.�S�B��8ooF;81�֑��.̵tb������Iy�D��Xod�*3[-l��Z�%�,7Q��t$����B`σ
-�Ygd�v}CΚ��] /Aޯ���2W�^Ɩ,�qd���Y�/����l>ZI�Â��g�e���A���ad���KnAls�%�@U����"\
Y�R	�8� O5�����k�y{����sJ�^�M9)��b��I���%�	3��sԤ���A�I��$�[i58W\�H_2R=W��hͅWݸn��}3?>��! �tK ��C� �isM������)���=#'M�ܴ���\��s�#���,}��'�a����0̓�WsyFe�P9�W����]���,}�!U���-���!���^ҎJ=KZ�3/���&�/�B��9�'�a<��σ�8&�X�%�Y��%���}���{/6FEi5��:416�Bi+(k�~�Z�w><r�G9ׯ�u��>���j�C�܏����K-��E1#4��u[04�C<s���^���byb�����ܯiŧ��|d�U�:.|/ �{'=2U@*M�)�ĒpK+�0�Tό���}�R�+:v\�t򪡇��r��?輼�^\���t��G����,����F��<��딪�3�⼙��O��U��\��>k���]�w~ض�b�95q{%���ٌ�N����e;���5v7��j���{��ک7_:��vcX��'�~ӳ�|��\|�S�q������|�:.LY��AK8:e+�.c�ҝ�]�C1�|�<M�?ސV��m�MǢ6�o߇�MJ��D����p���q�M#T����i�NM��k��R��2U�|۫~����/���.�)6���:�B௲��A�'��^p��Is�􎗯����a���5xj�j�>����Z<�W��
��\M?��I1�6�A�US�^j�q�j��V�����+	o7P{&׈p�:3wm4W����ք7bκ���f*ц?�I^ӃWOF��LSFϊe��26/��œx�R����T�����S����H;H O�໗ϴf�+7�2h�4�ǛmN�miԥ�6��;�����2��d����U˾�@P� _|nIM��6�{O��ӷ�i�B�y�E��a��X��yj�}��A�d�z��~����z5}x1^��{��d��b��!�9O_�e��m�7����:��Z<��4jԮ�q�FX5���Q6�q��7��#Z4ʑgM���I�X��Ȓ
t<�������kI�B�l�I46�L�Hk���D1Jטt]3�$�i*�բ�m$��*�z�Pʹ5�Z��"U�� o�d(�7�3b�dj[dYs0-��f���{���5�%�X٨�mF���h����ɋY;n>K���^2����Ĺ���]=�s$�@2eG-c=�^G���UW6�T0�-�uf�Z-�
[g:�jk���36���Pd�ٚkQۙi��ϴaO�p��Ҕ/7����t�^�ϥ�����8o	s����&��8e_��P�oaH��))!N4�r�k�7C�<Yھ6[U�ް8�Lo�w��ue)O�4�����y�5O�t��Cx{oﾜ��D߉���
��& ��1��'���r�|uv
��
�]»Wx�T�����J���c9��晜��b��<��?N��ϳy�x	o�,��ox���7�W�L��O����<�=�7��}�����N��J����μ=ܑ7����H�>چw�Z��h3���١2��k����ym?�H���X��m�ѾQ�oW���~4�eL���:0!/�N1^dx���ڄ�^�,wr`��#��lYan�*���Ff�11��n�����岼NW��j�HA�rU�F�T��tY$��8�}���"UQ�]O����x�XS_�kc�G���k`�2K�Hᩥ���JEKM�$N�IW��L�Z������t�4��o]�yԖm55�S>l({y�_A��4�\�jr�Z�r�-�s��c��0�\��o����҅�QL��?N��7�������8��5�36ှ�M�l��G�wz�����H������$xSύO�=����m���x���>�w�� �}#<CoYv禱���'�x_ߋoL���B5�qWߝ-�&��OҀfV6d[��/ϰ�ęG��}�<|�c7~����04*/#�Oc���2�~��G���] ���[8��"/��F1GK�d�;���={��v���[�kF�ϗV@qK~0~(����/?Z����ro?�~e��wJ��jG�`��1�N�G�˩țNE�����H�B�x&p�.�_�K
�[�p�*�G�?�$�kd>g|1�Е"�+���ݨf�y��v�� u�OkH�@ǖ���IA�BM{.�:h���5�^�󩖁/W @���&8y��%�Ԡ�3RQ5{$�/Yxi�l��5����J�qE�S�y��t=�Ƚg�:���=��~��=�h5�g����u,w6��dEV�U�8$�m��gW�ao�
V��J�s���+��[���7s�:h6�n�;�ٍY�o*=S�p`����������o
��l`��uZM�걋��{m2��T mH�kٝ��h�%O0�	�%*	��<����=�fS'�۴XX"Ks+�kzfT�w�P�����)�;���ͨ߶�6*Uy�
�j��[����������j����s��x�������_Y���W�'Ҡ��k�'Ze����~��^e�ʃ����*a�"|�ci�-��'���ۡ��׎��X���aI}v�Ο�'�|~3�;7��~�3��v��Ѯ�5��v��/�ȵ7�7��[�$5t䕂���w��۟�a��Udt�H��6�巢�d�j����sj\�5ͪfZ��<+����Aj�E��Kʥ�� 6:�3	7��?���W oD�ٸ��X���[R��������Ǐ���/����Մ�~��R�g~/Uc��*��K	U����?��#�O\%��'Fz��F7�"&�z��M�H Gy�p��uN��"�OAKm�O�Y��4v�Rj�󭍮�'�N����x[k2�,H��LO�z��a@JM�<s*$��Pk_C_���[���Z�����d��Y���+�-�i�i�{-�a�i���
Q5��F~�^�o�k(�� P�@o�$d*�UfUv�i~>wyGp8�1Z���H��Y���}��0���eZ?�ͅ��ظ)�kk�2�6c[�����ڗU�A�5�b�d:��]�'����K�Z�Τ&n����(��ֵ�X�:�ٹ�,(r��������{[2y��������M]L�oX�#�R�E��җ05���T�� +����&8;X��lK-';Bl��u$'�x{����e=���������Yy��<�g[�Du�9�hɻ3mxs�=���]�7�§c��$x0���N�?L�����t���������Y���1�����9����t^�8�׿N��sy����6_ r.��c��,�㿞ȋ��x~W�(�;n
�]�ǻ�5��o����
^�n��=u{�����b~ޚ�W�3�bew�%�ɔ�|4���5���vt�d^ym���h�u��E�5�����pz�����B��-�$��g��![�Y'�`�J�H�+��+Z��j�j�N������m�H��y�<jY��]-RqH-�-�}'�  �ȱ����HW�;\��D�mYWͪ���"<=)��K����e]y��um5���H���$����r��j���<5�B���.�:��G�s\�ψ��7tA�Ew�-���8�_7T�N˼��l�xPӑO�e��\�o�ݚ�|VÒ�j���5w���8>5Ա�=��{�0PM�7-��67��uJj���wMl��x(��@��K/
 ޭa/״�����<���g�na�G���Vc�H�I�j>�R�4r�K�Z�����w�jg
��&ƇVգsY��,���羑�0����J!/Cς�r��u��w}���ם_'v���Ű����˯�q�����|��W������7���ڀ/\�8�Τ�<�2f��0��Y��:�S��H�W6]�Y��i��|$��Q�۾�^;A����Y�_�%KA����J�3K$T_����B��<�I7?6��t���Zs]�F�}{�#�TKޣ��. xC����g�M����>5��Sk5���T��->5r���,����dn��1	���Zq�����a���A�jȵ��\t�Ჱ�\�F�1��ݸ�P��vu9���u���%߹d��.�)��nA��1�,Ey�V��3��d���ɬN�ٴ��D�e�Z��Xǂ���^�^���m�1��`�R
�pD��S�7]�po�Mx��dJ��AN�987���I>^9���h9�3
50�K��13������������xߟ�������+޾z�3���������}�>p��� O�E�I���,Mo�����+��.|B�acI-�a����hş�&���`2ZD��4�q�r�s��8����{�כAܼӊ��1ce+��ˉ]9*��g����r�O�{� y���@�"\A.�a��|��[�9���b�/]��4h׋��V8f�kͰ�*�61Om� /͡q��"�`y
�<Ssi5Pn�{�;�?��KU����o^����������א'������}�3!ݏ����/E=��B^���G�DZH�󊞼�s�!��(�â��j��2�b����#�F)8'�h�|��`)�^Ҍ���t�Xl�4���/zΎ�w�G�m�(tt&B:�)D�-��ʭ��S5y�}�T-��V�7N2�I��L���L��8T��w��'�K�i�rU��a��VK"�F~�QO�u����1e�d.��>�kR��ch�)H"��Ȋ���̌H�҈y\����2Y�]���~̰��<I̷XٳK v��+;��T�1���=Y��:�6�c��7i���-5�D��5��1���1���o�������ϑA����9�mI�j��X۔}Pǁ,[#���Q��T2[C5@Ωd(�Mk����kk��lq��6.�akC-Ws����2&�_ಎ5�0� ��-%�</����$��ޣō�fy?��������9��������<ޅק���\g�\���K�yu�?o?*̋�x�i^��'�Ó[�y�P��� /n���e�Y��	� �7�G�C��»{���(�����+=yz�od�՞�wǪ��o���B�S��}My�������B�Z��gs}ZC.�����z��W�-�BXө6�|��F��2"�#aX�@��A����VL�x/�=�pwa���4S3����Ԓy��-�bf�Dc�J<��`�h�0�Đ�f,�^���kg�7�4�+Z;��֞Y�������х5.�r3��K��b�{m�9�R5��&�^�lpb�g�����gD��)�X ���Ԅ�VRp��s��S!�J�oa�DV9�s6 ��;
=X}$n����m� ]�!�T�^��[܂�o.q�ܚ�6vvpf�ĩCf�v�e���h�n�L͵���u�.Ϻ\uἓGm9d��A+g�^�)[�[�p�ƕÎr�䤓/�<k�@ �S)��y�[��u͹�k�=�%%���\4��z ��P�� �#=>�q�K�/>�T5a_[{s�-���>l3�猫�t��h�+�����U;^͕��T�A@D��V�h�3[xr��mC��<��,xf�S���*KZx�Yؓ!p�T c�K-�ͻ9�m�������\΅EqI�ϫ�I��l��b���A�0�H8�>��|f���MW�z��4	��.�:o�M7�W��Z��H�O��]�Ok)4�0��5�%ݭ�i*𯯽/O�7*}R5Ń��8��5��\2�����SwV`L���2{r������/RͰ�̥(i�S4I\��眀��������ū����'�ڜ$����* �U Z�w��"�h��p8��}]���s�ԁ6�\v���PNZ�p�!������\$<���N�w1�h8����f#+�=���d݄��j5��G�i�f�M[��=i�0�N9��y0]�w#,(;yO:���h��u����dL���.)����</_��((#��)�M
	,�c�
$_͐�6��������U�9{�Bu��x+��l|*����ן�x����ՠ�O@�'�]�+�{��/!<�B��`�j|# ����rKOQhq��y-�Ʒ���g���4��Rw�k3~Ug�|���s���<��3����l~}:��G*�8���=�����G�s��Tn]; �\y�B�C�z�B�L�iT�WB¢?�>eٮ=D�n���-hN�N}hЦ�faZ3V�[T�]b�6�Թqn�ӱIL�9�L3D蚜Oՠq���~�W�k�3PU��ZW@�w��dY��cz�\5�V?��=eú�?��˶r�֗<}�R�K����Z�L�����G�S�k:�Y�"��Z��X7L�*6�8Չ4Sf
t�қP>f��̣AQL��0r��F2�R�li*N���F6x�������3�������]g����e���S[�z"}�J�6A2��5�[�Z�$���Ib��g����"�4�� n�\G5�����պ��Sە���m
�6�q�6e�h�@�2{o�4iƵ���u
c��?��=ٮ� $�8b��V3�	�.NNd�ԩ[��Mg1�U��3�ik��di�վ��6;#���	�����W����[�s��"R�P��s1�lN��U]�ljN� b��[j�g��d�����˹ME��xYY�ek���)��}�8ۚ�b#׶6��ʀ`{C���i�@n�=Uum��Б�9��m���u��-�����8<�{�S�?#�o�7֌	��2��x�>��k3y���v���ޖ�9Pɫe<?X(��Ɂ���2���H[�m'���Do��ԠM����ӝh���h+�n�Z�rw!�w��5
x���?ץ��~\"Z��wr?��sov*��$rmt�Fs�s(�Z��Y0�JC��Bv� ��.���A7%U���J��q�,,� �c����@Q-o�$�26-�9��,�/bvq)3
J�-��Y��̖����ljՙ%���-eeEkVW�emU'V7���R�d�����Z1����J��L�,faq+[�gq�V�*���6��Tі�����Z���♐�ɚ�SX���fL+i����eg˵Y�[ļ����c~�L�sM�jʪ�v�l�S�Ӗ�9%�d�P�$�.�-�ߌ�%-� ��E��\R�Ȧ��ܮ+�ZwbU~�z�ck��*k�ζ��}K;�aV���m�Ms�ߥ�=��vdC���>��=���cg�̞��$|�r��0v����86y:�bGiS�ǥ�OOL|�Iǖ���|g������M����]4�a"���ғ?,^���\�0���N ����_l�L}��̋����F���!�o����=�Ǣ'΁�p	�sy�u ��=�
 �:��x�L�x<6��WC_~1�O,O����>���F�}p�~q<I�t�Ak.��L׷'A��	��>y�V���Ŝv�\�I�/P�/�W��9��F����A) ���ƿmC��ٰ���r�t%�`:���_��V[�i} �����;C�f��pʠ��/�k9�䘻QAF�0ңb�١#�Z4cPES����G�q��32�qR�љ�r�d��Zf�W�l��L��|z�S+���jTj|)��.���lJ�2Z��~6��*8�R���"�r :W�-�\Z%����|�����\�j�'%=�������JYw�$�s�����V�Q\hދ��p�yw���Ǚ�8�n �$����p��nןc��r�E?�u��Y����LfVU���p�?�&+q��O�;	,]�_�h�
GѬ��r�i��4�)#3q�4Zd��:)�1-;1J�q��T
C&>��E�␜!��Gh�V�v�Nx��H�PV�y�pmR�w^S�o�b
��2|�|���[�i��Kb�����B�J�i��3�i��|\Y�x*L���Wz����j`��lR��A�:�6�Z-"<~���)L��SN_�H�!��T�3����|�d}�#0/���;;�g��r�Vt�PAr�����{L[�l�ʶ������K�Rͤ�2"�C��<�d��J�����mzO����9IF!�s\�I��W�gV��Ն��ӕ��j�sK��$N���b�^��Ϫ��U�x�:B�3@x}���Gx�I��I��O?�ƌ���uG]��ok����o!￝��L���G7i�8���� ۄL�O���M|�@n:��9�'�i��sz&�kB$��u����{s�>T���n$�[�'��a���νU�p)�k�>%�5J���	���ْ *�SZ ���Nie3��i#i����5�ؠg�:}?C�3�:�o�3��ڬ_��]i�d���V�9�J��S ��أ��>]�{�d#��:1�ƞaqY�r%���s�o1u�|�����ܩ'��!ZS�I��Ժ�YbkECgR�k0!/�#�lθ(#>��/��~C2?m�������&��C��u�Z],����k��'�&�vz���xD*�s�3���W[�\��!w���#�Q��Θ���@�&�f4��u���ӣ�!��m���Z�đU����1���C8�7\ӹQ\����ܜԈO&Fs{F��5���$�Z��W�
Dy��M�fa�(]�5���|�@��Ͽ[��ټ�R�M雹�|9+�Ϧ6��I1|<.��##8?�.�Gp�$�zF��C���XX�Ìl�&82 ڞ�~Ƥ��l����fz�f�&������'�D�<Ϛ�K�euE-�ԦwC/�{PY;��G�o�D������S�5z
{G��Ԩٜ5��c�rb��N]Ɖa3��g'G�����\�����6qb�"NMX��髹0m秮~�������3V��u\����3Wse�.6����شt��,g��\����K�p�Z��X�r�sWr{�n�X��s��`=���м ܝ��O�����~�1�;ę�8�y�7�`����p��[��o�Qvo9���G��~���ɽyk�^���;�d�R>]���Vn�ẽ|��0��Ծ��?q���ry�qn��Ń�x�r+_��ʗ�������~�����,���3�x�:�;��6�u	�:�_u�#�N;�s�֛���\v
�}-.��s�ޟ3������C-ͦ�y��\���_ǽ�q>��<#�($�K~8�S�+1����7B�Ґ�u�X+�ۑ�|��1�9W8�=�p�>��~1|˝�>�-��F\���ܫ������	ڶs�1�7��r?9�6J�Yy�� �Ɓ����ᇰt����Ѻ�d蚐��O���i�Ӏ��$
<CI�s�ZBz���w�>N����m&��=�9!i�k���0lw����j}�'p�LBH1U�RP�ȧCl*(��II�"&�����۷h'����u8���Ʋ��0v4Wޟݥ�5���X�ۍM�}X[Ѓ�}� З�%rl�6�b}QM��ע���Oo���V�ε�y[m��N,��ʲ�.������ެ�����m5Z��vc��l k�zq�j${�eW���;^��7pGF-���e\�����qi��9.���Յ;�x�~n.�ϭ�{��|7Gg����ãV�ISq�]�I�fs6`����x��$4wrG�^4�\y���$Ť�N
{#[u�[��4�i��[�ޡXI!�5#��+[R�}'B������fZ�+��f��5�DkTr�,�#����
�ӊ�Iȥ������g��w����{v���_���]75H����_I����?���~�p���-o��)����s��d~�m�˅�M9ۗ��`�R7)�!c%o��=���Ǭ���چ	��6�)�՚���s��U�|��<�;�p�5y��X���z|,Ļ��!ҥĩ�ƽK��н�-:hPg�  ����AS���\e�Wz�|�R"i�c'o~�SŎrv%z�)��[�����}�;����C��xó�/8t���n������+y���͵���Tp�B �Եk�H�ݬv�qM0����ac�6�*.U�iL"VI�X&VC��[�ѽ��Zc�����v[�J"�F��;)VZ? �DUC�t�2CcZ���SJ�Ce�2�2UJ�T��de�4�\9~���xj��?ͥ�7�\�ڭ���W.�,Xo��Ϙ�
��7[����zʗ�H߂���0�a��-j�o����V#;��Zi.�6�)S,6��sd��ru�B��zt�ޗ�g.����
 �4���QP^���3��Y���3��ߚxW+�u���鑩���訚�,����B~X_�wr�qC>�/��̠8F6�'�R�ں�_�>�w5%��%�t0����Ζ�8Y�hk���[���{9iR���`���@���ܗv"Ú8��a������{y�6?cB���
��$�Js)VbQ��-�kM�x[��83.ǋ���L��eQI0ˊCXQª�`64ac�`6	�mmʶ����6��ӱ�6��Z��
cs�ֶgii-���@�7�(�)M���I�8WzE��9ʅ֑��ZKFiF��u��5��V�_O⒞�"s�G���WC]b���X��U�ۅ��E#S���NGo�D�3�N
3B�Ǆ��L�`Q�VF�8"��!�,���"���1���Ȓ�,�%��4*��1��V���A�&���vc���.<�ղ�!:����4��'3!�B��%�1"��e+�ۨ�땱6\~քi��J(`S�L��KgKl.���ڰ����m��6��Ū�n�L*�*����"��s�LoJ�&UT�V�4��Kը��ɭ8԰����0�S'�3�J8[���lM�dZJ%��(O��uR��ٶ'Vq.�7Tr/���u39�˅�R�7,��~\Oi�e�羚�c��ی*�z,.�bzi%s[�eAe���ƒ�]YXՙE-:��yG����V��QՁ�-�2��53$�^�c �GM����Y��s˷pe�n�'���85o=��m��j���5웺���d}�/]��yKY1r�zb͠ᬓ���CY3d,����6f*��au�����Ū��88l*˺�c|�v������r`�A��?Ŏ�G8w�����۽Gy�m�����+��`�>�{���p|�A�9͵���v�&��c3���\O<���d�����Џ��f�%4'�Q�3�����>¤�Gؕ�Ƴ�$��N��d��0$�'}�tbPd7F4�O��vT�7�mݶtlؕ�:-Ȫל��J�B�RZE׺]��{�5�GxS��i*��hZ@��\څӢv1�4���Ь^��:Ң^{Z��@ۘ����DU��G��y�V�*굠�n3�k�S( Z�OiX>-"��\��
/�[�t�{�+٠5�"[3+�+S�3�5�WH	���4L�=&���1^��ٰ3�z�"k��37��S{1/���1=�m|�i�ڔ���f.  a6��sq�]�}�fl�6�æ�R<���5�'nu���Hۦ-�)���Y�k�:����}�T��֫���
B*�(n�gN�xnY�Z_��r�f�B�k�T�Ӥ���"zL���?����i}��]%ѿL
����/���=�Uj�҇J!�������XK��^����/?��?װi_G�zdQ?͇��N�K�!ydw��८|�����Mr�lRڴ%��I�������F<�Z�䙄ɳ�,��k�C�����'<��G�,XL����g+�nER�~�7�":Q����j��Ӛ`���u�T6�%QLh7��.�D�J��z�j���O�����v�����P<��+��}��g���F���I�^�>���n�6R�[b��IT��t�j�,�hR}�c����`;>��7Z �79=o�ⷯ�+	Ξ��y�ehE� �꿣�����o�j���ȈQ���4�e��%�͘(���������)���<e�bEM3��v�&MKuT�<cm�9V5ߪ��#�fY�*��S~W-eNE��3f��;D�Ş��{����9�ϧF�� ܧc�3/�����+��Җt?���3r�L�O�����/�������@J���t�&�M�X�n����7�g�����t�<:��U�`Y߮��M��������fL��>Q.�5�ͧ�=#]C\,���4���� gkc��?�O{slL�������}��_=y5�\
��\W����yka,`n)��T��FO;}]����5_�F�@����aۚ�9c�C�(�V���l����C�WJ}kR�C�w�J�t��ӧ̻%��ģE^F���k�b'�r�%٩�V:��PW�W׬&���;��`���	v���� `mn`���QR�l^��f��� ���N�ϑ��k�Ĵ ��;��ږ��L�d�] ì}a�(�P&ۅ1;6me��3�d��/6�җ	>����D�@&:i����(k���3ڦZc�|���b�������^�s�NM=�/���>��4�	`�C�]��)�E�Q�v��R�H�;�jZ�^�Y���va�[�=d�cK�$��C�����M
4Άv�մ�w���	'=���0�a�_"{���ր�r��^���݀�����i�\�H:��%ߊ��u��(���ݑ���gr�+����9�Z��ޑ�s��9������+��=��ɶ���؟I�F��Gw�|�W._��׹}�6玜��\=~�kR��~�#>��1W����ɍϸr�&�o�����8x�2[�e���<x��[��r�N����u�mێ�k�I�o?���شc/��d��=���?��݇Ns��Un�����Nq��N���'.sH��ܩ�8/�w��Yn����378{�#N_����>GN�=�:¼��X�h�Wm�Ⱥ�[���ssa���[��%+�<}��ld�E,���k�p��'d��(��R��������D[/ʜj38�]�� s&!�Na��:�-���,���\y����̢S���ϘM�I��c�R7�RY�m4��a�'�"4e,�i��K�IQ�R*�R�4�����rSG��0��FHOFR�&�$:aQ�FP��0"b�h�ȸ�D�'Q~��2����%":�/u"�֞���@K��FRLgR�;|�&/�;ez�+y$���7a��N1}��߃��>���H����ՙ��Җ>Am*�:1n �R�1!m0Cc�34�##{3"�}�u����k<��F#��`8��&Э�2+E{�Qr��}X�o�|o8v�yԋ˦�4
s����zb�E�X�&�*��O@Ϸ�L[V�ܲ���.�䩚<���QB`~u�Z�n������=U��?�<�w���������=�;���T�ه���F��x��篿����C�^���|4W?�y��ti��s��ܐ>�+��B��4�3���HjՅ���7����o��||�Uک��G�{'�'����k\�L��c�,oAHYs��u"���t�|�<%��|m����FxV`�Z�gfsƬܭu�Tm�j���M�դ���˿{+���rR���׼y����>���2��'Ր�����I���-�|���\f�لg�cZ7���Z�q�8��h�z���N��Kn�e�����WF=)���E��茕(�Ӈkʍ�4�;j����#�PVÄ���t16a��=�\����8/��:2����o��-@["s�D��T��I�V�Ma�ܔ��l�k��A��Q�wT����5��&[N
��ѱ��2�i�[.ܝ�S��rB~s�Ȏ��ʷ��v�Iɔ�;��ɛA�IWnm�fD���=��&y����}]%�!gSc�L��`ECS�-uhYǂy���jMSΏJ`P]��qoV	�V��3����r~k*|5��h����R�h,�l�g����{�kR�c����܃���J�-C���j�D����m.R�Y��j�RC�[W���<�'�8���Aj]mW�� ��w�}��ɿH��ߥ��)�e��P�o�$��d"Ϧd*�f*sK�>s����doi���5��Z�c�D�X��[25˃ý�q}\� v,�z5dVnC�<�o�Pc���I�;����ցa�k�u�d����aN��v��4�ًa.^v󦯳�\���EW+;m>�ݗ>���wrc�_����P9ޅVd����J=7b\]h�#߅0S��5#�S�:S��:��~L�eZp��C���O&�1T�al@0�£Q?�4Wg�}��$�vOSj�0$�İ�"��˂�x��ciL�c2?*����2�!��239��Rh�D�ƙT%&�+1���,�4aal��cXò�(6Ⱦ���w�-��YS'����Ց��mс�Z�ͯ�������.��V�K�^Aό
zg6������d�]D�s���]ɢ�3ػd3�*Hh@VpY��M^pE�(��LaX� Bͣӫ��nD�g]�$�sf��-�C��v+�]�cb1�W�+�%=Ӛӱa1}�`X�v�jŠ<���֔'�1e��\�Š�H��<,�l�z��162���9_���\�����Z;Œ/��lLSoFu��uǩK$���%Ʌ�6�ϗ�gvz��'��%�Ma%�m<����D�:�m���hu��N�������� ~���r�&�����Q�[�'��1����� ���޳�|�^ƣ�%�:\½��Z_ ��[�&��yj�9�G�#�U���ֱt3N�pn���-�ܶh-&YK0L��S�B<2�����e��-�7g���-}��3�ϝI�R�TBӧ�:��9��IK�Of�d����Sg�(iu�ڋ��n���&+~y���P�h����!���$i Mc�Q9���})L�KFb?⣻�ן������_�~�Zt�v�S|�"����7�[x)��)�nNR|v��:�`� ��L���XVI@IS��Z��_�YS:TS���x�j�|���^Fˁc�|��އJA�<���뿚T���`䩾y8�������#�TOo�=��׹��R���?�m��/}8q����$�� ��T��/* ���F=�u([��nAM���ªA����ڸQ�����*���?�0g��:�$�y"Z�'�k_�Ok�}��� {β�:L*����d���Z�H�^U����4������ w�_N���z�T�^�������!�ߵk�����Ԡծ������/���m._���4�?���Zب���?��L�b��~��s�9�sbr$00�(A2*
��((�0�"*��,$�������z�=���=�������:W��T��D�`��}J>6��z����c�W�oA9QU]pLˡ�H�nnyzR#`OK'��lI�
@��ӣ��C�<�@s���=���:�RceO��	��SNd�m4�["�>/�r���^���];�r�m� �s�?�;���5�ϝ���^(��^1lv�`�[[����ŗ���B%5�O���;���>u���"yT
���!�$��D���DJx!�����u�@�G��]�oiL���yi��4��3�֑�����M<Wc�Y�6���k䗵]�qM��(��+5}����3$Ґ2G	j���? G9L6�oW��`�K�܉��O�{@
�4�˚�f�?�ߟR��q�d�&=�6uh��\��HO���Dr�J�������Er��P�'�J�}��q�3���Rk.w�����W��3=͕�Ger��\N<���Y�|:���5�L�e��	���1Hε���F��wu�� Z@�}/�4�?��~}~!�MgJX$�cb�&����
�M��bjT��¤�0����Hd$����ECH]��a��EP�G���D_?�{x0�Ӌ1~�^~<$�۸��EF31>����
ACC�#����ȴ��C(��0Aҍ��*!���1��P�KCR,S��$� 2��I�o��"y"9��YL+,f|e���XUEK�"�2�c	�KJx��#�V�����g�YTR�ʊj^/���F��ԗcf�o�ZF74�g)y�����9l�J��3i�]�8R�B�[�r\C���#�̕P7����S���3Ȱ�%V_�$�݂���^ R�.(����FS-�y����pͽ(p��'_e���0�'�ʟ�Dz�dP�O�g�����I�O���A�t	I�@.@�N`��?�Hς*b����I�@@��E�ev��3+`�;0{%<��㣞��wU��Ty�n�Ā��_�N /�r�;���Cgrj�k,Kl`�S,�CY�W�Ҍ�4
�����赛��_��3<{oĮ�V�Z���]�h�n����н�����еl�C�����l�:4�C߯�|�!'�r
���9������ԡ����Ǡe�}7c��fr<k9�y�6�l°��lĭy#��-_�'���o���!��(��_η�z�{}����o�:�{�'D��?&�ۇdȶ��>#�ߗd�F@��n|��eD4,%�nqUKH�]NF͋�W�@r�RR뗐�y�kȪ\A|�<�j�%��Y�+��qqe�	�}	�NocR�����6bP�9F���=�gT=ɩ��]�����=c�P�#���XMd7y���� /���֍I�Fq)��"Gin��4����^HU#ٍ��xǁ�0�
�S�C�Z'����o��Z�l���Y俣vj�<��S��G���_�z���}���a��D*���9���J�#��Bj��Tޭ��S7b0���}d+Ϯ|�o�_�����ʻj�w�ѳ���$q�����z���:��RM^%5�\�=%��ź�Sag��c�{���߿���k7>�v^��vRi(BW�x]Ž�#����N*��o_��^�;=~��y���?�Mr��'�`��}j.x.�%��6y��Wa���gW���itr�����xI��g؁J;zzy�jm���*����8�T߽b�8=3�3���N�JyAgʋ��ܡ��s+���o�T� ����K0�=�@u	`��?3���f/��4K��AMq�e��'�����î�<���Hg�
3�ދ�N>�v��򿩞���K��������"'!���ݷ��#Gӹ�
;+sl�͵�QS}-M��q%�U5�ZQh��[ޟ�ʵu��25��2�X\���9%|�Z'N�Z̹7�9�z��"������˨8j=uD����s���G5"e}S�uP��i
�:�Y�����)��n�FI�,}�?�}����UMG5��nJ'��)��������=]���q����z�~�����g#�`S�6���Șxc����T>��ϖ�˒r�_V̾99��Б�E4�>1�e������ܒ,Krͬ�h�@�TP�}hv󣗣}<���I��+��2��!0�Dyg�:�3Hޙ.��|��g�:G/�9zj��HO���;#i���wą`[K��m5�����.���v����]��N��'��=�*j���C�KwJ�����C��/r�|���Au@q��y{��E��/r��G�m��[��I� d��� ��O�?����4���$�'�۟t9�$Orܽd}$�����C�I��bx@(C��'p5�?�Y��<ӱ��uݘRۃ��Քx�g�L��I~�8��O�f����ڃ���K�:%��eU�a�xj�c�R��j��<�;7re��}x|�Pz�ѿ�NS��
��7�RZ�u��WU˲'�2}�:����ż6s!Yn!(�Ģ���U*����
 v�ˠ�TrK�c(
��22�>���2�>R�����u��-&�K��f>{�u&�L���,_�ﾴ�esf���YL�<��Feѓ��f�|r�;�W�ɻ��%-�y��J����Y�sS�Xc�ZS7^������Tu|�d,���0l9�Eo�����oچQ�^��|�Ͱ���8+�w�M�`2�$�����P֙�ܪ�0�}a-˶��c7���c��7�L[��	x�і���t�a�%M��0���D���{�Ǣ�a,��R�Ps��"��A�KV��m�\K�r�;0�GQ����������������;qhu�)��y+N=�b��K��oĨ�'ڲk��6nǢ�'�4~�y�O�n���w�>�ۀ^'�ކ���n¨�s�+�a��er��\Crv))y8�`���_6���{�ԗ�.=��Z��}S>����w�M��/��unb��5\�c��])�5�g����NZ
���2^�O�ݚ�����5�x7Er�?ܭ(SR,q��9&/_LBs���Ѝ�.=	��JH]oª��H��2�4P7�;Ͻ�[s�2����zv8{~�%����Ȼw]~������<���J�;K�ܫ?iM�qH/��z�t�)�B�s^���X=�®���q�|��|Mn����KZ�8Ŭ��-xjY5����6�B�TN������N��8��I������r���T��� wnp��)�%34O�$6��L��spJ)�@�1�Hk�u.(�3�#ޙ%��c�����n�${�Q��I���vθ
�(�K07'��Y��|���>K+S����V�'�ذT���ܩ�qƬ��Wd�B��0sg�Ύ2�5Y:Kr�(4q�@ϒ<�������� @�Ų_qsMEz����ZQbaC��5�z�d���inJ��!�:�6�h�M�lH�os��m)����!<>y?=ʍ����U�X�9i���ya' �bn$0f�Ye�=��t��&ؖ�(=^å�p󃾼�ӗɉ:�����:μV���t��;�\][ˍw�r��\�4�0)̈́��ڠ?=K9/�$}9G=}3��6	�(�z�2��e�H�6SJ:��,lJ��mM�mj��Zۡ뿫��<�P۱�|4���˱ۛ�e�C[�;�N�f]+Yv5���D�g3#��V�ć#¹����K��yi)����VHfb�;��9x��̅kw��]H�u Vޑh[b��H��9�Ҟ,s[�(�q�T`�H��#��T8�Qj�D��S��5Ξ���Uv�T+������6�~����퍏�ab!�r�_.���ȹ�iǎ�w�� X���n���8#��(��X'_���I��r�#�I`N NY�����
#�7�0� �=��
&^ 2M��Xҭ���\ ��͇
o_���,�u��L�1E���@jH(��䆄�K��8�C����m��Lϐh����,������1���)
��"<Y�a_��H�fۧ��w˗L>��={Я�;w�Gy͵�<��d�}�m�^���ռ��Y.��?(��1q,�<�^�/>x�]_|ɾ/���M��j;{6�ﯶpx�>6���ϯ�n}�8g�c��6.Yʦu���sKx빥���9^z�YV-X��<��y����E���J>^�*O��9��GL���T��WF>�܉�<l u�T5U�cP�Lis"�Sɯ�g�����*��H�)䭵R��M��+�r93��-~����Ya�ɫFN�����f���:dC�A��)�|���s�8�Y�1�zŤ�a2w�蠖����	̙	 �	�9
�9�ڣI5�ڴ�úU��3x��'� �)�9��a"�1�T �$f����<��C�t��i��;�A_�>�D'0���&����k>"@*i5�9�:(@y��c*����n�4wk�`��kt=���� ������k5�w�އ��% �$ �m'��ߺ������v�k5
��omA�y+���d���!ǫ�
]�&;~�q��V��G�D�t&����r��S0���L*2�9e�v�ML���Uwû�^k���rSY�<K�P�A���]`O����OQ��K������ܹyK
���]x!��B��֚��N����	)NQqo�߾��l'm�B��ĥl8�5���u�5������}[�̧�C]3���g�q�֓l�5�G���'�Wr������S��/��=��]����t\MYs�=�/,�3���θ��!K(;�N��Q���VB;��Ow�$�L��(�A���_&u�p�Ԧ�h����~��Z��U�>=����ԉ����	��v���`��Qdf	�8�U`���6�� �k�$ZY���K�Z�o~!.)��b�쌯�jv�"�Ќ`#;h}��`9w0�^��;K�����k��	KT�v���u)�U��wt&����-Y~�Λ�&�$I�jj���9�R���gmC��Qv��hM��=і���e[j!�b:m�G��Iֶ$�ې$k��l/�biJ����Jse��j)��%>��#Q��Y�~n��\���?u�O㱉�C��'f&F��=tp�,��F4D��=֐g{���띵���-i��j'f$���,����o�q�jx�7߯��{�������#y&۔��
���Q�I����BA�@���X�;���i���AY{3�֬+˪�����o����ۮ�}US����T3���V��Y?�o��ۛ\����^�e��:y�
`;���'���E�u�g�#��'��ґjF&Y�|W/�NN��|�՝���7��ƩEU|5%��Ce�X_{���h���I��#�@+K�彲1����o']��|
�
̓
rw��ᮩ}Y�[��qR	��r'�Ǜ��0����;(gyw<�=��q%�Õ(7g��<I�J��'3(�t��p����J�������CMq��Y�&&R!�dq\2�$G�O�W��^)1Q$FE�+�FfL8��r�@R���.<�ԨH�b��#<<���Xb�	&&:�ܬ"d�����(L�$#A�)�LL!'5�̄DM��r	q$
�E�u�EőM�\z`%	�dG�Q��Ake5�j:1���z��OI=UI���2��V>��#����Љ�<{w�~,|"���Y+d�,M
�v+�*�Tˈ��s�6��y���&p���2�i6���G�Б�Z�xW�L�TÔ
��hY��c��>c�}��|�c+��BV]�S�^ZˠnM�_�G�fZ����܇���c�I�{G�K0��=X�ʛ�.����/��8�У^��G�+Y����[��̄n���%~�8�?���a��X��!?b��4�Yf�wcP����5P �y?��b?�V#�	��ļ�g��|�e��k�ŵ���ߍQ��X8�հ�0v]��t�u
�^qu_
}�Q�^ǃt�4�{�>�1�s
�^�Emw�j�m�O�K����Y��X4~�M�M86o���s��n���V�v,�b(f�|T�G�F}�cдS��J*-C@�JzMz]�С���H�e�n;D
���6���E���\O��Mڽ2�����phX�c�ꉉ/�#(+���Ӱ��!���}"����nZ�,�÷���?��U���ZK�m�G�{La#_�8�����K^��/<lJ��O�46=�ߤ��m��6�m`ǭ�׹*��w�_!�����h1{K�+��il/���ĭ;O�lu�Ϋ���g�st/��ʒU�Y���\����V��Ȼs�:?�; 5�'���1���(V�=������Z:6�/�'+��t��r�AE��Uv�1�3���뻋\�$U�fR�{�yjRǹv��]�]h���z�������I]��cg�k�)��x,�їB�*6
�aZ�h��"��VP�[N�R�H��*(3WO\�=q���Y
dC#��4�j���3ñ���{Y���
i�[9}�܎7��yS�J9 V1a�Z��3�Xz�v`=M�	��G�!�љL7o�̭	�0�c��1��fK��#66��klA� a��9aRP��b!���" "0&�efJ����	6m��'��o}<^���>V��zt:�N���C�>v���Z�s��G
gy6**�����dH���lH�XzD2�Ɓ���h��o�՗���0�Ў5M��ʏ/�r�:M�>���`}#��ȱ)�l�ʲ F��P�bN��m��9�������HE�P�`�Ͼv�B'`�� PY���mj��v���k8����Q�3�R�i$��I-���-�L4�����m�*�����o�#����7�*72�"��RQ��Q ��PG�<�4=*�m�ΜO�j	f��~y������r/[��f7N/n��<[��#�6L�������"�^��T,,����VF8�Z��AptA��FD�/�����h�Ҥ���@����P�#�
	#8$���$BbR	���'8�� ����":��4���%=����"�ֵ��ǳd�cl��#~���_|�k/,�7^b�G�z������<.���*�{.��� <����`_�_^�@^G�ƻ�gӭ�����XrӓHM@KI$6%�X9vff&�ɉ$$E��)�#�M�!^���H%B��I� >;���,Q����L23H��%	 �$�
`ƒK��+����ړJIL$��q4ddR��JE|*��y�,�&-(���*>��4��?ɞ�bޔx|�<��N�;�E	���Y�=��$�T������_.q���Y��̨l�鋹?�)^�Χ�\��%��>�s��.]��7����#'���M���U��1g�+���§�'������{1�<l�G�_8iYt�<�����=�Ե�i���sfy����ؙ�S۵���Kj�X)`wr�\�*SSKY������pM��*j� j�r����Z�, ��[D������.�L��i;3#�qȳ|@�m�o���]�3�b�D�:�%���2j�'`t]�)�Z΢�,c����<����u݊�� ���<�^g0h>)@�t�B�a��2� �C����]�"t�O�K[�q�rl�_ź�j͢�_�p�o�GT�b�};f���rM�X�QR�*u����a�H�G�mv���>�ԡ���֠��j?Ÿ�C�j���z)69c���&&./�h��|0���44��ڮZ0 ��<�:P����5�sn���W*%~j�Ey�֤�Q��������	��0� �)����Ϭy���ǻ�UU���5���H�=����Q3j i�+H��e��sv��V���x6�#�Og�Q<���g�罏���Oh��
y�.�_�o>c��!�����ӽ���P��e��b��X��7cf��P���RDX�\�r��^��ǨF���f钧󿁼��gR-��_�,���\��f��g!����YI-�9���ĜgO��|U5�cI��z�Rsq��+hs;�Q�Gf1���Jd<���8�{iV,}C����P.E,����i�<g=�@�Ъ�V��Ts�g/�E��+�>�,�`YP�yE�*/�Pm�F��'��ZSU��X��@��K����$	��&�e�5a%9���J��7���8y��K��;	�������&�gC�r�l�D���@�#�f��9�9�fA+3#f?����sgO�ÙcL;�`Og<]l�Q�6��X[��F��A��>����h��=>���O��'C�vag^k�4���s��Z�̭׻q�]��͝ag_�ԋ�*V��"v�I`E�+�$:2�߆�4�9R�lM��)���������10A��f��oh�G��v�3Ф��=�v)PT.H�L50�	��M�@���F�J:MƦ:L�es=M�cm@g�I�j�W������;�ʻb*s�Q��~��g)�z���c`J� y��9N������g��pC�M7����ws���Z�җ;;q����Y_.�j`�c%��3�E��P�#��t�6&]�+��J{S��:ښ��!'�NH���@Z@P0Q��vE셇�&�~�X)���ё�rdD<!q$G���JFl��],��1�P-�4.#�G
��[Y��%�L.,�)&����|f6w<���v���{$s��{7r��1n�?ʷ�7�΂��l�Ƹ���̳s#3J���Ϩ�**`\IC3�����^=Y��0�v)f@Y���t/ȡ{I	���$$���@J\4	ѱ$�'i����Njv:�)�$$��B�T�S
ԥfe���KFV��%���Fj\�fQT�o�}�ث�Me��R@��һ���4חлS)=��|�r�, ��w+�'>ͮ�V�ӐPDlz!}{��������\���5���\��:g�̬�/���C)5�8�%.=����R�+@.���V>�h'����������:s�KWa��\؄�k:U6iR��ϮeWmޗrcnN6�Ɍ݇%Kf�v�2��y|�f9_��
_��*������S'0`fhG^�zV�����l�L]x-��S�g��jf��sba'�;��dJo
˞ �u6�_k͢��Ҩ�@P�ט6�@��5���f/ūy�h͡ʢ�0D`�y?��_bZ�>�y�1I_&�7]�lt��j� ˮ�1n܅I�^�;mB��L��K��A��׼�m@���I/A�A��t�)����_ OI������E�-�w\�.Eҋ���%zD R>]�t�3��Ĩ��ܭ5����WK�A��]�����~�ݢ��w�&�y�� ^�yoa^�����U���%߯|�q�v�&�k&C��^�A&�Y����=��EC�*�GA|�:�W���^x�5�[TÛ�7��vퟙ��W]��A�������r,(w�<�����d����x�'|�e1���>����d�zs��d�s��:1��Gf0zJ�«��=|P�ȫd�y� ����ϛز�@ ����zp��\�9���gq������L��4[k^��]ܗ��z2t�X6�=��{��q�ߚvI����c�)+��<{퀩h�;�?�v��{�=$��&>���K���Ω|���Z7�^�;S^�]Z�P�-���B�2��R�2�R1�	���g�(?k[�T)+�+;�FZ�{���n�hP��J�EEU�_�ć��YW�������4���#��4����de�q,:�A�D�;��A�-X��R�iqr%F~�&�ܰH&�ȬAcxl�8��#�F3�e ��b��I<2�a���C���B���y
�<H��+�)����<�OR�*k޷'�0}�CD�y��d!�'�ja���)���x	��Ӛ���7�E�xu�ީ�C��v _>��c�z̫��	|��3�W����R�~� �a�{}��F��-a��^2�Y@ŕ�Q�
����9����Yik���'�� l-p�����Y�iS3�$��؉��β���P��rLޕ����Y�L�X���Z��i�NԲ����zD
��"H�1��"�o�&#������,u����u�XSjgF��	��me��)�<]���zG���³��^S
{îAptw����V.�ى�T�~t,��yoH<���x�]-I��34!��7#u���t�" X*�m�)�UtD41�p����I3:2�U�׀(.2�؈HB�C���'V�.6,���rC�)�N�2:��E
�UR��i�LN�b���?"�n��t�u�����{|��|��>x�)^Z:��?x����dh�JRc蝑���������ɘ�,���2�������gJQ1K��b�ތo(adU�j�ZS)�P/&�jaH��t*�Ћ#1<V`O@-)���,������,u��?�t9fvV.yY��S�Z@jl
9�>16
{[#�#�������W?��3�l����8��zY��{�����yg�r>5L+�䣖��Z��+�]���'*&[ .�r�~��LJ��np��}nH�yEV=6�EB�c�"��ŕ��i��l���������*��x�۲�ߤ�}A�MIG��j�I��'��Aw�">�=�����~�����S'�������|w�8o|�o����Nq�����^�������w<`�|/VdIey��W(O����q�0�=O���_�B�p�;�}3�{�U2ߖ/����Ǵ�j��A�w�,���y��@@�f�G������?�����5
Un¬z#M;p��)�u�aR�*z�/k����Ǣ�^����*�C�<���0Κ��FU>��� Ө���7�	��z�O!OY�:tߋe�����a������m�r�b������>�a�׽�M�ڠ��jP��?�g�+t߇I�A�z�¨�����+��6���gQ�ۜ��&ג��Jii,]��>���_��K��-~��Җ<b:"�)��>�u���ទ�O^��ϵ����9s�)�� ����*�ۧ�e5��}�f{߾��ڏ��H�K^R���ߝ�w_��_�p��[��F#O.����k�p ����噗��wf2��/c踎<4�/��{��۷k�R��Ԁ�+���6ole��j~Sˏ��p��8�]ño���ŉܺ?I@n4��>M�o
�}?��?��55�B�o�U��Q��T�T����nR��#�w&ՙ�_~���9�U�=���ϗBNPui�s��~|��^�
�a_�FYK"6IQ8�*K^%�R#w�ڌ[N��O�(0Cgm�m���&����`b���&R�[�
ؙhsSe]��U�W�@?~d!��])`7�}-8�:���qv���8{�<������^�D����@B���
,^ދ��������j��ꉇ&��9,|lON��S�a�C�Ȩ�̝��f>��E/���7�J/!��R��t{W2�\5�����^
BlbB�X�`Ǐ�c���R a�Q$G���n#�����Kc=�,��w#�ݒ���̩������;����jn|�>�Ʌ�,�saB�)��G�iRg�/��W���Q�6	�|=A�e"����q��f.�֙�ϔ�s\2E�j�/Y3?͔i��գ���ή:*\��`I��!�̌ cC�͵�o7cS�����hՄn.`g�3ɳ�`���5v�vZx0KC+l�l�u�J�:sM�����G�����Z�cc����M�
gL�������F�٘Q�lC�����8���لZ79KZ1"В�~F����� �ni�o���Ӂ����Ey\^]ȝ��a[�����!8"���!���g���eB"��=ywH���f��<f�y��Ɣ�U�v���Pk�v05��˅�� B#�		%2$��(bã���JMHҤ`/Q OIA_�R~BC�2�Nͥ0"�<
���G��5��ԆGRL��%>为���Jy�/%>��S-���J�+)�Q�@� VnTI�r��n�����C��;q�F��?er�5II��SUSh*MY9�/.��t�23��ɡ.;�.����ݧ��M]��PK~r&I���$呐�E�@\BJ*�I�.Q�.)�?(=)�\)8�2��)))!;;S��)�!̞1���.�M��q���b��_����9|�36mZ͑��g�Q����P����;�"�����Խs{�5����+R�(�y���~��w���cO�XٙA�uX�&_�_B��tb}܈	d�s���n��=�G~�g�n�wֳ��yg͇�8���Lҭ}X�w4g�}��J�%��[\ʣӧ�h�2V���^ZɊW^�E�?���,a	/���1�@ ��Ђ�N���[t�ϦHg���\N���y��pr1\�Xd��R�X��� �x����v�Q̇��b�	�ì�0f=�¬�e���0�iܺ��i��`�S�'���͜��Ơe?���<�٠��\�來��sm䮮�!t]�DW*�f���H������T?�.jٶQ N@��_����=8U3o���kޅM囒�S���ƶ�'��ۉe�^,Zj#uUB��m ��ko�}P�yY���S��u߃i�MF��!o�y�]6���3:oB�~� ����T�q�Z��ڲ�%����/���Ɠ���yum&_Ӆo/����}8�]��j�~��ɳ�0������ElI"�	�g��(����o
�H�zK�?W�������pe�S�v������� O��9LV�2�����#oq��Ra��8��L&ͫ$�>��?͏�����4���'ߜ�G�i�[�"f>:��7p�
��g�H��7���&o��=��>R���-|w~4�όb��>��n8�������z�NnN/���8Op��AIE���V�E�)<S����M�P���M��(?v���4�-��{)�דs��$��S����1wyWFL�d����:�4�CҰO��!��Ϡr(� �s��bl�Vn���6Ύx����A�H_dd������(��ي�Ԁ���"���*�׵2�/����,�*fy��Ob�Sꙓ\M�}Iv>��y�l$pb�G��?]ρ���7s�@�U�6�ͭ���%Z
J�>"�͍)�"\=�~@V�x�8S�]ƂY�ѐW����1�!E֧ۺ���p2�@bx ˟{��'
�}͉�6��P/|ݬ5�s�7��� ksR� )��=B�Y�-�!�:&d���tw6��M���Z֏�gb�9ӓ�X�)�O��rxa2��^������7׶��m�} *�??�t>�÷����c�z(��[|Y�ٍ��,ȳ�,FFX�lGws�M�r3��Ř[}��:i�G��>VFcJ&��Yh(�&s՜���K[gaN���G�+����v4#_�-�ր/9��)]܍��O?3�X2&Ҏ	qR�92!ɚ��6<�n��'^(taU�+/ر�ʙ�:��qp0�%���.,/���r��A2��#��w�ǝø�Q#gV��gf����>R)XX�O/we��T�����91�z��y�;�*��`���;�!>"?�:Nx@a~�DGh�׮��M��1�D	F
�= �4;!AY������}�h��..�GG����'�Ǜ$'G����<���&�ǝ\w��}Hts"��Y�����ȉ��1d�ES��A��BJR��M� ��(5�ʌt� ��Q*�PaJ�6��H�<-���Q��ir�Y�Qd�Dj�6�
��1�gW��AQV>	1ID���2��MLN� �Ai�'P���FfZyY����r�r)*ȗ{�Kj��J�ztd��F�g�*�M�ͳO�`��xa��|��3Lh��Z�ytY=�|�f�����Hm�RJ2r��,J͡"�X�Q J-gh�!Ft�A�<�7g�a���5##ė5�����sY�%$�Q��Cir�2��t�"�->G�� n���oА����9�WTW즓��A�@_I�

�����'*6���h�"|	���T߂��"fO�E�d�\x>8[���ϼ"�A1]� �9�X&%� ��i<l�z�QLU� ����)7#^=?Ƕx%����{ǁG��z}�ksc3ռ�F�*�*�ӡe�����m�=�&�-' �`5���ļ�y�T�m�%O�0�q\ ��z}�Ao����@�&��E��T�����N���j,4W-}��4h9e�3m:�!�}�a���w�%�'�ڸK�A��tm�;]���5|� OW!`[��y�e�a���%/�����t����Q��a8�Ǐ���Z9w�̵[M\�m?�{��=ͷ?>Ç_�a�[C���3ǕRѫ��;�p���B{��?��~������y�������c
�A��~���p���������@��Lg���dw���O���%��I�^�����x����������㷸z�w���2���o?�c�*�lƞC�8z�?�6���`����y_Ξ���c�|���7[�~�����s��<I���,7�'���{�_��?���M�!���O���9�m��K���S��򏤑�L
�w�8*/h'�rBhՍ��=��M�Nj�
씿<%;���<��t�n�X�i�:R��ne��K��7�Q�.�Ǝ:;j,���H���c��d���ɩgIH
�5䩬b�]|��t�����C�7��C@��ΙpO2�l�k���Pz�;;��H���6��U@�EO���1A6V���W�pqƶ�AN>L9�.��u0�FӦXٓj�@���6��@
}�<��%.ț��=ɱ�{4�ۻ{+ݻ��jo�����4�(p�h8����J�ʝ|-x�ʟǋ�Ӂ�Ƥs�S��mR��L�˅U,.vf����a�<U���c947�s+����r.�ו����`�@�n�9(���87���qm�`.|�Ĺ��8���cs�80%�=c������;oV;�Z���e[27ՄY�FL�7`R�!c��m��H3�ʹ�
4e��	C��fɰ3�߈A�&�~p����ϸ(&D�0#Μ�)��M�dq���-YQd�+�X[i�{�6|�`���l��Ʀ>n|��ͮaA����r�����h�>���ݯ/Wp����؛;_���>s-��/�5������l��w�8����S�x�W(�5���|n|Л�5�nx4�Ý�W�*�O�s#�,M��p���� �B4H�	#<H /0H��пI��G�!���H5ת�l�Q"/�G{0:/��h_<u$�YQ�Ey�?u�TE���Bf������?:���R�C]�U�ɘ��Lm�̬!M��������̝����E=yrb�����0qT?F�odp�N�4Vӫ�D��֣�����248̊��F��
���г4���w��:R���"�JL��� OY�ڕ�����33���L'3'S (���,r�ia�]^���ІLFw/bTc>���2e@93�T0{t-O���K�ZY�A��+%~�dڸQ��Gip��J��V�K�P�@�����9yP��O��psl
e^�MJ�wt<�6������G���6�ZY�s=)���#��.~��{S�EKr]�"��RV�A����N��Ɔ&���ӵSW�w�III)�e�t�mm=l�3��E�s'<���&{�&��ԑ²95d&G��;=�#K�"Xj��b�x&�6�T�,n���|��ä�� �ql�}���x�ۍM�{�Ʃ�&�������)�Q�c���;��{�����0My��W��x�n�1h>�Nd���}��A^����{����4ƽ� ��s�ּ�Dxz�'�����j.`�K|���q�[����ª����ޯ���u�D�m���e�c����@P�׽�T�D��mvٌa׍���:��C�'�uz ��>}�Y(�*�J�ǹ`*��uw̤s���g�K�<܅S����_;s�~').�Ia9��w���ܼ;��#�H�s���'Zپo�^>�J^���*��R��/�v�{pRi�������joݿ'B�7'ϱy�[���2�}?��Ou�r`>9Raх�~�͞��xr^��.g��G<.����͵��i���>y���_nZ����wPA^7~�:��?	�o&r���\�1���"�����y/J�i))�R'���=����M����M��ҥ+|���;wN�|��m��M�8���ݽyC�u�<�݇O%��3>�9��,#CqL��>=O@/�|wYy�;?s)t^nX`���*{cd4��.x��3fZD/'f�ZA]a'�(�eAd2s�x��x>(�ʋ��x�)�J��;!:�i�2�l��3�ZVA��Z��y�o�:�3����R�ҵc�2�gw���Ck��t-̡�$�Q=(��t���VXn쬹�H�`��q�(邯Έ(ɰ�$�O���F׶A��y��:�C�X��)N����=ɾ=�4��tu���KS}���,��r�r<ܨ�0��
V6�2:ޘ�]�8�Zw�j�ޖ\��/[�&�P��rs��l�Y����l�ɉgR�qE%���ĵ{rgc_n���m���o0�������(\�0�BÎ��^߇�k��J-����˂B�=�ǱiI|=!��##�24���4��/���o_�F�y�>0z�����C95��k��x��'ow��ݞ��#�w����%�O���Y?Ic`(�FE�%�}T�&Dsrf2�>��ͅE9��4�+��sgU%�VWq���(��O`��m��6���twʺݭ���ʭ�}n�rk�@����sO�ϥ�zrr^9�'�V� ٰA��Oqim�YV�G#��D����U����Wks|<����$ ؗ��>yʚ��r�R� �)���S}��d���6i�Mb���Z
�*!����%��/��������^[�������aoH��-š�tJ��{�+��d�vv3��fË����<�HƸk�2���=�,��ƕ��d)[?X��uK������B֬���sx��9,�7�y��婙�yl�`fNĘ����ːs����������S�OϊB�w���P�.>���D�+)%�Oȋ�K���ed���_�h2��2)..��$��x�2��?��#jY�Pg捬e��:Q���c��Z�S����L钥��5�'�S��/H�C[��I��;��~^%R�+qq��݃:�L�{��՝|Gg��ȶw����Zo?�\]ȓ|��Փj��Gkqd뽃�I���Au`4��!t��|&ZX�lgO��/1����=�N4w��˞g���VW3��1Z�mvY!��NZ�wS'-p�`H��w]L�x.(�c�s詗�W���1�9�1��$���c�X:�Q�a����|�q,���v�I<[�`U�����6|�u߶~r�_��u��U?9�>���h���1�_�]�<tA����Ǡb=F�N���дq#FyϢ���^�Zm@�r��|ҩ�x
��}T�����$���)G��y�a����ob׼3���~�{��{�,�i�[9C>���5j�/�ۭI��3�s S�A��E��5�.@ڼ��m�v�U�o��s�:o���3P�W�]���G��w0�z۪�.�NDF=yR�t�c��P^}%�S�p�\+��֏;���y�3wn��ޝ>ܾ�U���@W)K;II[ϕ�}��{���!���2�S����J��O�S��;����U^�oɵ���*�����^�[_=IÈ��������ّ��>α��xhF�?�ȡo�1uN1O.�͊W��_Oi�A�� ��_��m;�d�[��rZ��ᇫ���� ��\�6U �nޘ&j,��M���ɍY'i���іr[�������q5Тm�}�?����[��o��"vm�?a��8�����8w����I/�OT:E]2)hL# /��*�*�ݵ	��
�
��H�<FY�\q��etr*ϥf�"9�q�dYSb`ǚ�46�E�O
[�����G�,M/竑3y3���>a��87o����b�j��ʘ�����o�>t�֍��:Z��hm�N�n��ף��N�z������̋�=ɻ�-�6?{��n.�gg�A�Ժ�OMv)�z���[{)8���!J2�@#Cm0�r��#׹ჵ����\���]4Ԕ���3�V�XYY��䀃�)�v��6些�P�=���J��Ru�|6�{�Fr����ɯ/�N���u�P��Z3<Ç]�X?8�m�dp`~?�������y�@
U_=�"����sX /���S}���{R����č����E+W6����-���|��:~_U�����Z.,�|���:�ӢR-j�r,���|~\T(���b�%E�����/�sae%��Zͥ��4���O����^\�| W���1�>(�{r
|;�̄����\/̗�s�]����Y��C���Z?���'ܲ���_5sw������������,���$�<��{CYP��Si�,������=��N#?����!��s��`I�N O�vr�]�|=����%8,���0BBB4�S�g#��Q��W�ƋR��'P� :<���B�B�Iuct�F�Q�i@��>��:Bmu�Z��q�sNݒ�H�1$�֜"?����u�g�;�(���/s��'������_N|Ư'?秣���N~=���Ω}s��Nt��  ��IDAT���#�ֱ�{l�l��J����y|��b��h%/-y�����K-e�f� �+�������U@��r�w|B1�{񤤤h}�ғRHNLҔ��$���Mrj��ʲ׵���iat�r���Y��ay,U��+yiJ��k5�<��5Ӻ0�4�G��%o���ֆt� �<Isq"�Ί8se���D�|{I6�r�;�4՚�Cm�	����D���VfZw�T'wҜ��r�!�Ƀl7O2���rv%�͍Xg��<�ӝD{[���I�
�r��섟����裏2`� ���Ì�S���D&�b&@jk錵N��8sIG�*cs�J�@�d�?�<�:��9�%���������d�-�w���
�5֚i�[a8���S����袧����#��=�����8��p�]�+����ƪ�#t9���{��O1h9���im[��wы� �V��Ҭg:�~�5�-=�`�!7P
�=uT�!�bŰ�9��0i���-8�ϥC�`���9@]�^�WY�l�ƦE��#�އ帇�c+�k���j��m�k�=7c�C���FL�uڀi���ߛ�P�]� ^�����EW�F���*��{�8��;i��nՑL������w�8�M#�.�ƍm�;�-	Ԩy��  M\�ۅK�%_��)wn��5]�������������1�]5�~?��n~PV<�w����ǻs���`���R7f}f?Fv������;�������({�-��#Utӑ7?�ƞ��x��I�^0�GwJv�AȻ�O��c��ٴ��-�*8�]?��C9w�/�_����C�AWo<"j&�e���)B�˸y�sI㪐c��j��K�3����W�k j�
}���|��'lٲ�˗�jM����y�oܒ�*4~�>/��٥y���Ѧq��q2�U�t�|�W4��Q /?��t͟���G�LG��\
��*���=�:C�$S[l��;���ȋ�z�l���/��k�l��70�#�¤|"B����I��gS���ƍA��/��θyx��卓d���vظ�cbm���+��ϝ��]�г�y��e|��JJ32��|�^Bh>R{��` %@ڿ��Yt*�!D2�D+�5)ȋV�.�����ߟ����G�p��=s��[7ҩ��@o��1�0�Bdgc���	���[��nAK�9o�K��
WF�Q���\�d �O�\0�܍��D�X�9���O6ґ�`FK�-�r�e��MLd��9]Z�ϯVr��:X'𳾗��ʍ�Q��s���\y�������ye�<�� �ʫ. uA���gڠ�W��_��Ot)�	 ����rn�̀�Z����d���;<������d[����~�%�Ζ��q.�]yN^|9�M��}^�GYЗs�������-���E���un6�OM�Ɓ1\������v��n�I�o����oWp�jN>���9i�·äp�ʔ\wZ�M؁����������5���
��R�hK����y�zڨ_y~ʊ�O� |Hx�y���Bރ
�� 42J�<լ#���v����OA�Q�$J��9u��s#ס	�KB\H�� �F����nT�8P�eF}�c+�Z�L��0FU&�v�P�۾���>�֯{���^�_8 ��0���¹�\���>Ε_����������?���Om��ѯ8s|��n�â�_q��g�=�9�6���_�מgͪ��Z���S�RZTMea��k�UN]z	%I��'g�/@� /C*y
�2U��(5])�Ԕl�RՈ��	Wd��lc�;OO��)��ʢY,�ϋ��¸r�W�rb5+&T0 ˓�U�ZoJl��p��S -g}\��.yF���̭�!0��хFYW/�
K+
��(�2[-
I��&�T��P�gO���̭�5lS'3;��q:K~�[���݃fW�����5q���[�j����GEE�zt��%���/�g.y��=�zV�^���i��e��-�}b��o�y�K���R� ^��ebb/�+��g�W8�?��H1�yfCOi���IE�/���ս�M�>���t}�Z�ӡ˗��ϲ�EtY���6�-�0��.4G�j�}T������t��X	Z7�F�w�5ϸ����5�M���������V O��1����ί;����ۖ=ڠ%vM�ZVp�5���� OO���S�,��mD��@�\�a�O�F��|�i�g��w�����G�\���E��oСt�_Īh.c4�+(L����F��~]?�ԓoN
�	Oܼ=B�f47���uFqC~�f�h ������;{�ܾ���R���Ԫ�{�����b��7T������A����m�x[�
-{M �?_�΂w>%������.�BdM3!���/.�����|i<�}����g��^�]9���0��|}p��������]l�j&;�6��H9��6��������ޥA�xk�������!L�⭑�~w��-���r3�����Cm{��<5rDMꁫѴ��v���?vJ���_Bޭ�Z����9�1�>�������C�<4�Ԫ|skpϫĽPy�.�5� �,��� �cemF��;����͇1*��:Kf�ر�Жw��x���u:#֚;�4��=���Ό���:�'f���勗���x�͗��P���r��
��1�y{���DFA6~���j��:+$Г9�?��g�����d�a��zz�$5���H��1�n눒�6�ڎGgR�m���jp�*�� ���4>��=~�����S+���愭�-f�fXZ�Km�L2�?���Ht���S�ŝ"Y7$�Y)������W�r����������%�G�L� 2"�ЈX#C
������.A����������siU	���p��fm$�]�{t��M��/�r����}Y�I�����n�x�\��<ϝ����n������+2Y�K����.�6�-�d~C~ߔ�n4�Y)/��5ɶwDwe��2���v��"��˒����en�{Q�-��w�����D����Or��OM��Y)o|؝{�ؽۓ[ou�ʫ���r?�P��g��?3�=�X?0�ÙT�M�H'r�u�:�x8݂]Odsu]w�no��OZ8<���������K O�Q�T������!��+�kS�����"�C		�}D~~>�o�f��s
q�"̉� w:z�kV���4f�d�Y���\�^ɲ�4��̒�<7��5���_5��~  /Pw��|��$�� �Xu1Q�w�&}[�sW�$��{���U�R��ĵ��t��\�Q�� �_�}�g�ݐtn���oG���Q~�n;�On��}���UL��(�{�SQg�2���Iiriy$�)�K�oLY����`/%���T͟^Rb�5/Sk��MK� �g�/���u���!),���ޒ��X>�X��'V�hBGgz�Sψ���lͯ瓰Lֹų38�}a9��d�__�F��)��>	�Le{@2�e�mA)|��^�l�I�ˀ46�%����sOd�{
[<�d�$sY�Jb�_:�C3��̞��E��{v'~H��tV�7Q��xz���˰a�xv�|���	�񣱾�B��,K��"�Sȡ�r��`�W/:����8v>���I��w�`�y ��J���JT�SZ�<ǁ��(��z��� ۦ/p+��q@O�z�Q����5G���k���+~	㌹��?�C�b{�ƾ��?�nŲ�~��U9/v�#@X�������4��>�y���1|�Y5r��������d;]�#�ϻ��W�B���G=&���>`�6xD5�*)'��}��e*Ъ���{�ưQ����]��y�_bR�	���0�ڀA��^y�T3�~���*�BW��@�k���A�j��y�����%s8���e�Q��ʴ�A|�>��g8�]w�\��3L���Z����Ɗ�K�6�����7N��Rq�|�me�XA&mY�{5�}Dlk�&IF�n\���b���O OK��!�+�7��a����8K�#����>D���9�/�4� �n0�È��L����O㔱|���ַ�Ȼ���6���	��U�ׇ�8}�+?�4@=e����0~�;��w&r��.��o������\��Yn�� y���A�l��B��C�� �8��u��k��7T�͊��vj��C�6�����ڕ��ta�L������<��O���sR!.��(!*�y�9�%%K�W��>^<��2�`ƛ9�#0�Qg�3k�Y�����۳^ߒwl�Y��϶1�x5��Ѯ�tLH 5'�ԄB}���ϲe�h��DEZ��� K�ٹk#�u��7vb�h)|��@����:/7���yxL�=9�ܤD<l���%��/���fO�MC~ş���kllI�s�b��Ѥ�C�������������W9��9��o��n9:�bkg���5��X��le���1.V�����l_ƫ]����c۴T.��L����;G'pnQ=�{0�р2�M�����:ꂌ���3��xc��ˤd���̒b~^U��7j��Q7n�~k�ԠI�������g�,i���粌{�^ঀ�u�_��|۲�ލ/q�֫\�]�_��<W//���^`S��.m�yI���U��V��*�xG@��J9�
���_�»�^֖�6�U?�{
Wp��b��(���nO�9��z�ƽOzi�ȿ�X�/+j�vq���kV_NM�ݡ!v>�-���dz��i�zc�"�}��㵁�|�J'Io(7�������p�l�xW��US�j��6P�gIP��6�"0�_SPP�	y
���)�S�LX�������D�NcV}��(�#Eޗ,7S�E�)Y�c�#�̒�0^Ց��Ĳ~y�4����f�~.wTޕsr/�B���I�3W%�qWu~F�-`'�v��^m��5�h�HU�%'j��Q`(iݾ������{9yz3l�_�_�hJ3�ɏN�0:���mD�r�S$�)�1
��c%��H�����	�JX�@`��(���5 �G[bxzP"�e�i���䕲lB	K�V2J o��#_��md>?�s�>�3Q��� �E������y�D����27�d�v��*0��l��O"�x����T.z�k�߽�d��o{
��t7���	�\���O��l�J�hG/��p�Jdiq	��ͣ��4551��'X�`u|�I��W�g���46
�����.~<o��ަ��x�9��C�Y0�C+��5�Ȫy�݊��#X���܌X����1�y��QM]��uޓU�-����uߌ.{��'�N}���B���.�Y���χ�vۇe�o�hjĩ.p:�\̽�Ћ�E�*�o�k�)l�F�j��r��]���d]�r�~{���6"��!|�6�AA�E��B���y*��
QfR�%f՛1��\�n=e��u�W|@���ykГ���3(X�q�J�r_�2w1�Y��+CBa2s��T#y�c�l�ґ3�v���-�]����\�-��qK8BIu��}o�䁓䛜&��*�?hE�*�۝!��^��r��Z��)&��L
YD*b���^�w�'{�ܿ!9��ʹf��FL�e�St�0J�����B�;u��{'bKK�)�MZ5��U�v�J@}=����CZ�����ܗl�4�]{*9p8�3g����f~:�ʅ+C�q��0�]΅-r���IM�ޝWl�șJm���WLm7�oR7@=�_���O�g�Ξ�N{�jRN�/�~�BY���V=���S�e�˱Uj�o}5���c����(��+#�̎��Kf��Q�a���CrV�����1�����3O����'��&�	��L�fi�R3�qra���[񾽗���!�X�X�HG?�T�?+���H|\��(a��%�)p355��љ��z�k�{�&�Jil�5���'k#�TӮ��53&g����dgbcdL���&o����hf��A��j�LI�S��b�@�������DA�j�U�<�{�O�ľ��q��q(�0�V��ٚakm����ak������)�����W�bM�d��Μ}^���7��q��P��@�y��l2_=�ǼD+�9�Hwl�e.�W��+ ��oŠ_�W��J�46M*f��\�=�ǹ�K8�J�|��>k���4qZ����s�s�c�\$�T��j6UZ.zA^��"���K5ݹ�h����Hdi����#�{w�dt�qSҺuGY"Hޖ����+iޒ嫲NY
/���bυ�*�
�=	�`��������'W?�ʕ���mU5�/.�g��=3��FF�b��w���P�g��%ҎT�6�j���΀dSs�lt����ɹ���4H��d9�4~|���O���!a�N:=��#��8�$�@p�?�!�k��+)+���@0$��H�7/T@&���Dz��PW�Hv�'��a��%P�O�|/�uMU�I�������CǨp�T��pe(}Rܙ�%�����/^�ҙ��z����`L���pr�e�0��/��S�VU��^�T�}�_���(�p�Gͱ���ͷ�r�����9x��7���5������˴MaN5q�1$Fҭ��~����P����_�OYq5%%T�h�OK'):Z��C�ꓧ��Vg'3�&�)��%z�_
��`��L�<T��KX>��E��Y2��aq�<al��8�
p�s	�s �l�8���q� ���rH~u�〕��|8�������΅�xN;s��G я3.��N�rB��8���!��O��瘕�Xq�7�ީ��wb�G(��"(�w"�ʆP����������;9j�����<h:	Iit02���+�!�L��q�J�����"R91h"��Z������9�PV��3<���N�c?p�6բ�)l�|�Y��'�������G9��0m؄e���Nk��e.�(F /n�1��E�������8�ҷ1Rּ�5���H /B`г/&a�n�T�$]�~_�1��6�C�dQ�Y�� �K�3k��k2�{L伵����t�Ä'��[�s���)�xJʅ�_����h�F���#�E�)tَQ��W�Y�+?�{�J����"���bX�
y/`��<f9*�ٳ�gN�;k)%��w̢kg_�.Ngێ
����]\�>�+�{q�F/���K�7E�ʊ�|�N��o���T._�|���:�}�ԩJY{H2��#���I}��X����-meXR �F~���6��.y�5�z���J�����<�r�Ͼ�'���%���,yc:o}2��1�4)�~Dg�����9���|��c��]Z��� ��}9���*8x,��v�K�9��߮�p�v��k3�޼9HNh�d��v�%~��+IH���y���P��|������?k]����e�]]�Ãm��g޿wR}�k7�hր�/-$ ˖�O��S�J��=���R<
�4��b���U�SZz
t�h���I_�{���+�+���
�}`���F�l6�a�d�K�4d2og�2�3�ڔ4��	�����^
�^z~!}��bok����j�Q��|)P�s2(�ޫIj`yt�ы��
-f���#sgO���5T�c)��1�
*����g�%�B��xS�m�Qs
�;���Ԅ ���@�@5A���i�����\��Xj�l5ȳ����_�/6t	1gA7��(����,*�`�h~��̍�c�3�������x3:yv ��X�ӧ�U(9���6F����bϐTve͠6NIc��y�����+5�����u�ҧr����{(����葱�>1�[�������l�E 𗧹^��,_�M�w���鲜��%�os����S���	�}��O͐t�F+�~l
7M������kw����ù��P�}8��o����=�qU%g�rt^��d�������1v#��|x�ދ1����RfE��	a:�6���:}��m������F��}6�>�������������@�����_5���X�p�ךZ���)jּ`hp'R���^�~@h�������N��xZK(K�&�ےJJ���rw��Ɯh'��(v#�ΔkҼ)�mK�L�q1�{b #K��)�G5��1�^^~��\���`�g_�{�Q��:��'9v��?�_��sx��l��_�_�����������s�X���_��y_d�#�2��<���N����WP@VVyYE�Ʀ�GqR2}�j�ө�Net%�t��Va~6��Mt�ؑ^��4UTѩ�H��'��j}�Tӭꓗ-�yMn*C�ٚ���$��-R����9,���1����aP�)����j�~q���qG�q�e������:/�9�
��i�>�sㄻ/'=���9.pw�1��]�9���IGwN��q�U�w���󵝇ȋ�
�,����U�,��I��T"RM��~x!R!�U���j�=�|����M=���*�uMey%�H����CcK�M��0o��#y�s�I��+�7.���l���f��wbD�@«_�~�,��x;�y_����n=�I�M�կáj-M��v`'0��S��F\p���ykO`%p���=��ź��j�Ų�X��h<�Y����މC���X��E�0��1&}w`>� *҆I�#���rJ���_�F�>(��^�q9�#Xtۆ.}9��%�V���U�:�f��<�����)�k�6�ۊa�\_��*?�C��w�6�bՂ����V��U�{�c���܅X�<�M�h<�ZH(l$�(�n��,^��W[�8t���~k�@��;=�t���7���Gs��~z��V��r}��yRl����Z�I���׮%�)��Ze����<�
���i���W~�ˮ-��g ����L�G��:��c��3sn$��ȡ�o2��ь~�7�G53p�h�nߢݛ ����9;�����z�}S�o��s� ޭz.�������Qz��)sծ~��~��6�n��~���_4��ׇ�v��A��xʢ��w��V]����#�Sӿ��a�޽��[WQC��\�m@&Rc�H��!����;[Y�Jq�-���y���/�]X�uup�/^�
�#G*u���LXbf���Yo`�:��;��d��2*�7�	>�i`����B������^�ʅ�U��t}{u���XZѧO_ƌ{���B2�6z8��T�����s�(���䅇��Ȕ��ܵ����فX)���=�OH�I��]N���_,yI�Ŋ�-,H�k*�, /=�̔�]�����C����je�ӂ�+K��g/����^�6�H�^ḧaۤ<-����|���+�v��czs���h>���x;F�[Q�dC��)�r]&"{*�� N����t�s`T���}X�;��%�eB['�q�1���
��2~]^��W:s�n�\ۃ[�6q瓾��П{����ù��(��o���C`�P�	��3�{����Frw�Hnom�F�FY��@n���}��fo.���/�����.��[R��g:r��">���i옘��1q|<,������g8�k��)fT��3���%/��xW�q1Qa��B��غV:<�;�lN��!��Ƭ�	���t������C��f��F�ې!�N�Nq��Q��S��lM�quj���$�`?տ.�/ּv�k��]�/aA���㏟�����%�32;�4}r\��FM��6�R���ވ�p/��v�#\(�xwБmeF����Q�K�{�?���L�âQM<3�O��#��3u�$��:��3�l�<V�[���cՂ�������^�,/>�K��ɲ9�X��4��:���L��S�=}"���у=�/}أ+#�tgXsw
��݋-�ںAM�hj��sm�6�Hu�P���R(���!#���R�����CRRI���6U��)�X���)LmLdFc�(�YM)���'�yCrY6���C�d�"gw��g��;�=�nl��g��5���>���8����:e��R�l��+;,]9��I�@�6t┥ ��3�y�w?�F�o�(�s^q|��w������$޷c���'!S�����C������;j˹s��������@uY}�[�������#֦v�{�����;��,M���	�zf#�s�n�J����è�Q�-�I�ξ�9�1o9�����?* ���ښn�PS!ώjf��D� ��]�{X��J@lF������)�t*Z��2��,˭�kN�u�5��܋��6	8���ʢg�r@�堶�?�v�j䬊Eۧ-T�a���ۚj������ڭ{M����xj�E��!Ϩ�3j>֮OW ���&��7&e����E�}�yY/�=�.��Lrgb�2 ��n��5���H}gW�/Lb��*�����@�]�,��,p'�߽�������y}P�mU�<�%۽5K��{7D*"~̵C���A��g'�7T�{z����5#h&˶.i�w����͉S+�vw��^ɳ/�1yN?\zQ n S�`��!�����?���C4k�fOg��/䚮�Ւw��Ǭys��T�dM�}ؑ�?+�/Y��������������ͽx��&^�l oY����h}Wڡ�/��Y�9�?������)�S��}RD^[s�j����\����_���`RGQ=s䵐��E>��=�j;㙔�mzVE�d▙�����@O�O��Q�<��?�664�z2'$��!���񤣁�^+Vy�'�=�&��>� 6$�rn���,����BUT�������������h�݈��%�ƆZ��2)<"c����gIqqG2�2q�����M�0���?�G�NZ�U�8��Kj�vI�y�Ï�#��P#K�e]���H2k�����P++�}��^]˘aØ=�Q�M�L�G�jS}qL�5Iŭ���F�ZZh�����A
|_W*#l韬cE�Gt�!�,��b��Tο^;�p��H�B�IU�5.�3��{'�,͓�aT��(� �L�A�tm�fU�M/�(K6:�}��dϬ?�,�de� ^����|*�U�㶎N�,����i9�����J8�D)�̭���嚯��9�lG�pd~��cJE�~��#O�r��B?�ǡ)��{8�����56��#�04��r���'�N�HVw`e'��x0�������t{����/ܚ?�M�s�ks3�3�es�v�Z�]=4��a�O�\{��\���G3��=-��*2ș1p�a�
��[Rϻ-�4�k�#�Ȑ@c3l%]KI���ow�?!Ou�W�� 䵃ރR�V�����c�`7G�{��0�c��~G/k^֝�eIx(H�w�Y�K5ն��1�&������A'_7$&3�k��R����e|4o<�^z�/^���U�yw�V=5����w_X�G�V�ɫ���Օ|��yM����V�奬{e�__����%�>~m���uo.b�[Kx��gxw�<�>��,{���>ŪEO��ʅ�]9�g���c�9e�f)�3{
�Ǎ`@��t��!.(�h� ��R�_B��R��V��KNV�dR�o�<;���1����HF7$3�w6��2�&�{%0�g<S��ՒDOC��7��-q�4WW�%;�������+?�؈v���'�/������j��vagZ?w���
6
�M�w:��ϤR�Ux<{s8�֑�eJ+eR	;��9�^�Ş�,�O`Q^_��e���[���O���v.d&�ѽ[#qqq2k�t-�ȓ�b�g����TL���)f�tIȢ������92���dj �RX!oW�`x�8����:� ���ò�{������[kVY�,z�Īy��պ�W�ڋ�0����h�lُM��X܏퐃8���=8K:j��A�Cm%z�@��Г8�8���X<���o5�-止>G4_uj����޵K�O��Y/�n*.�,��x܈i�횏<2M5ٚ7�͕Ϡ�A�ee�kډA�t�]�/5�k�la�E@�~���b��Bʫ��J��S�X�3&��=���ئN�6y)�c�9���t�y�쩘���%���Z���|��g��r[5��t����zc�����F�zw����5s�^7���fq��R���uuUV<z��m�v�SS��vj�v~h������~?�rR�' u�n[�_�<�R�����r�SΞ_��o�fͺ���N?_��[�52j��a��<%���71`�8���$�^�kX�cǎ0|��;��RBA�Rr{Pҿ���RJԑ�RCv�rZ���WC|�2��Lg�韴N~��������ӟ�'I�ä�n�6����)3��px�S���2�=Զ��<��M׮�K(�w��	.]����F��IT֒*�s�s��IA�uj�iyW�Y�QH�3�����bDD<��nR���n���!q�,z#4���x�+����ͬb�ĹLM+aj~%[^�ic�:);��ҽ���KЯ�3���Z���@W)�Ml0upA��#c=���137�ڲ��&x��0c��}�j���7ꀛ����*�΍�E�:~5R ��a�H���v)f��N�99akE���]*x⩙�y�e�}���c�����ű46���+kl��d/�hc%�L	r��0Ȟ*
D����}V	��y���V�0�������[���Ʊe@35؊L[Av��a�3@_ �X BY���:�'�a2�{m�O��ua��J�gd�S�C�Z�̲��
��p�-bIe/�G��k,�5��G�zS$kz��<\������[��Y��׺G�r����\�/�J�x�ċ'
ݙ����4�%:0"مIyA�L��K��nf�:r]MIw0#�ڀH}|�eN�,���a$צ'2�ӓk��"e�t0�{kc�=��/u�:���~t W���Қj�o��{�wJ	Ox�k�#�J����\��^��������v��h����Y�>��mM�>�>Z�}g3���*�"�\G����+yy|w�\��#�߁w��z3�2�E��Y;��?ҟ5�Z��ɉ�}��6gw��ܾ�8������|ťS��t�N���g���	~��gl���-|x�����;8{h;g���_qb��g޾-o�s�j�oYÞM��w�+|�����eM�6�Ƒ�������!�6�a��ر�U>�`ｹ��_~V�޻W#ə�G�����G�)t�(Ԛg�[���Lr�3�w
�Y��ԕw_�˻/�a����<���O���ԫr��lY�ޟ͋�������Bv5bMt*W��7r�[~9���/�d�#�Y;j"o˂z��Æ�O��\ܻ���N���������'ds��O��k�̜���CY7v"��eu� �?<�ϧ?�Ǐ>���+8��:VM��غ&6�����l�M쉲�$��gC;�,�q�ʟ&��Z$�*��Ѷ�z&�W4�ܒU��fSn�ļ�T��®'�2*>���ἒ\Ū���{��n�j�����ٍa��5+�U�=���.�t!ЅN@/b�)3�*��]�s8t���p.��gJ^C?!NU/�P�
��E��.��B�R�=�U�/���!���ƺz���a\�	���q�{
���Z�Y�1LZN`���R����Q����ѥ.�|�	����7�C���~�Y��;��'�u߇�I��lܦY#Z����%����Y�ϰ��|�E�"���cI?f�Ȋ9�Y3��^le�SMLљ����%6�7
�§�Qöُ`ӂmH%��d�ePX���I�l�\*�GJ8�K?\ƥ���ښh�7T
Zy�4�xW�'���ў�L���R�j!����W��<�M���鵳����;Ǐ?�� P�_(ݕ���j���2�wR�W)���	X޽�Z(/���^x}2������9{n�|?�)ϔ1|F��Ng��Y�XNi�b��+i=��G�r�΍��5ۻ�(�C�Z���n�U6�QX�Oq�R��u�������^xV���������+\�Rf����| �t�ԍW�����mM�
����7Z�������/\�t�o�{@�դ���+����ɯ�X�� "�ͱM�%�L ���6�Sr���օ���%��s����-��.�[;kE�x��{
����<�a�J����i6s���;�)%���|g��n��3=��-[Y�p!Eii4��`�T6�탫�U���� �V����+Q��R`���M��/��AĆ�2c��|������,	�2?��]��P���F3 $��8C���rQΐ��,�Q�M����T�����w���i>|�Ur�Sp�k�4������V OIA��y�y�V���3&Ï�v�3,�����L78���N.����5��?L��9�i9��������s�ʕ�`���)�=
N��M�1%�چ@,����jj���!��D���nJ�@_��	��fx���˒;}J��tP�0���	�>��D�)���@cz������jH�c�cGK�Ma6t���ה
o���(ҎeMU�+��.��Y!��dI���Ύ�{���F��=�r��u9�ah��N ]��Q�K;=C�M�	�kN�7���B��;#ה/&Es��CR�>8���G�f����h'R��HVbH/CC�$�v�s�����w������+, �؀H�"���k#)�u�
LV��P�C�����/����V����#yn�^�5���d��~�q�ߺ�ﶬ���/�6����Dw.H�}�k��k~��_=)��y�������B"޽̝��s�Ə�e��ܾ�����W����\�x��~����7r��GV�ޤ��w����v������wq��q�_��s��kٱe_���Lf���4���G�(<�Tl\���̢�c��I��%���NnZ6������C���U���a~��?����_����%?�(��\�r�/��J���X�־#X��G����/8{�&jl��K����Un�~�s�N�p7o����s���[�{�	O��u<s�r�9f4��;�r@~��;���w����_�>|���v����ɔ��0k�L=�_����|<���� =$���2�����Q��1e"�͚�ܹ3y���<6s�[{ӭ�P{�Ҋ˙;�y*�o�3!�:��O<�A�D�P^L�di�p��&�n9�2� f���׬h���
���ac=����Ď� j��'��v�v���Kt٫��<�.|,��1�b���Y�e.¸x��D�n՚=���{]�l;]��yܳt�{�m���[B��m������:�����FW�Q oFy�c\�6�M�0��n;q���٫�\bP�6f=�ҡ��{lk��s7i�,��	��_�$���ՒN�<\'Q��1��9�O��̙��qm[/���ʮJ����lZؙe7ѹ����:,q��cBo\c�ͪ#_�˺� ��g_fq�d1G�o�ۋ��F	%����!R���oM*�������g�ԍJeଇ�V�'�z�k7�p��u��m[���Q���w%�����u����KZ$�v�� ��? �o���L
�Ԙ}y*}� Z�ԏ���+�͘���|�4._�-�2��{���ᎢN�=:�3��fݣ<<g,�[�7a:GN�&�KX3���3���:<��q/��#�~n�e����xs.�ķS����� �"��6�/���݅!��������]wwwwww��]繫:d��}��9��[�;����W=e�p�X��Xz�*���/�S���|�E�<5�VA���[{��#P�R�Q���C���?�o_T��O�߰�D�y㒜_ชt�i���<����/O�<C��zc!`��섫��������֬�li����R�U�M�`g���)�%;l*��Ji���$����^��r
i}�R�J�G�B\�d�>D�'PW�חZ�adFDQ.8�bᑤ�E&���H�B�T/�!��Y��P`(��7an�ALlҒ��;3%�m�ܨbbM��9�PjZ�c+��,	���dZ2�'c� ��#{�q�'%��S�.�N��Xbaj�/�gkm����l�C�`��dXqfe�rnlY΍/ü�~��hǦ��y�XJ�����lK�?�ʑ����҂ݒ�\Ɵiqδ���,�� Oy�z:l�谓�8Y��Ⴟ�=>f��-��0��R Q5dv"���]K��T��:��k7��*ǵ�y|{��Z���mn"oIh��
�r�$J�<�ٚ���ĺ[��M`��BbK"�L~��@u6'��I��>1ȃpWkB�,��0U׭����F���+�ڂ'�TkIs��Z���=��QM�&%j�u����ؐ�s겫u�����e���	�����S~�	y����vJ���W�� )P����&p�9�V��퍤�#`�(����I���#�΂�NkX����|R���Ʃ��8�w6�w�Ʃ#�8z��-���|�z�����#^��½�G�s��_^��}���P'fC3ڂ5��(�y��(���N3��hj��G���|x�7�/���޿9Η�g���4߿���)w-W�㛊ɺ�<}r�+�ױg�t֭Èa-�VY�Ӽ��!��$S��8��#od�2*������R01ESFj:�'R<� ujU�W��ҏA�;Сc-kż�Y�d�ƌié�˘b9^�b�2: �A�:r��C^~����W}�X�d&9�/�|�\���HL.F��u��g�ubR@�C�ػ�(��I�'�P�*R���/?x���%�y�$��fR6�2=�{�d�2���3�!�œ�m�ٱu5W��܅�ܸ{�'�����5�>>ϥ�Gػu����Ց�"E>z%�V�4�alh"������t�������Q��R[\q�͏���*N�.cY����h�eP��5�bS}>���>˄^�?<�"sp�ڇS���җ��7�B�1/���Fa���e��?F�o���0��]�(I+��6]��'�+8]����~��XW߅�jf��ܴ־���,�H���<�S�e�fȱ
�Ŵ�r�����ܵ->��c1�?��k��{Lk�ͣFW;���!3ɵĲ�<�·�6\�O$or{F��������77W�ܒT�oJ���(�����h�/ț�1��β��tkGrZ)\�+�S�ز�*G�"I���I�>��ۙ���s�ZY�>o��o��k)�&�O7�o�� _�~�F�����t����vW~u���W�<{ɫ����3�'���,�WͶ?|��o���-T#�o�;��!O�3�U���O(7*o�%�9A��c(S�k7gKʑ�I�v~iU�iҵ��� ��M�0r~�kG���䛹#��w�S &@ٿ5X���!o�jxW��K��y��@Q5y~��.T��2����o�8g�$�qs�o܊��U/���%�3��2r����{f�0�o������y�_���7S~|�����(A`��S��-Q�_ O�.[��U��I� ��'�6NDz�/����o�5����al���P,`!���.��$e�g��%dU�K����bI��P�����@s�1���n�y��nm�u�WS�U�q��_�-��3���Z��R �� 'g\l�q�2$>8�0gwb�H���JZQ�U�bG�~l*��栂4�'I@E�E~{'��l5'����lX��������?z��7i5�m�7�	y�y9͵�����^�ͳ6� �J�+�Ն��A.��|q�_!nͫ�ɉe^ޑ��4�wjb��۳�yi���#������p�O��ew� �%��"r����k������<�m����`m�Ӭ�/0�G��O�}�JՎ�ty4�e}����`,�K-���:I��W����*VM�f�������!�f�ؙ*��J&�M�����U�T�c ��dY�X�ٙ�p�5����<xI/��!R��]$M��1���]�)�O�o�F��V0�G���p�3�O��۱6��P����q�S*SJ��!�#�C��k3m�� cCf���Ԉ��p�2%�oP��������-B�"���ɍHI��An���Tow���hoM�����](���ҵyu�vj̘!;��G�`��L�օe��r��j�_���['�v��.m�Թ-ܹ�w�QU}y��U,�2�_���S
�r�|�b^T���C���;��5߾	~���w�4}�|I�Z~��� ���ܹs��g7q��
���L�ڛ�=S;�i�	*T���J�/�$~!�L"6&��y�@B�D��
h�W2��6ZDX��l"C"(�X�"�S(T ��%+���ũ^���ׯ�(j4�r��l�L���@�{M�;r��mn޸Ϛ�ٰj3���w�q��}N_�M�A82�N���Ɠm�/@Z�%��{p��]>~��w��y�n�9���o�p��E���I�t�"�f6.�JBp�fv����{�w�:v�^��œ�;_�t�d~�6�1��ѿ_W��J��5�J���b��	������3##���~�ϡk���q�gfZ%���E�R�	�:�qir��W�	��Ī���ˤ�E�CؕY�.�'���r3�����q�{C��<��Xq>��Pg���;���]�dL*,æ�2�
�ô�,�lŢ�~���­�^쪯�t~)�1��Q�ä�y����v�����b��y�,ļ�t��.�ܘ�|ڣ�n�~� +,�<s7yj`<���	��<�Y�Ql�N� ��Rs�q#ɗЉq]quC�,����_���پ\Z΅!��Ʈ��^���Mf<������?���&0*��B����X��I1H2�Is;�e��T��O3y��~4�����|�V[[���2���-H�O�
�ظ���.���W���g-�
���9R���AOA�����M޾Q�4�,!�0�xJ�<�����A����A��Q��֋7]���Z퉭P�	����4n=H���$�O�Ϙ�<x0�����sxE�ʤVǦ�7�'ϕ��@ޓG�;r8	�kT���I]���#�DC|S�Lk�{�����gB|��Y�ճ�1{�Z��R�<��ʭj��Lں���:H�/Tsk��U��e��
�L�O�k������j���g�"�`0>	���
����j���S}�|J�'�R&�e��7��=N&����Oh4����+g�^b�jbGIIW����7u�Dr	1����h�'�`ШI�4�>G3|�TF��A��iҸ����lѪ��xb�3!���6j"o)�g9�3��#:o>��,HǮ]>f��-d��g�~t�0@��f�4�����0�$���o�@	#�ML	�w �؊h��]{���^����G�r��q�^����=������	ܘ�~��V��)�˕�	���L�t�m�?Ê{��U'Ԁ�Y��۽(�J�0��5'�
�������(Vn������$x<�����}<�K��5F��������91)
�$��30R}�4�ˣ��@��N�P��)������5�SR��)�1�	�<z�����ʅC%5�9WF
����MD*�sJ@�ӓ��ղ�ί�������:S��kdC!;�;�S�ޒ^ִ	0�gDF�ú,>�/;�éw���p3��l��s�p�s�2��L�(GJxx�Yi���;S��������Օ��`�?�j�U�*rk�TS�Y�zʅ����'go�]<H���Q��kP��U�h��B㲉�-����i\�0Y��]$��E�Y���T�i��4�P��e� �4��mҷ]z�k̐�3�����]8s�M��\<v�G7����=�߿��Gwx���}���ϟ
�����ϼ|��׮r���]��勧9�'۶,f��9�Z9�9�G1i� F��Ψ=6�7�{w�_��߉�b�۵nH�Fu�W�e��`�X
� �P��26.�|qy���9E.�T���BP5y��R�p��]}?�^�l�}�1>����F>� �B"e}�XX�-���gmp*=-��@�GhD��b�L�5�I�qf�An���٣'4W2��̢pl:m�W�����h܂%�����JBI��ʩ}�ٲt#��b�9\<,���]�_O���$�&�pZ��$�~+��$8�(ߐj�(�Q���KR>���%$=1���x
D�#�/�����8�`�gI��Y�3(+�n���n?�cg�5�<���Q�YY}�Y���W`��0�h�S��95@"OSQ���5��Y�m��b���:���1�>�a�x6����<t�ô�:D�* ��<��j����8�̍8�X�.n�v���Y[uΐ����D�f������Qs�5�J�z�^j�3�r�I�Θ��Gy�Ĕ��"�a�<ӄ�����fؔ��m�}�>�.����6��Y�:aS�&���[v���\YY�ӫ�ui$���ڲp�N���� ���ހ0n���Tw.����eE��*�*��)�7�D���7_��ɤp�f�-㦅��h'/��惪����g���{�6��������l�/Jj�H�R2q�|^�qJ�Z��s~��A���ͷ�@�Z�@J�?���倞
�6�ٳ�?}�>�<^�I��uuMS��=�s¿Tj�ETǉ?8�����ƷLs�զl�����G�$�z2�J�2{e�~���]���-Ϯb	R�d2n��y[9���y��'��|u�JVūp<�J�[�0��i�ο+Q�n9j5)I���:��w����m|��N#_��A����۠ O5��8�������L�O�k��}�&�_�]��ҍM�hT	1R���q+� ��� O��ET�IX�؇�b��A��-��@/���s0�$�.%zC;W�����އa��Lpa�s�l�(�Hʹ�tlڞ�r�t�ԲNKM�뷡EVzd�``�~TI,#F�9n�d�-u6,)L+s��ߪ�1�ۏzkб^K:�mF���Ӷ+][t�U�6�kڕ�-�ӦQ;���MG� Ny'�4� {����̉��US^��H^Wꖫƴ��g m�5fD뮌�Ѓ�R5_x
f�4�|6VfXYcee�#Y����j�"����׃�)�L�������8�,V�ќ$�I7czG΍*ɫU���1_4�ݩVR� c|��{sg\e��H`f� �;��ל�vz�Ye�C=\��d�vX�j5mʕ�0V9ʁ@����jĪ�����3)�S��+}15�7W���"uU�j����0�7���}c�*�dZO{g�j�`S#��L	11���E���FMG�{[�.̎~	�/�ˊ�a�l���|]T�����k˗�-���O�Vdw�H~�0aj	ƕ�V�INj{Gs���B�\��U�k(�̅<5%�6��O�S�/�	y^>�x����)�Bd���f+2sX�M�ʺY�Y9�?˦a��ᬞ5���n�TV͞��3X;u6�'Le��q,�0���'�r�x��ܱCӷ�������Lٗ���1s�`�O͒�Y�`��;o��y�[2���q�B6�Xʦ�+عi;�lf��5,_�����fLe�ԉL�<���3F�;lHw��"0מ�:jq�nmڿ���z3zX��D����ѥ#];��u����%.6�Ԕ$��ŇkR���5ۅ6�YZ�V��JH'`(�"b�T���cb)�D�r��]��*�f_�v�*AG������5K�g߲u�9v�W������}�;O���݋�\>w���ʐ]�$7�N�Q�n�����3-*�eͼ5ܻ��{p��en��ͫ�ox�����z�LX|.vAbCڱ~�zR��g�D��I�A䏈 IT(oeR�)!0[<>���x��q���\�FdG�2�?h%�
&��f!q��5��c���P�z^��)߀��Bɾ�T_�E�?g���y˻6��i�[��*�
]����N����M����<&����2]Xo+�������C'�^�qt����ƥ�*�*/G��
]�`����8� �M/`�� �	���Ǵ�q�O�8�:j��/M����9�.�
��u�*�/!5�c�6]h�K�Ư��iP�\c[ܪ.�&K O�N��I��� ���~y�v�?�ҙ�80�����(.lI�ئtnm(���^ܬg��2�<.�ĕTN�udai��PM�&�:���Q�����8��W�C��ũ\2�ڙN���=霽\�[*��M5^�Ƈo�5����>_h��?����5+���E��,\;�ן��d��������A��b�
������X���f.7��w�<���Z��_'w�R�'詿����G��y�?j-
{n��b��xV�ƻB�K'�|)"*T!�T)b˥���~���{o��jvc�g�g��r�/����!O��8e�b�W&�LY"Jg��r2E�FR�U8�`��j�:Ӏ����}g�~�/O*�>����9m�r��߿kC�s Oo.����PՋ���k�}��O����ܠ~J�?���~�����~��XB�.��,��WZ9<ҫj����@^N���
5.QS������om�TOV{�Dߊ2�qv�Y��#�c��w㨓G]8��u^��cIy���:+�9S�ԕ���T�5q����Z.a�F�gYցr\s�籥���h��'���+�%�T�lbNqSg�Y�P�܏����ѳ���-q����7���Z:maK1#S�����?�k~���G+7���0
vv��z��N�"�	�r%���&[#c��[c}�<#�<,-�4�Ȗ�y~:I���'����B�|���oÌ,��JӦݺ8�[���Ĭ:�Y��+j�zCM��C�O@�\Wx��τ����������,��ΘzDX��˒*.֚�4g[m�F�����y�0�1΃���֏��X]�fFv"s�<�r�>J�mɯҶ�kM�J
��ZY���7���R�C�����������6"��1��M)aoBo32Lil�9��fB�(3F�Y2��%�+ٳ��/Ǉ���ڼZҐ7���}MC�ސ��2�~�6������\[�UM��n��z̫�ɠb��6$��X��	2���*_��&ￂ<�O�ޯ����OA����yn�������ꭹ�)�??��ve�ql�?�c�Wq��FN�$ڠ����\����W����In_:����cܾ|���s��n��':čsG�vF��=����WN�ܱ���ř��9uHi''������8���Gv�5��؁�8�S���ʁ]9�g�w�b��e�ܺD��Y�i����ڼ�}��r`�I/�ۗ˺el['�f)]:�%R��̒�	��ͧ9@�Ml|$��oٞT �6ZjZam96>��@J��b�dU,C�aW�<�kW�K���؇�;�ri��gvaW�6K�L��3Qᴂ,���O/>hfZ�q����������?�����4�Bi�����ww�:0Z�OŰPf͞ƻoQ>BU�"e��'��Ws�֞��4<,<�ْ-�VQ8$�.�t�V�V0lh�V,Iɢ�)[��RR)������FthI������Z����;���	Zmr��S�g޸�$&��ΓΕ�+{i���Wu-��Nc���6��y��X7�����"Oq���b^ev��a��"y�_D��El����jt-��6Ŭ�|L�\A���5X�e[K<+-¥�B���]p+;�
���*˴Q�Fe�cPy�Y'1�5�����c�����>]0��Mp��+��0y�P�7t��:♹+K�Z'ѯy���{�0�����%O""�3�'������d��Y|�ׁ����ejQ��N|�1��MO�ƽr�h��u���ϲa���o}b�P$w{k��iS���GP��}���lm'N���r�V��o*j���~�����|�.��SC~|k-yi��hÝGy�q߾�޿ˏ�]ȅ.�
�rA�?B�z�kǅ�׸s��b�.V���n�sj?(gj9כԗ�f�UM�������o�3���:����N]�����TN�w��ZW9�B�f֠ߤ��Z7��;f�nX�un���[�� ]+A�hY�~%U�W%�Ke�N�����r�����6r3�OY����߿4��n�{;As�ݴK�h�Ǯ�)����������t���s����ϯ��琣_��l��9���Y��*Ot�rڠ�Բ�tf
�
�� O�ы*_� �C1Pfff�tt`�_+���&Ʒ���ΐ�&nl��_J��$ާ3�eK:���ɗyblg*�A�����(����4#0���y+�cd��~�a�_,]�����
�HV��D&3;�(3��dU�JL�M`�s,��dAh<�Bhe�LEc;"tz�q$�ֆHsS��3�ݗ~I\�Nf�K��\��{p�ףj��L�0��u��Pѳ"(�nF�Zs���g"0cai������>��N�:LU�<++L&�;�(W2��hmˀb,n�ѱx��Og5dy�h�Ы��x�P��|�ؘ�ۚ��`;���7
�M����Ps�,��Ց���"��E���F�HG�9R/ā>�s1��}���P�5g�mwK�Lu�j���D7�o����|Dj4�R��Q���R���m��
�47(	��$�R�N@�ΈR�FTp4���15|��dL�:�;0��;;2��#��qezYW�d{�0.�+̃�J�cW3�Ȇ���� �݂/���1�[��fg&��T�����δ�nt��{���-�1?+����D�=�XZ�쫹��0�Y�7�&O�%T͵�jԬ�^XX��'O�]�O<��C�7^�8{y��!��V$��2�S[VM���3�#@�@��>�R��v��6�]�ˍ+�s�(O����%Mj�٣�~q�7/����=>�z���?�χ���	��=�|�*����^��㛇�{��7�?���{<|��On���M^�~�g����ݽ��[�w�$wo
\^?���ݓܹv���q[ ��}\�x����s��6ΝP<�Y�p۷��n�Z�%1&��M|R^-�M L)������E��S�v5��fҭS���o�1w�hL��ֵ���.i���{�0�Jk����d�;�$=����a�:���š}'��$�������<x��[�r��&�Έr�9�~4��eV|1:U����G���sm�޹3g�z�2����ܹs�=�[w�j�::6�LzH2]k�a���D���ehJ�5��g��մkےRŊ����(3�a�пK?zv�ż��٥��	䍦xd�6�����f��988��`lC��M��ai�FPk΍.c��
F�.	�]Ʋ�L�m0�I�4�+.����5�~�S�Ի�u�3�0����U ʯ��f`^�<���0�y��[4���S��Sq�������E�I��F���|=�E�i�����M'���'h����]���Y�;������f�ĳ�b�d�D�8�ҋp(3I ���nxg��6��:M��3�����-�|���:Ӥi7_���p�xQ^?�Ȼ�8;0�c)�v�}s;��Z�E�˻�&\Jt�H�|\�^�;
�kE��	��QG��]��UV<�+Xк��燱}O
'Φs�^�M���wUy����|��c}�|ņ�u%#n�q�w~�ӗ������
f��A�U|����w�r�T�w��������mo\�'��+r9�\r�C^�+��bw^i}�Tzuܜ����f�UZR����<}�g��/�/ek�o�NUp(Tǌ򸗬�g�*�%!�lJf7�^�4�߂.#����.�_߿����+.�e��F��Q��+s�EC^}iƇ-x���E|�ڄ�ߚ��c��l޼j˳���&O�žӀG�Xy 9��3
�?��
)9PѳjkWᯇ����� ��� ����ۗ�Rß?Ǟ�q��*e1Lȋ�@���&��\��%�a[0��E�͟. X���k�����>vZ�9
�켩 �f����.,2�ә�V o�h��Td�vY{����#n�v	`�d���}���n� v{��E�y���ڋ�f��-Φ��,�+�h�6��gwcu�6,(V���
�;:�5��,K,��"���^���8�k�����֞��^���b�M0�<���:���!_��΋0r�45l�����j ���%f����/�E=�<��DK:z�:�?���1y�064�j��ݨ��C�$�W�f��|\��"@W�[Ӫ�*;��%��]%��}�r{f5~_^���~]=�f���6�q����H.�.��c=x��%���fc�4f�h.��T7F�eh�-�"��eM�ps��R�FG%+Jˊʘ�(%qi���m�uT�7$�Ʉڎ&�w����--��i�kF;o���5Ȝ��6t��g�=��3&��ȓߊ�1���y��]{�%qxh:g'V�ƬڢL.L��ͅ���_��&* ;n�3]`3�E���x��*/�T������ʼ�D��8��[�����>��ٱ��q�4��O��;��C�w�vN8	�+�S�ۙ�h��D�H`�/~��Ss���0������oO��q�����3#��<�Ң.ۖLfߚ�ݱ���p��&.��̍k��y퀔�Os��y�~tM��W�n���]����)}z+0��w��.@���_i���5�>���_^I�Rӗ�9�,�(}z��������_t��/ _\��3���Wx���@�e�9�]���~�8W�;{����r��6�����(Y����D�@���1��I��$&'
�%�\P�J��d���Q�Ju&�Ǡ��<�?�Fgޤ)��m:���f���ݻ���0g�DF7���F��R��e�X1q3�Lbt��h۟]�0��P�t��>��<b�Vc�j�Z����N�9�c<�+�dV�L�����ә�y�gr���8��}ưz�B����6���k;��cdv?z7�΢9��n֞b�Q�b-*H��~��Z���R�l5�j���Y>m˦�a���޼�y��a�v���N�_$>v�:�w�X�O���6M�-�^�6]���h�	�gn�f�PN�-�������NWr1��~�UX�O��5ݏm����=�ai���)�U]/�7�GS���ؕ��}�3�e����a�J	lٕE�]��q��Eη	��K�L�������EBW����5A��Jk�eC����ʁ���RFu.bQ�(yR�h�u���T_�Q9�˒0+'י�:��r}5��0�:��e�EW����qt�wb��W t?>�ѯ[[���ͥM��<%����1��3L�f6x�=�!���N����<y�Č���\�Í=���l����"L)�I��
4���Ŭ�Vτ���X�.�#�ӹt�W����R<{'��/ux�����0��Ň��x��9���ķ�;$�}�������W��Or������\�xM�JU��U �[����k�>~ý;�xp����k���\�0�����ʩ���Qk����w��S徸�i�g���d�U��pY\�
���G�r�T�Nt��$֮AR�
t4�ׯ�|���V����l�ٌ}�Kɭ ����u)��*��w�x�NJ����c�@^{�����n�|9�w��=���,�I���~Y��N�_��ۂ���Խ¢��I��=Q�
U�3��F�EKc_�(VI��x��%�)]�ؒհ����^���ɇ)���;SZ>��b�����Xߖ�yLY�Ǆ5y�ؠg�V��R�ڙǚ��V�hک�g���F�w�h�h���B�my��ةg�΀��|��N`e�,����&�%C��іݘ�4s;��-��v��Z�>�-��%�9f*���2�ڕjFf����֎{o��=Ȳ�`�{8G�8-���Ε&��n���8�6��$iʙ9R^`!B�Z�-AI�:�@Au�7âfgP���Ƚ��g�"�w��5��L��SA�6����$�ϗ��r\_�U�#��΄�l����ex���W����:|�وO���H6�϶���po� �Hx����x�4
N����<�Z�K�p�[;���f~�U3���ܙZ�E��\ćIތ-����n��(�ʐTgF�y2�D �K1�X �J�0�t8��G��l+��z$��b��0?[�f_���]�{�Z�`RK��k«U������*����q�f��R2<M��k�:X�_��#d�?Ov6�����ؘ��+*�1�pNIN�(����nL�'ZY�&Ċ�բ�8�&G{�O+ʻ����L�� �ʛXw�0�m��������S͵
�""����@F�W�����Eb{'�~3<��h^�2N���ٺ�{6q�����έ+{�s�0�^��}���w���/T�c>�~ʧ7�4��$����8ro���[��?%E�I5w(}��>G_?j�����_���=�Ǐ���A���>o���ݛ{�yyW��&�?���GW�}�,7��^?����8p|'O�f�ڥZ�:5��r�M\l��F�A���">1I���S�HN*L�ڍ$��ƺ�f�l�f��ܮY�mۇMcˤy�7��=F���D�����Kwru�6��Yϭ�{84i)��.f� ��8<u%G����o�91i��ss7qy�V��_ǫ��9n;�b[����?���G���d����^���{�F/����l�6��}gsu��M^;��9��$;��ȡs��|����x�F������Gؽ�[��d���ٲ��vsr�*.�����[��r+:���7	b���1{�\�N�����N�kК=&�V}��6���Eͱ�r<l���M.�_i���Ѹ
ȹW� �]���	�%O�F��Y�m͍�ҧa�6���/�Rk\j����.�#�egc]{&U�cZf1N%��Tx�������(I�PY`��@�r���r�D��L�.bW�����l�b��=Nu�`\���G���)�9�Wt�uq�8E���#�������{�(���������ȦNt���]9��1��GK8p7��r <�u|��;��ۊc��ٻ W��sjS!�t��h~'ңB�*]���Ѥ��\�-=F��fK!��+ɥ��t�W�����<{SC��&o?ekR�o_}n������ď���{�������:|RΑ�=����\�z#��N�Ī	�û<~��[7h�y�g��+x�	��?OD�;�G�zx��W��"�WA�8r)R�����El����"���ƌ���GZ�	zo�����.'���᚜�X���x�,�_��:L��&����}6�?w���|��O�D^��ė/7�ܼ\�"���V��/�W�ϟ?�ӯ]n�u��5��
��hM�ʅ�H󛥦"��/$���7���&�9�,n�b_H^qR
a���9DVͶ�%�hs��%S�����^aL򉢹�������,�pX3g�Δ�y����`�@��M���o�Β-��:I�\g�R��,�7g����B�ϊy��̯ ��f��\�`�9��<&��-�2�bc
��Q;�L^�,��9�N��|���������8��!�ڎh+;�QN_�I������|�t���s��@�Uj�$�L���c��'���DE�"�ī�����䙨�"jz+o����r�M���2���E��!�3J�reE^��̵�J��A�RW*���O*w�T��e:˫�iu}�miG;��DG�8�.�ɩ�z$��|���@M�����R/8ם�����μ:ؙ߷���L���5�O�V���ܜV��S�pyR)N�N��rܙ]Uӭi��?�O�e�ha#�m���;����h^͋#�xwf4_����[���2�UR�{& �\������̕�[��Ӌ��:��V|ޑͻ-�y��ϖ��֌����qlk�Ȓ��)A�p;*:��ѱ�e�Ge��G��x�fC��� y�!VDZ{��K��^��X멩��`�����n..D�G)pAH� ^h���!24��@?���/ޞ�xy{��텫���.X��hS�U/[�3�p`�bn^%����'�s�����Z��㇗�n���^��z-���V���:���n��j��f���w�F�;�i����,s]�hz#��J��O���=|"�GR ~���y��>O���޽��{p����s��Q��ˡ���0u�6���ӗ� �g1������G��/���뚔T�������զ'l�^���[��A������Y]�[���`��n:��Y��U�#g��r��4n�˭�s��&O�w�����q3{ �Z�V�!<�>�=�C?���]ƷA���y��,���S<�v�#C�s��>X��ο��d��������ܼ':�A�q��5�/�����v��C�݉n}3n�,�w̠��m$}���o�ں��zХy7�g�du���ۙ��p�p=��V�@BYV�G1�:�ή	�����M���L���趣(_enu�b��
捯i·��9��+��ۉI�%X��8����b�;���a�4�+o����6�"Pu,g~ׂ3���t��	]@{L3fcZl��ߌU�9�9à���q���w&:KU�����1�}��w�S�����@�u�]���@L�e�-��5<���nt�J�;���}�%e����N�N
L����A\J,�@��t�Ƙ��Lj�Ɏ��<ߟ�ە��ѯ0w�����,��g}����!ˈ~�n��Ƒ�Ǣ�>L�H����I��d�gT�T�D
&zR����I�vA�����*zո�6~���g��}Z���y��-/�u��Χo���m	|�*��Nc�_����A��S�w���ѫ4���翿�F᪚=�<9���y_?�C���w�5�/ǫR\J�ƫDm����]��ū�Z��zv�%d�,5ꐷV}�*W'�b�/Z���osf������������ٳ�	��q�B��~��M���������ؔ�[��Kg>���o�d��|��V��I�A��l�D��������Q#f�����O�W�y9ʅ<e��҅�.-��;�~�q��b�P�B�p(P���,.*�u��ȌKj�6ř���&At���#u,��x�hj��TK4�ʖ�fm&�����B�}+���Hߖ��v�׳a� �
پ�І����0w`��5����q`��'K�UceVC&{1�ʍŎL�bUݖ̪ј����I�ʢv�Q�2�\�X-������^��	�k�L%3�k-llF���ĚR�Ҋi���	H�F`2+⋳�q7֗����"܏��ED�&0�҇�fntxhm�A�����k��J�m]�i�@Kg�-��k`H��%u��ҭDm��3������2|�T�w��q{RE��J�j�F��3���{&sbh!.�����ǥ������5�˞�|=؁�'���t>��ŇK��~o_����/�5X�\#��z?Y P`��p�,Y�`���}T�:���^��e�s��g��l{*�/��$?�������V�q��E,��b�>���r&������|�)�tm������|�ߝ/;[i#�?n���Bݩe�:�Gb_�d6��Ҧ��Rɟ!��������-�_��
stH:�:3�X�L���ȫ'�' l`N��=��n9��nn�����Wi�g���n�n���k
�|ߩX��	��7���@���+n�z����3V6�ff�(T��ㆲm�llZ�����vr��An]>,�w���.���m��LA��7�����5w��Nӷ �V��S
�T&���.�Z�R���h�wr�~�d9>�T����/� ��^5����=zO�����k�:w�������tjI`p.�>�)(���i�V#�C�5%$Ē��Lބ��Q�p]K0!0�.Y�V��^�,tKb�g��
��+���ql�NaSp+�ҙ����+���v��pH��38��$�CӸ_��qe�僑��S�E5�<n:g���#�6�ue[�1�g�W�Lt	ٿ8G�S9Y����o���r1�*Gc+2�?��.�Tu$�ڕ���w���E�|(d�M~[�]�Y�3�5�-yMݩ�̨��.�I�lйp�ԏk�Q�tOfqXI����~i�A����oڃ����0s��b���ٷ�hrK�<��ױh~����/<���X�96*0���por����7Ʈb��@��F/~�	��/8J�O��9��ls�{
s�O��VcFc3�<�}Щ�y��b�4]�`2f�\�Ʋ�I���׽.R�R�U�&Ϧ��M["��e��+��+ ��8z�O�+�Z O9`�A�Y��k�j�Ԥ�~�p.>���pkO/>���b����B}~���p=łw�y�؈bۿ	�a���<�
�aV1��t�y)��t��a��9%��V�*T/^���")Tԛ�՝�;ȗe+�9z�<Wn��hȣ
�jh���]��iϳW=E}��u���4��rH��C����+�O�1*�~��N�Ѧ<ӂ�Z�	�]5�*�ɪ�_���=������O����] ��(��w��t#��x�~xE*�Z�2���qY,��h��YW�<�2(�ݚm�����O�S+���wn�d��l�"�@$���ɛL��͋�uy��1ﾶ��.��ҝw�z���P>|�+��EJ���h_�����E���/#w�\�Ԩ����c���^Cn�����j ���/_˲�篿Ҽ�h��`_�t\R��\����@^r�b�pL,�o�R8���]:W7����ǒ�8���S�.:��e��FS[���*��z���Xk�b(2��Mz��ֆ:+��f�����9��ȑ�ZM�5k��R�U��0^2��y��-�㥄�\J��J�f�{+}�XZ�13JVf�G� ��y��<�e��>o���	 PSgI������Y�lhLI#K�y3/�0Ë	TJ	~n��L
�`�W�bY�d�XFyF1�+��^at���d�=�X���͜����M	;w��0P����=���K� z%:1��;Ǉ�����|ޘɇUj0F��NbZ'X2:Å�Ճ��&�34Wƥ�pF)^.����Y���1�v4���F�q�	?��c]��TO~\���k��q�/?��珻C�
����x�^���~�@����H�<������cY��J#��~�,ϕ��fPN��=��`?����>�qC`�|>��ȧ��Z�/[�mo;8�^@�msޯ���Ee�=��V{��["�E3�n(�*һ�� �C��kBV�!mMX�:�M���>?�U�g{�FYR�ފ ���F�K�>�ȄPK�<�B��;^V�ZM��*MM �G�I�0�
Z$�
���_X��扫�����R���憽�3���XY���˸��ظx;�����>��˧�rM���r�{wN���y>�̓'�x��Vs�j�h)�Rͫ߿��Y���O�9�fN����M�U?m�(Ǡ�U��I��PY��f����5�>���G5#��y�$x̓Ƿ�{�*������;� o�g��_� ^���~�Z���DH>���7�0�^#�J$�sH&�Ű�1��F��4�c�U�-��h��z���:�F���M�Y_�;s�6��V~�7�d�����9�s�3�;>����׼2�f��@bF�|W3���g�n9��U'�@���1e8��e�@��qﺅs�5� #@ܿk.����u�a\���W]���ƍҙ*P���)�.�Z���/\���T64%���8+�-���`)Skz��&0��Na�s�Ξ]F>�H�f��8��х��ƚ&}X�=�&���x/6�n���.���c�}��w�hu�&'ѯu(g~�z��l$ˍk�ܚ�&޺�1nx��1kv�z�hp����jtAk�ի%i�_���>�� ��9��}�����~���8�;��3�v�z��տ���e�%�a���Q�+�1M�_Ƽ������Q�3�j����ս�Q�����K[)Z�q����.2�j(���4�~��w�Uj:��J���;w�.���ə�|9�	��r��}�x��i%/��$�aj�{gWv8��)ڀ�yud��(��OF�^��	�q�*4�^��eb)��I�Zt��΢eQ>Y��7Jq�IyQY�����}^��"yi?~5��z����I���)�x_�-������VY%RͶ��>�������	C�{��Z�a#���_vC1��
�_ȟR�Td*�����:x	����_1[ /���.��L뜮f!+�m��8��!�z]b�R�ae�Ь� n��]�:�:��!O������8:��;���`>�_/����j��[]��h����|�ގ�߻j���}o޾��7Ũ����*�WP�C�rK?o��6���� s�?���U�9פ�0��~��M�s��=BK��PJ��	��&�j�u����\Ǥb8��K��Gr:~��@
� �8�ik�H�>!45p`2f��=�-�X+n��P$�'%�_�fղ���6l�c�=���i��T�/�t���Yb`�5�.�S�q�$X�Q��m���]�w�Ρ!�XѲ��Ue�[4[m�Xg��*YV�k}c�b��vS�;+/��:��đ��^���x� �n���8;dfI��ie)��*W�æ2�\3��q���k F���=��!PZE����cI٧����Ry�L(kdFis+R��1��O�H�ѦܚT��eh�$��ү���rql���y��-���.g�f���?C�$��g��[�T�bs�p������$�L.��9e���nE~l���Z���#��� �R'���.��˽�z)���ѭ��q��V��@��-1X7��U�}�;��7�h���� ��=��
�	��&����J?�"ǻ��w�f�PӋ}=���}M���Y���MMy��o���բ��>�w'�������i���5��W̍�)δ���^�9uC�i�@�TO�����n���/�����jO�|�!�$�
ԉ�ךh�MϓG ψP+�x�ܵT��̵�xj�5�����^���z��A��'�v��Ο o|���������*r���E��A�����s��ޚ�0�vn͚S��
�-́���=�	n_;��gx&6���{���T��LU����|�*V�W��)�.W�5{9��_%A��\�uZ3�j�U���_j���zo�����ޫ��	y/�����;�8�xGO�צ��ר6�a���&62�����!!6�䄼�O�&�@�
ʺ�Db�K�O�]t
���Y㓏���3�ḥL�إg��G�[�gh��!�t�\;qN
{��N���qJl�	�-ܸj��5OMguN��s�qRYX������M���C�m������_�9�n��S�sG��3w�\����]c��{��ؙF.���]�H�	<>s��[�b�n�C���=�,v��*(��88���^�.P�Ԕ��AJ䲜�{��YZ����sv�$��K�_L64���z�iVaa��`��vz�-�hΐ���b��
z�a�X ��u�'�a�%t����ð�5��ϸ�L�]��������W0�V���a�'�����W�<zu/jR>���y�j]¤���Y]���1�5�}('�״t&��)3ٖ+��Y�"Z׽�U���׾�^�+�70ʼ���k\�(�UI��95y���*�W���z�v�>�F]�q�t)@f��J5�Z|�E]�q�Wz�r��=���x�乿��!O#f�л��*[R���z�i�L�(
�zS�Xa��.C�r���R����1gA��fp�v��{^�'���k#^~l��/=�'��s�~�ʇ/}������}=��U��!�rA����\�r][�נlF����˖�\��˹ney�>�L߹������m�.]���*QY�<m �@�SZ9��JU!�~s��mLh��U�Ť�kx�>�zr��_ O�E�E5s\�����*��P<'.�����wUx����[=^~����b�:��Gg^�k��w=y�b,����݇�y���s&�͡�������ϗ�{�\�O�h�jr �'��><��Ë_�9n��i��)� ]bn)i�)gȎI%4�)3���R�ؼ�{����@���b�(Ƭ�Ί�:w�م��Tb}SVI�v�~� �}��Էc��=b��:m���ۥ��61؛�lY'�Y)дT�B�Ϸ�ؖUPk��y3�`%V�lˊ�5Y�^�-]F�(�s\#�f��1A/V�h��
�Y�zk;��;��ڕM��l�c�vcW�۟#���0����[�('�mm�3�Xjqƍ�Lۚ���5)w"��DYXajA��9a�&i~��M4�h�G��cC�M̰70�Nҩ�nyt�8��5ş�%B]L�lh��1�y��,��;�T����*�i��iE�kN?���EݘXΞ�R���:T�������.�퉅y0)���*�vQUm�«�����_vՖ�W]Q8�T�e���l8&F�t;8#:ن'�o�|�-?�d�㐤=�������7����|�SW�[��;� o���~��N�
)�.��Ӆ��;�<w�W��o�8?R�<)�ѾE��%�M-Y�Ŕ�~�,|��J�(;����4��v�F�+eʹ�A,���N��m��Rt-�JV�e|\H�3�|����$qL���g �gA^Ow���p11�JҨAj��(?�����P�o��q���	���P	b�U��� M�a~D�h͒!!��y�/&�f��1eL_V/���ʩ�ݼ����r��A.�9��k��}�w�����<�{���_��ͻ����?���R��W��o��6=�*K+���c�sL�2�
�r�Q��?�xr��ߞ����޾��W�y����T{��En�8��9||;�lb΢�ԭ_���xJ��x�Z\�H��P6� �K�R�daʔ.B��ŨS��ڶdl�NLk�͔
��
' �0��p�؍cFN\���@�	���u�]�$@vM �Ε;\�s榡��<�����<�\�9
���@��^2�	,�ޖg���l���r��|l7�K!����YqE����7le�N���#K��x*����C Ӟ�־�>�����5�Ӯ�@�{���`�]0��^eX9P�ޕH������5�a�g�R���q��-̙��92v�yS�P�5�0���T���]���U˫m7�~p&��c��V˥$+w&�u����E���´�-�]�f�0�S�h(it�c��26�b�}N��kxA��Z�[;5����L�����K��E�����j�ƪX����:MM.a#�7��r����>8���V�6�}���0�:�i���G��̌2O��|��'�,���҃Y�L
�z��R^,ϫ�ո������*���_���,x�m̻�!l�����6l����)L�eM�f�4��E�/2�C��^��5�Q�jQ���O�2A4l����>lܚ��+e����W��wux��	�>���&_R7�~�̻ϝ��_���ɷv�_@I��J���W�Sz��.\��h\�}PRԣ�s� ^��=����晻.R��d�����\#�K���NA���S#k�Ts��^�>I�[i/��W�f��Ze����՜g����囚�Q��#7�oe��Flݛ��Se�t�
��W��皼�ZK��o�՗c���-x�����x=�;�o����b��k��j��GN��vc�x���?���\�˕Z�?r_�I�����9��sW�+\
����..���y�<�uJ�t\�˺�TCC0�t!�ÍF�<AJ�t��4b�C��<�TO��Ē�U��8d��A';j�g��^g�J	y��#;�����ٳAүѷ���),�E�س�*�y�k�>�+s<�$�$S��eq�&��Kf�][-�Y����=�Y�9|�Yif�z�ŝ.�����Mzr:O;�2�ԍR
L�	��&��V��<\!K�Z�p�r���/3<�-q�s0t�S���(l�����J��zؙ�633�%���!�����g����KfF�$F�adq'ַ����~_V���k�YYx�$���Y^#��qtӧ[���qy�j,�g��
�,�����ln��n���������˿ed�sob&��xF	��.����2���<ϗT�ɢ�.�ē�?���fi�ϩ��ie�9&��Ӌpcb
W�&q}|*��'qz@'{�p�_�{'r�G��ư�^ K�YV'�y�����;�x22Ù>q�t֣]�>�M�e�iD�?Ӫ���U,�z'��S$[�2���y�cKf�#iN�D�Y�'�$`��HG���VO Ok�U5y�n����j��hb���Vs"�)�L�5ܡ5���Ô�Ӫ%���HN�hJ"%
'�T��
ƅ�"I���`B4�y�H��Z�3�վ!c�cʈ̛4�e�&�-dۚE�ٺ���qx������{9sr?g����c��y��*�^����Z�����_t�7�����޽z�ۗk�7/�jz���������R�Wzt�*�]�@�Ν��];ť�G9{� Ǐ��'�پ��k��z�B�͝Ψ�Chռu�T�Q��4�Q��kҺ~mQ&-�֠E�4�^�&�+R�fU�լN��mY�h����܁�0���K2.0����[$'8a��E� .9s�9��Na\��薝�!�K�~�p���:���%�{��V�\-����,-X����:s=��,aCRe�'�bwh"���x❗���r�㖋j��c����7�v<���g,wC���m�(���X�=	H��W�l}y"�Mhq~���u�H30'ElF�����l��3&�܅!r/K=�1�#�.��9�m��P&4��)e��ݟa5�P��<nǰ�e�[45��E�C�[>â�]�d5�髧�5�s��71m)i�a��>��
̮c��:f��b�Jֵ�)�w�Ƨ1kq�l���0nz���ѫ# ��j�ͮc��
y�ܺF��or[��S��I Ӽ�@[�+X6��T-�i�3�w\�ET}��Tk�M�`�X�OΩ�I��ӯu�<��(�jBWm?�Տ`\��up+ù�Dz���-�:� �����K�92��-�֔����g�w#}���Vh[�{+˲Y"{�Q [��3��7�9R1#��"�)��ڥ�Ҵnu*W.NF�P*Uv�G?˾�O���͊�V�ǯ�p�i#�6���^��%o>7���VR`j��ʭ�@�m/I����j]�T������័�^��y�n��|�i0�vJ?���Q�W���JPN�o����V��|ѵ�Y���W��tv�[�)P�Բ���ţh��mN\�f���HT٪�2�Wj�59�����}��E�1զ���e��ž�5ٻ������~ވ/js���Z��ϵ���:_�W��Jr�My�j׍�ל�y��Wro���_�H= y
r%97��kN��������)�S��O���j����S���8U��_/)�ԋT�V��}��u����N��	J�6�6�i8$��ũ@�&�d�\��4�e�Q��1I�=�rs��_0��S�����a�K�-=Y$��Z�l��3��=9o��Akw��yp�-H���s ���8��1�(��DrH��A�p�I�z�ѭ6~�0pg���.�|�k�6fu厬
*�Z��,�-Î��X]5�����$����X]���g��7Q;�!����qB��P�!W˧��)�o�D�;��o���>�Fڬ��gp�a4�P_��g�]�73'�։0k7<��p7��%�)n�fx	ܺ�1��X P��J?�6���@�����C����4�����=
���Y��1��%��raTͭ��-Yp2[@Ot�)��g_�(��dF�+����j@�hS�Ę�7ΞA�I�bH��J{2�R�jD07+�%�"Y)�_�,��-s��U��}�M��Gs�k�;ư�C,{:�k��66�`]�p64�fG�DYeU�@V��Ѣj�̭�ͯ;���K�28Ë>�N��gC�h+zG��'^&t�1�+΄~I�,bϴJ�,kņ�qln�ц�,�
aff�J��1�#���(�kOA'+b��4�04 � !��C���{��Uն�9k#�uv���B<5��IַmP�!��ӿM}������0�S2�#�H�?ըti�,A�ⲾXQj/J�R��,Q��ERi\�-kU�s���ʮ��vM�ѵ5�{td�о�я#$��fθQ�?��&0k�x�L���)�Y0}*gLc霹,�9��Ӧ�h�L���j��X�h!�/���s�~�
6,�K[V�b͂E��g[W�`��l��;׬d��5l\���˖���˗k�Z9޲ٳ�\SX3��ߒ�S��2c�h&���a�-@<�C{Mc��ax�n��6�[W�v�B���Թ#�{�dT��L4�ES��a�"��=,�4�y�2�^D��$:���E8��A�p����/�3ɜI�DD*'�
q4&�cys4:?g��ll��S�#!�+�ټ�J�H|
�R�R�:�g/����X�Z��b��/H�/�8W
��lB1����S�E���,�
V�|r9�$��D������
��JZ���))�.P����-��6�ckdQ���P����Vv䳱'�����51'�Ԝ��{�'��xVL���q��w'�?��*u�^������j���9tu/��� Ϭ�L_ ��5�5��i�Y5�ɶ���Ȣ�#���?�8�f��wD���@��Z����6�����e�;�4��m�X�@l~]��V��s�TM���6�%�@������-��VM���Wob�膀�,7<G���1�s�:r�VK�uQ����<�ɰ�1�k���>�+�ñ�*
��L�b��\͛ó����'�GplKw���u�X[	�Ys)�_&�șme"G:qx��F�0�C~��PK��E�
�HL��|�fQ�FI

�d� �`�� ֯�˕�����>7����.�x�V��ok��Mu>}�#0�X��1o��cש��t����_a�A�Y�Erh-���~��ϭ�U�)�3��E�իW<{�����߾H"�2�S�H����/Z߽/�?��������:*O?��M�)جa��R���jY��6�B�{�X�+�U\q��9�k5":�)�2�ݦ3�/_�çpT�Uר��/��Fb(�y9M�>=���ymٿ��q�LI�?��ɻ���kH�L���)�ϧ�-9~�=�'6�*���`��=ܑ{���J�'%���O���
��3���C`��Vۙ�#S�}�.X�]B	,T3�)��"u���>�&G'�	���\X�N�4,/:W��<h����$����Qg�xc'�ZH���Q�gw@J�Ǽ�"�s(o~�GŲ>o[c���P��#�X��<��n$N�d������3�֏��Lp	e��'��h/k؇mG��p9���F�-�ڒ��'1�I7��a^Y�!+:�be�a,*X��.�L��e�c,�F�@��g�|�-<���t��%V���8^R��7!M2���2��(��hDv���oׅ�-�2�eG��oK��MȮ܀�ekҤBM�W΢a��4��)pX��i%�H*Dɔ4���,/�$� m
�}r:m���"ѝA��R?��U�4 K�Dp���T���|;��+?s-agc>/�˹^%��0����(�ҁy-�aM� k��Y�*ȘVa&���c�=]�zF�0 ��!��-h�iX�9#
�3>͖q�m��nǤ���=6Ֆ�S؁ѩ��Hv`H���[k����_`�k��.�:��s�!mÍimA�8z�ah!'&��dA�V֏aS�=��gk�Dvv������S��=��)����YPׇ�ʹ3,݃n	�4w���E����`����6����Y�-Gz��<Ej7�]������∃@���W��m��޲��֥o�:ܲ�û��b�\v.]ʞ�i����)��i���n���f��Y,�:�M�y�<�.�Ƕ��ey����ڔ���毝��3پd[�e���l\��+ױ{�f��^����9�Y0m&���aŜE��������`��-r��ٷI�q�<�
��7�uK�:/g�l[��k6i�ܱj��=�6�k�:�o�̱�8�g?����#��wX�O�9��Į}ܼUKt�N.:ʙ�4�ݯ�;�����n���O��+����={8�{�Ϟ����<�t��W����5_�ɣ�7�y�"Oo��̓�?��E}��>4�6V.r�a��������pGoƺ3�3��ޑ�d�|ã��x�Gy2�+T�c�g8#\�m�Fw{ZN����>�&��u�c��?�|&6Aͬ3�#�Წ�bsF{E3�7��/��Q�.��t�g�����/=�D�@��3�)�.6�T5q���ł�tt&��M��8Wg�\�1��N�6��c�������'<�0�{��l7M.���UL��è�m�)դ�ym��6���h�fXe�ź�]-6;�q����8U#�+�w��Қx��� Ϣ�=,���2�f�r>5Us�_�
r-�fP_�̨n�T�n��.k}�T����utT�5tu.�ߗeYTW���dq���t��.�?�)O�c��8D�j�Ы��2;���@D�@֨��%M�p�-�ϖ��|�Y���N�{[�.&��}^QOb�<o���ڶ4&�N�X�?%R��<�=�дhQ����e�Z4�]�Je�I/N�2��o�ƌa���|�.�n5���l^�m����x��<oޕn��g�p�vc�-�L�	dul̩뷵B��LU"}��3��?�+K��b�_�)���{�\)QӘ)?�
�>�����l}����/�ii�J�F��T���V�H�~S��ׅ��V�Ih�*DU���~���Y����#�hӣFW�C`�z�C䴚��8{�>ӮK5����A������%UG�/.p��hv�,ˮ���p�(���޳^|L�ey��g�5d��&TjS
?)���",�;�G���MԼ���)E�ڙT�k.����^�A��}A���<u�߾|B9�~*����E�j��PJ��J�K�V�8��i��w��V��	��N��+kgW2����d�p:���o�r;_6��_��ysN9���7��^��q����\���Amg��:Q�����5������6��kJ5����%�[kjL��>""�޴�@V:T�J��$�۸R>� ��u�C�4/V�޵�ѧMo�vB�ZMȊ�G��Iz�$�Hx�74"V� �ؘtKkR��	�L��@ �H���N��6�#�VR�=x#��a�)̚��9��;ks�,b�y�9�2���&1e�4Y�ȴᓘ<`#:֮�w۞��6�@���4H�U����ҤD�1�z<�2�rc2lYX3���Ӹ0�"we�r{C�k�ZÕ�p@����ܞR�#=�A�+�0��$��;��t�6���%},�'��'ؘn��t��K�%�%�bA�P+�ǖ^�V���{�)��M�nH�h3��5�g�1�#��z=I��^�y4�S�7&Ŏ��j�����]$�������L)��e�y��6������Q�7����$�ˆ�~,j�Δjn,�@{���v�r����nV���j����0R�&�SŹ2�+'�*���Ύ�XKkh����k���p�e`�ly_�X6}����o���E>�~r���;>�xΧW/�Zо?�����R�z��?޽���|}�\�_���c�߻��kxr�"�����;�yt��w������z͏����-o�����w��?��Wڈ������+)I��)�!��yz����s��������?%����?���&gn����^2�b�$���-�߼�e�wɘ���J|����k�C�^u^�9�u���J/'�=���]��$�J��?>����_�xÎ�(�/.�N�����%V}+cE�uF���̈W�3�5(�q�.\ⰟR��I��#DE���s�.f������J/R�ձ��K��ZV�-�D��e��v�Vm��OI-+���?f�1Ԭ:abk��S,H�s�Fz���SBL��12�ߦ!��b���d��E����FTlq�Jw���&����\`˺�}�C�[�Ʋ�ul:����-���`"��-ob��z�d٬�=L[�4�����
$�7͉,�6$ ��V�s ��-t���VWO��׿+��տ�A�Q�;6�F�N��f�~�$]��ս�|�$�)0�% �9Te	f	��Ы���j��CW� �
�0)}���8'��V��?0��W�p�TE.�����8N�D�3+3.��y^,WW���JAxֈ��S�bq|��^��ueL�.t��I��ɮ^��M�ҾQʤ%Q,5�U\��?���Jr�|M.�������ex�1����%�s��&f�\1�qĖ�H���x[l��D�P����Wv��?�����%�RAq�r�j�^���j�4�S��s��ML�G>���Tّ�9>5_����c�L\ElVO�2�Z�1!3E���R]spZ)Ks��C�t�Y����p/��sjq��h��Eiפ�r-���\��[939�ʳ���ر���%p�X^�<(ēW�xK&�?�c݉*�V��U���m�y���bk�ju�ɔ���0���"Ԅ�
 �/���i;V�z���.�E���&�#�Ũ��Ӝz��}��/��!g�\T���<���Z�Wy���:_�!Q;�K�ӕL�P&�2�ԕ~bl'�:�BJ�[t6Ȼd�f);P���<��ѳ5�#��J�!S�ۛbgl�}���g���b����X����� �.�9[;������v��/����]�iG�݈�̇w`�D�u�
P��`%�up�C��O-̌02ΣM�o��'g��<XJ	�M��斴�c����6S|�T�%&"6��$b�y��"9_��J�]���t
�g��BJ�t
D�R(.#g]lA)��#:4�ĈDR�
��Ͳ��C��i�f�.Ŝz��V%�A)V�V֓5���ߧ'U�����؜ɗÍ�:���B�ݫ����x?�
G��J�v6�eC�(�T
`v	O��efqO���0��C
:1���
�2\4 ֚���Mt���6I�eDaGF�;0��c��1��3sk���~�Ű�E<;�'s�I./��)Y�\ؐ+�m�\��pH��\��Vp�����Q���qof*�FŲ�K�����'�jz2����7lMYo[R��r����kyO�������`.��Ts:�-)�wo,q���t`˪i߳�o�ՔD94���Rߘ��d��]���:Y�:�ȷ����n�C���R2{����Z	4�������4k��6��Q��ʁ�f�U.��.T:�����(���t����>�V��Hv��r�U��Z��V��yJ�����sY�G��}���\ U��,%w��W?^p��~�Ԫ���;�.�;8�ꎟ�#���;yj�I����0'_½�	��HT~R��Hp!�{0�^�󍠠G���T�\��w2z�"���t�t��z����CA?�]����K���6�q�g�]�Ir �=�4�`J�DKHaO?J��*iJ:U���O�W)��$y�P8(�Tg?�G$P3o�|�b���JFp�p��^fSF�����=|2�M:Q�J6�w&$s&�7�� �-���$���t7���qm~X�������g�͑,��=�O�x�<�{��86>�ɡI��[�í�y9FN���ޭ.���*��i�W�+����k˫85��s�+�k84��]���6��c�˸���S��8���}�Em�m�Kش����<�<��a�檬���0�{��4�e�F���k��0�6�֨�>�Tل���j�Ǽ�Z���ކn�پ�{���Ԋ��*W
	"�Zh�w.^��U�㹊\=W��S�)Z: ǰ4��(y��L�۟-�ɮP��Ukлq��oIˬ�O��dQg�6�d��X�/ƥ�<��8�_����j|�&��T`چT*�%���P�:�b�~��яyK��P
m�|�~�����W���<�l[
�^<S�yb����	٨�����_�'�7b����ج�go�r�

6@x�vDg�"�Fc��eQ��@^M�g5&�zÜ���k�|�5�[��6�6�X9���/�iע�K���Z����9M�ܴ���5����4O�[��A���F��݂��3)� ׂ��$ƯTe<���#�"�%jb_�	��;�f�JN=��{�K�
��+�{Z��D���s�Z���ԍ��w���C�[Q�R9�V�	�~��I-���������5��D�k[����/������*oA��T �TU|3�i۬l,�������Q����8��:X�j��K�\Ye`��	G����Fg[
���4k���%�zFD��Lpx��ѸGFI�� WB����%�:�/�`�|}Ő�i��	��",H �-��0������OtLA>��8�	�p��Y�����N�x{�CzbEf����J����"(D .��b
��������d�
i��"��H�~��{��Dbx��xKf�����g�bؕ���۹�b�≩\��d\��.XX9`gጳ��6S���5���J��bG�p7�bt�H�Vddi�ف9�Ѣ G���*<��ɓ�Ux��?�ԅc��^}8!���6V�뺚|\^�������\�Z�3c��_,��D��c4��F�C�u$[����e�ZG��U${��s�W~N�΅1�\�\��s��lIe~_U�7j3T|ۣ@N�� �I���|78�]�%>��f�}K^�u�>�O��5�L�P��ln��1��5C�XڗAi����Ne{��ْ��D��+~8�[`ah���=N�؛�346����or����Ņ5�jT��nؘ�`��G��3ϣ���Cz���э||}K����7��!���*�r���-X*��-d�.k�,I���/�e���v4���f�d�jQ~�4�ɕ��D�S�+��9�
�]s��������g�E�f�T
-3P�ͱ)�������1\�@��.�i�
�iM=Z�Meꏜ��:Tf���:�
��J���]�������#�Y2m��f�I�3�q#�2l�(�O����<f:��p�bfL���YK�m��.\��+;{�<fL�˸�3$C^��YK5b2s�lb��KlX��S�2b��X��+Y�d=��ob��̝��Y��1c�2���Ă�Y�p-�b��_�n;K�� ���E��?cKn`���̔4K�J����X�Y"�n\��u�W�B��`�|6,��ڥ�X�P��>���ֶϙ(�:e)GL�O���jѓ{P�JW���Er�nDjOxzg�:���B�(����$��9�5��[�����vI���B����[j���+�?�����{��;c�E��^tn��Qb>���[~.E���>�b��0�Z�9_�O��Y����Um.~��Q�E^5�`�&��Kp-�������z;dy~5V�S}�h%~U6�Wu-^5��Qk�u��^e��7��2�+ԖJ��]�"z���\�o�Ws3��4�F��`l����S@�H��MBK�Q���T��k��޽�ԥ3}���M�,�Ԯ-�3�K+2+�XQ'*U3�G?#�o���E_�>�ݷ�<|�ɶc5i�?��jy�N�çdI�6+��K-x��o�aמ:�:9Us���g��W�����Wʅ�\�u�%T���1�?�/7�c�ڼ���h��}�r���B�b�nE}�G�<���u�k<��j-�֐�j���\�(��ʵ�[%����i�Z1���4 ��X۴�x���VӖ���(�'�俺�yB�?Kߟ?������<Ѐ-���d{2�� {p	b+e`��mRm�E���J�[�n%��P�6V%j���l��+yrXU��̼fT���rQ�t?�?/27�u��?y���?�ț7����Y{1�gp��#��CryL�KaU@ O�]rv���)y��Ѧ-�/&��Rۄ�X��<*C//���i�p��v��Lr��+lX+��Mg�)+_�9�PE�?����bl!ZU�ͨ��X6i6Kg/d��,�����3��8~�1�ɽŘ��^#�m(�;�g`��L�;��'hF�Y�<�i&j͠s��b�ؙ�8����d��)�2�q}3}�0��Ĕ�#�;h���f��U��x�\��_Ȥ���X����ߖ1g�,��Ƭ�Y<q+�-f�1��=�iC'�h�\��ʡX;j13��eB�!��:���1�}o����6�Ա7m�[Ӹqc�6jJ�f-iQ�	��֥Y����jF�Zu�[�:Y�jШBM�,K��I4��Y>7�Tc\�0��aL!7ƥ�0�l �j�����^	��ՙ���8�W���q_%��&/��i)��*�y�� ���p�5�7��Ά�ٰG�[��	lm;����M�d�mGd��o�����X���d��SnU>m����y��27f��ڌ�\��3M��!�����Va,��+�g~u_&��dDQw�t�s��C��s�����@p��Q�1��R��p���M���� �|��*��_
���Q6-���H����6��#/{�w����u�Z�7�E�$ �;av��H�I�){�ٜ��0�A����>~|��o���J�f�y�����$������OZ���k s���j�䨿V�}���`9������?�+�s}��V���y_�+�(b�AiA U�/�:�jm
.��uʮ���r�_5(Ů�9_˹��x�˗Oy��%�޿�����Z2�g�=�P��\����k��jr3,U(}�������Y9��3�k�jv/Z�v�KV�j�rvn���5[ٹn7G���c[���Kvj>�.-���5��� ������-\Z��kvsn�.�.�¡�'8��4ۧ�������|����p�	�8͕U{��f?W������v�[����}�X�]���r���sn�6.����i�89oǖ��������#�W�o�r�\���80a	;F�aÀ)�=O�V�/��O`���7�n{�Uɦ}��4ɨJݴJ�J)G��$
�Ƒ�E
��Qxڅ�j����6�X��`a��Q ��~�����K��:#_t����4=�`t�A��LB02���4�p$�7�D�2
=�(t"�-����#�]~�;N���8=�tn�\�s�*�nE�:�"y��ԯ&��1�-�i@y��kh2��Ep�F�ڋ�b����9�e��θķ�9#��kc�P��U0���Uhu\����_�����1:ځ�!�|��Ҋ�1��5��me��Gva%q����W�-$���btkܖ�}{3�w�u�C�ƭ�P�&�Z�`B��*�B�T�dFv;3��r�P�.����LX�B���L�'�!�s�+�6+ʕ-�˪ɇoe��!/^���E<s�__h��?��W�
xJ�[R�'��~u�)��x��Sΐ?x��G���V��/p�
qS��PV��W���������J޺��)W����	+]����4 �R�*fV�QUjT�*�IE0�+DR����ח��.���w Omȅ<��_U���f����Ђ�≯�B��5�-S��5E�pMOǫhQ����JE�
�&�|5�g�S)�|%�^���I��aU�J�?���5�z�J�Z��������߅�^�ܦ$����֤:H����v��P�z�)�՜Z�/���S3\����R���^��
��fZU�瘐�eh�Q�xxS�՛qa�Y��4S{��Ykj��9�I����\qf��������V�~Ӡv�������l�1��������9i���۴}��je�Nv�w���9�w���<�,�F#�����H�F�}�n����V���񳰍z�W�nMZ������i�K������maQ��XP�s��`n~,�k��eݱ��`��1
+;���ñ�|0����#���0,o�+:��
sVu�u{ak�>� @��c0�C��-��-�bM� � �m3�:���~�N�vV�Ί��Z1�kFas��b���}��� ��4�{�������ֶ�%]������՘��3s�cz^[L+����֘ZT��%m1:�C1 .O�#���^����a)h��"+G$j�#M[ݼ�06�c�M��O�����_C�1/�
k
m����;Z��W���3��hi4^�N��aO&p8�@�w���b7R/��J���L:ہ��t�#�$�9�7�0�W��G�[��	߭�ëeYb�[^b���8���Cq��7v��v��U�7k�,�¢<K�ΰ��S	�COoT9ȡ�F�frH5�E��<µ�*wŖb�A��-a�\�-�a '�����g��
�!w}U�+�~%�o��B�M�B�Ic�R�/ۨdC���7��M��ѫs9�m���/��O�$0��T��?I���d��wx��^�z�wo����������[�'O����kx��6��|�����ś'x�����}`Pz.��iP>8�~}#�?�
>�Ľ�7p��Ma�{x�¼�g������B��w�P2@J����"d{W+^M��+]0$�J?��_�x��߾*��/��νK�z��]��\���w�n߹Di�#��q/_="�{F��N���v)�8/^�~Ba���<��}'�x��V.���٭�:2�Yh����I�hOI��,tN�G���*�ؒN��T��>��g����)8b��cv�8l��ݖ18萀=�!�ퟅ1e��g����L{�뚆���t\8����C�d�4���:l��.I�b���B�)�=_���j�m��i�����Q�f@~����[�±�([L���0+4��Z++5�1_�c,1�����z�����-Z��D��	�[�!LF�͔��D���è���C����z=h�T��B�:�-�5��O2�������4E��MQ�~�Z5h #Ԩ>�k K�[Pg�9�R�\��Ѥa4n�L�~XN��ш�6��חEc��7hؒ$+Ը�Q�l7n����ߠ~3ԧ8�Dv=�_��r�G�����2~j�F@�Ln-h��Dv���b�Fr���۬%�4W@�
h�H��94�7����jsn�i2y22����br3i�Yu7��!:2��.H/F����N��C�bр~�1`Ft�^%TO�bVF�&��	���k��=�0x�=FL�BV�`xe����46��q0%��H�s\(&�J�/_z��T�z�G/+�����m9��v�Z���v�u�#ȓv�������W׏p�~�߻{t�	^<�������`�g��A��k�V��i�L*�CJ!���a��8�Ƥ����\[jی�%S�����o(~�q�ap8
��1�OW�;}����K��ǽR�<~?��?��g��݀V���^�{(�
z�&��"ӡ� oh����R��F(~p�X�_-<ɭa���l��gP|>1z'9#����͓��nx�'!O6U-�q�x�U�~�x��o?Bi�q�L��G�|c��=�ޡh��u?J+O�7���sJ64< k�u7?41����)\��Qid�9��X.k�%MU��@oG3l�~w��8����Ԡ�#�^h��:�X<|*�����IX��M!X���־g�>ڎ��t�׵CG��4rE_#71�� 7񻛑:�ء��#�i�`�Q �j�c����Zc�9�5��`S_5��}sѳ�(cW3p� m{�Q�Dw%s�%���b�����c��;�h:b��&��`��'�;`��=ƙ9c��a�!�vB�u�bV7A?m3tW3A7��E��I�ݴm�Y�ԭP.��j��e�e#T(�J�%*��n��%�r�"��X9D�j!���j�mA�	�j?���*z�[�>��tP㡁��Tḫa��2&E�cn������aCK���}}�qd�=Nw����y���\��3#q�咮Lƥ��29�����(O\���c|qr��sÑ�8�����aGW�l���X_d�e�fX�j�9	������Z쯊ޞ��謀{y��!�XIzr�іE�zSx)6�S���j\f�����~�-�8h��6n����l��A�a}�5��F?A姟�X�����@'$C~I<W!�VjD�U��䟿��	��=Q:���6:�+ŌYCq��^|��!��}��o�����O}x�o^<��Gw���\8{�~>�+�����s�{�
=$�w�/�Ӈp��^\�rZ,v��9Ig/�<"(��^��S�'�oS�{O�]�3ۯ	
_��/�;��q\�zF��+P<xr7��ɳp��!ھHvA@��ۗq��iܥ�<��7��H<��t>�Ǐ����_�y &>��iY�?��?����G���Ν�k���y�x>�C���y��ݻ,�/]<)����k�q��BpȐȓ+?xtMls<x��ga���qb��>����[A%���PA����Y����(��Ƥ*$
]��P�s�~^H��U7��B�E'�U��N��5���(�mc��6�Sq��L�.�i�Q8h�&!ج�N����X����m�]zA�e�����n%@o�Y ��Ē����[-���$�"��(;	�ZGb��?A�V�xc�E$�Q��b�nV���0l4	�
� ̦�j�_Ct\1��UQ&o���zHj�� %��[syX7��i��ЗQ�VEh6V��Y��^3�&�^�y:Y<Z݂:5MI�=����c�xO�ܰ6�|���=Wvo.S����$>��0�-G����m���~�S�n3��m>F����Ȑݔ�qi��'�bř��O�����W5$�'wT�a�=+G�[���ۍ���W�)A��_���*A^��@3���B+rӭ�EK� '>��v���#�p�l?+Ŭ�=1��0�8�;u�h�O	O�X�0��G�7D��DP��`j� ?��ï�5��*a������еZ�.���x�K>����.X�7��������<��5�6�o�P�
Zҹz��
I�@��Ŀdt^��0�c*���v�>�}W;����g�o=B�%�a��V$���τut:�ᚖ��4��=i�	������8"��1�ahh��^�.+ìa1���V�>S|9?��?<��>f`}�D�#����Y3U�
J^1Јʆiz6l�2`����`hDC5<��	z��	OKo�Ǧ@?)�	ep(ꃚI+���M<�La���dMIxT.����g>e�D�Yx�W���xV/HN����x~G�Ł�K�T\����_��/��:z��  ��"�m���N��s��g(T|$r�.ED���-,��_ T�]���	y'[�ؚ���U�^�i�*����V6Q˅���^�S�a%�!۠l�H�pT�5���5&�]c�c�W(viZ���Y����&����]���zn��Be	`�k�?��%�%4��h$��,][�'��E�
ES,h����T1MN��c��&�ȩb����y&�W�DLS��|��y�����IM0��.�*�a���������&�7��$Y]LQ$X�U��J�R	Ú4�(���Me1]V��*R�J��R34�0A�@L�0�����Qo�=�J;7P@�v�sVRO9�^C�Q�C��LꡦR�7�ܣ�C� �a6���O��߰1��5B�l��D��

tP�@��
Z�*��\m��޲:۵D����o|�&&F�aV�&f�aY�V�am�)��ak+kl,���R+lkm�5�F�n"�2� ��M��w��	��1� nF��X�bb���ʣ��<:��D;%���C��"rL�j��Xyj� �kw�&�o�6͛�˴i�4k"&�6��E�߱�<��N�j �����n V�u��d[R��:�I�(�5h�FM�G0�+'K0��ͨq�� �)��1�M��e̴[��z3j	�AkF�UC:������1g�?�����[�^������ݻ{���^��C�� W�������ȡ}8tp/vnߌ];��̩#�x�$N݋c�w�ɍy��#�w���}@�\���/�����Ť�O�� �@� ߽{	�.��� ��u����e��0u��9�:s@�?~f?�؊��6���=8w�0�s�ۅ����~&;!t�
"A����	�A���#�7�ٕ˧��7�s|�߹$���9~t.�?����	�7�]���։s=�KL��q�t^rNN+��'w�4��p�<_�q�O���#q��l^��KKQ�@p�S�.i�葕��YB=sr�%=�2s1��
s�������� ,i?�z�Ö�3�q�T��1��L����6d:V���Sb��EX�oNLZ�cfcjy{�*¦��qx�bl9G&/�Xw�^�CӖ�䢍�;c96����WcόX9dVS�������n���s�����4��avN_���fcA�	��s,V���b�c~�ј־�v�z�O^9:��}l�}b���������	&�0ֲ�u"ը3�$�5�cT[�A��6���ϚQ�[�iK4m��f��A����m�H������\��t�4�CK�h޸�6�Q�Ɛ���ՠAc4k"�f���	u��ӽ��K��MќG	��?����?5�uoB�k��b�B}�:��1�Q'�'���fߨ>Ջ���z�݄�Culܠ	��}ߘ��������8�ɡ^35�樤8>�� ȫP������uD}Uu���!*8y���^�S���Sqx�"l=�GNîK�s�,�2����XQ^�1ř�uԁ6շ
��s���DG�*#	�U%p*͇~|���`����pl�ӏZ���� 
G: 0��f�ìM����:\���_	��	g����kj����$�."a0)c��E����r�{xa~�C�ʆDf����7��J���d�|�n>F��p-���6p�o��B�%�
���˄[&�NɁe2�_Z��=&�A���yֳ�zj2O����zc�_.�XH'	����;y<��tʐ'������So���X�`=|r*��'ZD�z	��
��!mkDG@-"��	PJ�zH
�"R�KP��\�E��4��F���q��'��s8�DD�q�1��Yyx�uȓHR�<N��8/K�����a'���$&�;�^A�~a�
�����C�7*��P�
6_��A��/�AP�60�����T��`E;3h�#��#l�1O�
�dԱ��"�6Q��fZ�'�+߭���*�b�������jt3[��b����;n:�{�DK�&�9�S�n����d1�@�{uTɩ�TA%�CJZ�C@։����6��顟�!�(h`��F�kb\5L'��H፣^�x;��
�BS�t���Q���jbά�����Y:Ƙ�n�IJz��j���映m��r��U�1��m��>��`���F���j�M@;Z^��1��:�(jc8ŏ���n�Z&�D��M�L��uV5DG%}�S�E5�4��5Q���\
+G]Yn
m'�i!�*�pU5���D���#��N�#��m@2�D��2�,t�l��d=%d�tZ"����9��Qf�ef2��$�tPDO��<=T0�_�}41�O��0�SC|51�G}��o��Q�����Q56
(��G��,�!N�>�t X�>4����ξ���I N�	U�M�߼�x�jL׊����#̔��_l�(�o%Uڧ3EUX(k�I��44`�!����aAy��}VJj�&�+(�BE	-[�DE�J�8��j!9��LQY�"�XY
�����\S$�Re�q	޿��׏���#8{n7N�\�x�Õk'��χq�����8q� ��Ia�<q�����^9�S@��@t����}B����wRX���\�v���8ǥ��q��	�=����Ǟ�q`�z�=�G�̩��3?S��w߁-ؽw3���Lqچ=;7b�V��}�p���'�:�_  �*���}��y�ӧ�����x���]����"Ml�d9���<{wm��=[����/���5�xz�����E>/�R��O���%�t�(MKf�G�R��4��+�R�),B�B�~�%��C�+0�S7l]��V����[��Q=|���V/ۅes�b�­�3u)��^��a��UX61�._�[�`P���wV.]��;c��=ض� V�-���o��e�1k�JL����l�܅�0j�D�N6�f����k1s�L6�����1{�2�ǘQ��W����¤ɳ1n�L>ݺ�E��}0��0:c�NA�n�*���HJ/@PH2�]�`i�[��{���Z:�� �SR1RV3���)���BY2T�5�N��O��nl�H��O
To�6Wj)���B��E3e�2��fJh�\	�d$��*GZM��Tu�8�/Y4j"��MZ֊�KŏSYɏLE4�S6?n���i!9�L1�5k�9���7h�	B�4m��T��Pg�u��خG �sc�	y?�ǵ/�M�����Sh+{;�{� �?��(�MŐVm���P,��+;����C���4������C={c}�^�����1h���3d���Dn�1�0N��eNtb��M�p��yN������.ǜ��/��E�3��
ժ���=Gp��;��B�hI|P�-��<j�k!�{$��Z�cV�*)�}����<<;���Y�����a���#V�@z�Ip.���RXe��9�
��\�K��[&�:g����T�5���	P��"���,}������0}�H�K�*#Gܙ�D�=��G�ǐG	g�c���x�K{������y�Ztܟ�.
���!���4�%g@'&Z�q�$bWI�ZX���E;&��/��q0�ޕbl+hduEh����4=z�Wt�~�,r���z|�ɂ�8N__H��k��aH`Q"ix,�n�"��'o���#�m?�ض����4腧����$��;E�1��߲6�� ��h��A��-�������Έ�pF7/̳v���Z��Y0m�J��?�\�Z�c��&�<=�w�V5�z2Т����-��=�fb.��.��k���a���d��M��	�
	h�M��cl�#k�2&ws{�٢�����ptA��:8����':z���;zY����/�����g �{��a�o8���w��E��K ���b�w<�x�aA�0�(�D/�a��B_�X=z+�;Fg�Of1�aX~+��/�جbK�È�2�O/F��B��,E��RtM�C��V�S�nIE���Q�h��6��h�����h����xTE%�5��е����@${�#�;��QH��"�'�^�H��G��� �gk����KO��P��>*r�
�K�)��e�-�~�M�"+��Q-�)�$]E�i�D�nK$�+ FWN���Bud��jM�.�fpTl {�����	-�P�'�5m ��)� �M��ic(�4�B�PnҰ�1�ZsY�((A� L� N� O��M������TR�����&�x��\uh����~���,#5�?�C^"Ζ ���^�:B��'�&p�Ԇ��<u����t������aG�l4�ڠ)�]��t�d\:s �N���:£p�p��^><w�d�������3x��^����Oo�Ѷ�����u����o�eä#a<:�˅�x�!��9��WN
�%��7���ޱ�`c&֮�#`�ݡ�� �;���#z�_::�#���+����m\�t��sG������0�ݾuQ@�tԎG��ܾJ�{�S<H7����_�ͫp��eܻuU<�����/�,t��a~	�����g���O�<,@�왣8rh���}{�	���}����|�,�jW.Y)�$�[�cH�R������j�Q���w[��h#��m:aր�ٹ?*������%U�jP����:!#�5�t�U�v`�Љ❬`j�����t�8��4,e�E(-@�WRܒ�闅d�d�;F �5i��H�C�c ���e�8��zD!���6~HvCj@�In�H��D���� -��>QH�D��?B(�U>��p�L��H����i	' �:#(8��w����+�-�addshhI�m-]�U�X|ѯ��Ym��S�N����Zʫ�y:YU((�@��c(*
5k����)nD�&�5!#���M� G�aC3'���T�I35�8�=D�d���Y
���\�V|EE}a�o>GK9]�PG�ᯩ<��W5�k	U(�=�D�Cy�ͨ��B^2-e�D�4�!�k,��jHuN=9yh�k  﩮6(r@S9<׷D9��(�DKSk|DS{���T�&���k ������$� �Pu�=[̊�Ŧ^ݰ�cg��zZ����j`�f^P
�VT�%¡ŀ(��# ?��RU����hKW�x�P�\ ��x�w@����r�&�?~'8�x�G��=��0  O���U�ը���	tϮ!> �12+�/����#hFAn�>���@ۙ��V=:��`��Fy�Ԏ9gV�����2J��U����#��
�%���F�DP��#M�5�C�թ'����U�]���K�,q�:@b�@J֏L-��~�\)�8�l~y�֭�����9ߵ
��@'2��c�.y$����$hE$	�ӎN�QR6�ҡ	��8���C/���m����mG���mX��ܠ~M���˒̕��q�Ҹ��EI��8M����&�.����t&Q��~��e[�]��~	h���,h~�c�3�Hۚ10�t�洂w�*�>�c�B����/ZЅ+oe//T�8c��#��Z`V�f�=���[��R���?���e�_E��u�z���-�SSh�9��`ưq80q��D�5)�4Q�bE5L��Ŝ�4"��E��t�L@�\�&pJ�A��\����&"N<�XZ�aU�ۦ��t��N}0��+Ɨw���&��i�;f͢^�n�0�G,�?
����S1����:S�Ō��0�k_���Sz�Ŕ�0�O�NF��m�:��ٕhߪz��!]bl�a��c0�w�~��su7�k�	�;�,�9qy���:��w��H�rH
�C�Z�o0���P�	x�u�yz�?���	�p�t��ϡg'S;8[��� �����0�Ӂ��"t嚋y��2�M%#g�(�*=������SCS�W�z�?�=�`���[=�կC���wݚ�I��UՃ�
���|��oI��R���5&�bT�I�� ӠSXM�Ӝ�M�7K��6��{��o�&?II��#���?-e�A�ia����)x�_��c�Ѭ��rB��d�(+s�h'GD8�#���VB�v�mM`lj"jg� �@X)i�YO�ј4�z�����ѓ<���� �Pv��1�%�㑾�W���x��ׁ�������9~TI�v� ,�}�����q�?{H��<�[���m���c�w
�۹y��4,[8[7,��]�c�J�۷n��=�q��^1�x���;sPw��6�wo�#y<�v��N1��ڿo��>~�ʣw}���QI�����c��9X�hvl]OaP;��;�a��%X�r1����V��a�Uؽ}#V.[��3&a��1|�X�v��7v���#�`@�^�Ю��>2�/jZ!3&�
20�CVaHe�V�cp�J!��a�	���TV���з��`-v
�ph��[Dh� R�~ʶ��t@NL>6�ށ����PQ��U��XQJ�S�D`#mx�S�O=���/���!B��--�C����T�'�E�@��9b-���ͩsA��o}eD*� J�����Ҁ��*����a/ym�;"���f�0��jYO�9+�!�/�����
����M��� �ۺ:�0$p��5���!4���N�*��AI��M�D���m$��rj��|q����#}-�uɯ>����/�6551�#�t-����n%-S�TՃ*������i�S�!�S#�R�5iFP&����M	�����2P�5ׂ\s<E�TK�+�C^Q�V
JjP�NKAQ*��"�J�zP�ҥ�����"��7o
�\6���u��,��=��$ȓ�#]c�f�B�:����!�͈͠@1Z'e�"!���Q��.�>l�E&�ب�}F^�iP/�Ύ����2L�OC��=t� cj�fn�P��E�0��!���vl�bSa��~���=���8y&]G�����͆fd	�òa�Z�xj���߈]�/�.���;1 ��%X�$������w���xH
x�ѡ����1?�Qߋ	��.<|��;O w���~fO���qz��a�TǌVp�*�Gv+x��'��t���"*���`_Y���G@�7ɕ5�8t$��텅�ا팵���:k�$��D�@ޟϬ�Ү�A�J����Xl�E*zX��#Ơ�}?"�4��GS"mՈxv�Y0� �&�ӎ"E&C-,���ЈɀzR\t���S������f����Xx�.�����&�h�N=���[1���'�6����2������
��^�܉IV��#�ͷ���Q8ll2*���@��X(PŧA=V;�گ�g���BxV.pw?����׬�gk�&���H���$�,��Ǫ��X�X;�5��z�����&j��	�;A�
/�A��tc��ZKs+L9	g�,ņ�L�5���ژhm���)�U�C�K�>4	e>�(��-$���($�)��B����Q�*���dD$"�z�m2KQ�Y�6Y�Q�����$�#?>���1H�BA|:j��<�5���$�r#r�Ky���<�R��L���x{d{G�� 4�-a�^B��+��qC��3�I>��p5v���;܍�`�l g3�Q�f�f k���HYf�:0W��]�$�	tuU��L��1��M��R�~���*p�;P��Y�
uYu��*)�*@��,�6�ĩ��A�Y(�4!���l&��͠�LN���ﵱ�5�*��A K�`L@K�q=(�H$O�
M닗��%j^]BM�		��ȍA�'�V�/�4Z�@L|�ڌl:�m��N�������o��<TdZ���W%��PUP�����lK:��)]���bDO�*Me1�)�J�T�.�D��ܴ1��=P���?��{"�����FId�#BQ���$T�%Q�G!/*��h��
��&*)�hW��3�bǞMس;�o݈��V`��Uز~)�ـ��w����8t`A�f�:�'�o����ph?�׮;�ţS�޹}�p?rp� ��6c��UH�����uK�c�J��q�"�]1�W-���s�f�,:�b�ؼ��B<V^�j֯_H�˄��\/��m�w�Z�ݻ7`Ł�{�&�ܱ�����k�����X��f�bڷY���Y�'��̩�|�<lݸ{vl&�[���)N+a��ebߢ�3�`�T,�7Ml3�M?
cG!�$@o����&����h����6�F�Ĩ!1�gW����F��	C1� L�������}��������~}1k�@�<�����cF����^F��h�����a��*V�T�D�W8�_��#�#��=-\�[�m�t�]��!�j���Z� 8a�FV�U��K�=U��QN=	���裋�5�&������o�^z�h���
ڟI�}��zd�Z �:�a�'h	ҤN������c����aT�������)��p�t��C�`�������Ҡ�B�ښ�PW5����Ս�i��umaf�	C^"��-��v���jNP�i`e-s��-Y,eM�Tф��4M�kaUCChȰx[V]C�z�BE͔�!��)��R�ք�[9���~U�zNIM-u�BN2��Ѩ���UUL��o�*3�Sbcu3�+�msk���i�f����)d���W׆�5����_���
i�������1Ѐ!�9��i��k��A��vv6�q��;�9�	(�KBijR�"	����m�'jw�1.,윱T���L1�@s5];��0���N�0�0<�!Cm�bx��w�0(��1p�ɀIVtb|���y���Ë���Kv��B\��<�a[�b� :�٥��1m�-Ă��p��}����>Og�!��y�v�_��l\,���[�
6b����shP0zp<[�r�y�f������a8�;�&�v)�pH)&N(p�W�x��p�FRǮ����E�����&�!��<��K���6���*�$��v�e�4��ՙK�$���!�����!�A�z+7l��s������>�QXRywO�s�@c�P��$�:�H��H|����B3$:D�yZ�	Ѝ$X�ˀvb!TRj���F]�e<��X�9{���7xA��C�b���TG"~u�������		���ܯ={���/�f�b�W�Fx���	LS�O[��/:~'�Šg�RPy�՝�0�Ċ�N�Pp��O���DBP�x$:��
+Z(bSU��Įfj�F����5�O� �e��<�ۤd����~jSkL:��-�2�tl7p�������B7YeX� �<g$�9#���T����#�`*��i��b;��C�$�L������@���&�P3��;p�Z����ԫ寃}���g?C{�9���^T:k���	���x�{�0��lEМ��x� )>!��A6���Y�;N�GIb�c������f�� )0��Aԫ	�FRH�}���xO?D�#ԕ �-���s!7wD�Z��B�~q�F����=���
7[;�XR#a�?k��S^�P%f`J?�爳3 ��Ӈ��6,�x^9-�S��DCK��f��H %}U9���0�P����$�V���:4�&G��(-��`��+-5�~�Kg��Ja�B_EY�.����dy;Km��j�F[6�z��҇�����`kbL�5���1l�a�ogS�X��������Q�.Ɩ�RZIN�����Fev�w�@��<L���:WbP�Vж5&���#b��X9mV���5�����1{���5Kf�ì�C1}�̞=K��������X<�V.Ī%����wnYA���@n�mY.���AK[k�e�!����}�n��k��0�P��`�m����}�v�Am3��}5vo[Eи��]�ի�b��!r�]�qp����3���#u<r�����<���o[[�>����E���G�������X<b�#wz���������������Q?�����q�7��|Z'�f���}�؟���J �	���(�v���]kq��h��e�E��
ٺG���1Ӄ�'��¥#�pf�,���V� �q��6K/l���j#7,�	Ĝ�|\���FO�T�wPq�s ��xc�W�{����ξ���m��K`����=to�u�.[p��a���~� �s��p�s�Q��p	�r����	�t߅��!��qVVH��(��-� �*�!��kŠ��k("�3b�`_8������v��յ`��m-�MP��c#�GMM�ab�}'h�����v�0����<`d�c!e];(T� �$ n�neU1���iu�7�t�M�J:�����E���h���>�7j��KaYR����(,uM�al�
K7���CÀέmO h
Y%s��P�ad�#o������Z.0�v�����mj�U5(��ĺC�ڎ��j�V0w����� a^�u����Ѯ^c<6��S	���77���)�C��VTo�;������)$�*N�F|l4��̭M⃂�$��L��`L�q�l3�!ȞN������C1-(	.�������#��7T����8XQ�Ҿ(�i1���GvE:]�UԂ���b�~G���>2@�7g�Q��\f�,�-�2�X�%#&b���Xv�g�zO?�Z�!����~�|H!����J��"�oh����?���CLY�]g�AҀi�6v�z�,�-ls��6�n)y�NχOV�x<�#x�EU.o����o]��V��m��BX�fB�?��=��x$�VaF���7j4Τdb-q�V�<;l6���y+$ ����!��p��<v�T�#�SKc��V�b+]���q����BzA>Ԣ���'-�SS`����Rإe�($�~I0�L����j����2bS����l�R�njk�Wÿ�0�O^���`۹�x���P&ð&;����a(��q��$~z���L�s9�����;̓+a]$C��B?:�~1P�eB���ĄVI���Ϯ��[�G��	p�/�A^C�(:y�$(Ia�F��rcg�T��J9l�S�ޖZ�%���U�E���	�L��6+�!��O0n$'�<�ǭ����p�p�4��=���L7oy��;5������#��h� �v��Kb&j��P��aI���B;Jo�o8���QL����xį0 �ZUTNm�R��3�T!T�x��`���	��n(s�B��
�\P��{G�{�<$����/�ҊЭ���zb����6|f���CFa����>b��d�0����a�1�_?���;�@��.�,k���jT�V�&�:䖠g~9:%�w��&d�Gr��ģU85Qa�BYh(ZQ�R�����!?$�A�(�)�5��Q�v�D�=A��=��,�ca/���^W��C�km�4�j�l�|)�T�%�UZ@O�)��Z�LG�f�d�����Հ���-�	 �a��H�c�y	*5��+� i��#>��U*54����zZ��ׁ�������E�|̌�cl7����.|��O���Gy����6<5u�o`� �x�Z�!���ζڡ�N���$  ��IDAT9zc��iX�p�M�%��c��Iسnl]�]�H�'0Z��;�bú�X�z6A�*��Mеm���s�q���X�r�n[�}[�V/�k	J�c϶�ػ}3���жMk�6�'�#�c�[�j>V.�%3�_=��.6?��m�cp��{���ޭ�wٳ;7-�p�`��I`�y����ظq1��؈�;��xp|���m'��ǴR1�m�B��u�!O
x�}{�Pڗc��cdx�+X��ZH?��/i�_����Ƀ�=@~T,}�P������GHG��h��-B��n��픇[֊8�޽;v��Ν+��::��nā}�c�lܿ�N�����94����T�g�mq�����q�-먎�3v!�w����8C����1�����	8M�v�9��~v��H����]�-�q��7�p�%7\q�1?���Q0��e8�K�A�x�4�G������j�tꄕ�١�ň�L��ĨD��Ŷ�#��� ��SQH��dd��0������O�:���,,�ao	'��Z����'�Lal-C(�A�����P3���������:BA��*n���7��I(�(-j��sndNPT%PSw���3Z��@V�-�!����z�h�捦d�({@^Ǐ@/�f��4���a���e%�P� ]�8�&A�8-U}�|!���U����
7?�h���,���I!K��YtM�ĺ���V�a01��M(�-}ї:�w��� -Z⺱5:5W���3�(�L�C�hg�`�� ��#��_;wX,z�#�-���T�ơЃ�^���@O��!���st��ښq��(��r	rE�_4�,�QJ1�ML�SQ�hcm������+p�� j�K��C$V�Bz{����2����MʃYZ+&�,�Z�%�\����aΎ�8y�}x�{o��~� 7�>��w/p��+�x��=Ö�O���m��z��D����>�eC`Y��ٕ�ͯ�si{�Q;g��J,S�P�_�l9�?��)�@t��H�v-�mg��A/2���
ɅfsQ�*���� ��;�ꀇ�iڨb��T;Ԭ���W����~`���;o�~��O�pr�b������jةa��nxH=��˱�[W�@����<4�9����a� �b%B�u��;{ʁ���)�EF @�C?&jU����&�3Ȫ�Ev܊;��98v�6E�����=/��O�%�s%��S�r��W���V)�s��}�똵�(�/݂�^c���� �#�R�aW��|��d��:^J�!N?�nr�+�_��zr��,��wFdu/Q��.�h����NФJ(� ��\5K�7�zeln��}-5����4R�^��2����z-�R��i5#<�^�vesD�k�&J4�Ŋaql���)A7K��� W��j�����]m�����'<�;
�c�? Zhht
���b@J6)cr+0>�
�
�#<=��0<���1��|br�Wbzi&����َ���3�LKW!�l/����b���l�gg�v�%޾(	su�,넾5��&�5*r�ѵ�
��ۢsQ%:�W�"��������X䥤#�:�!�	�E�O<BH���h�d�E��*�v^��FyN�J7r����n�t�G1[��%
̬�kf�,S+d�Z ���6������H17C���|	�|�8�j!������ӄ��:l	�l�T`��
+e%���ǈ �H
��T�ʮ9l4��f�Wc��h
���J]�*r�R���a�&OR��R]Vjj��Ђ��>����m` g:����5�km�d'{�S��Kaz��	tO��j"��.XM����;@Q*{tj"��Ɏ��=�Q]��v.����X�h��'F�VΔ��͛1J��M��G���I�1c�HL�1'����ѯ_;t��
];c��.7���킱�za̐��ѡ�+�QQ��NU�ҫ/t�%����c���}пG7��#�ńQ�1}�(L7s���xL���#1g�8�%s�a���X2o:ϝ��s��ߋgK�5K�	�\�`:�-d?S�x�4�X:��MƜ��|�,l]�
��,���3�h�l,�/���ӱp�,]8��/�X�q*�+7q�pL�4�P�f�w��f���93'cŒ�b��-�\I��v��Z2�6d�^�u+cӚ嵿y{�Z�Q҆��)�Y�bd�x��9b�t��Y����h��_8�i�|�9��`��YX�h�-���K�b���X�|&�.�!�Ϛ7���,��}�Ga�w4�X��q ��{$d��)��	�Í��qj�4��±�R�ɮƩ��
��>����Ń�j��(�~�H���q�(w��1�P�r�	�@���A�4q
�1�X�tL�i�h���a�D��E��#�̐��(��5��0&9[aeI�W�ǔ�|,����QX�Ց�(	NGzP:ڗ�@yi���>�`/������@HP|��C�y��̀���_\<SaF��k #K%��}$�-�a�;w&���✊@�bD�W!2����	(��g�\3`m�(![�v�O��el���	'�8x	9y�ٷ�e���OX����"<�3�R�!>�'"�y�����ABV/$��Ctj7Ĥw�����Y���?��#��? �E�Ѧ�H�UD^qwj����j�+���`t+鄹�����5����K�RГ�f8��n�ƑF�k��h[��emQ�U�V�9h�\����0��7V�ưnC0�s��=�����6=�6�
�����8���¨�HDG��<*�a����|x4�"�-�(�Q0��)���Y�x�Z�6�������紮�ͬ�IJ>l2�`Im�Ev��a�V�⮈���#ƢϴI5f�[*4�:|�6-���K�g�t�6��g!k�L��������V66}a��z�]aMחCA%<J��N�]z�Zó�-�
��Z��"�UuEn�!��1 �t�F�tDx�j8�@#"�!�bIX�7��sl;����u�������nV2�V=lP6�C\Z��r�B�g�I>������_>��9��h�E��X�f��ͽ�(��S�f����(��[3*�\\�"*��;!��@���
��X�Mi�����"�D��,�'dC'&�<�U�h"Z�_����sk�����K�ۯ���<�;�.���[���><|�7�ní��q��<ܾ��^�Ň�0�z�'�GB�Qj7�=a��f�0&�6H/�Qj>,c�`O�K�]<ݔd�\3
XR����pHJ�uL<�tBQ��Hl��Y����C��Sv�GLD &DDa��6(�b��.�� �k���r�8�@�~R�����Hka[=U�V�������d�G
V��TI��S�9��i�*�� �n1h��~���G��Qt�B�G�g��AX���	X��ٶ!��M7n���b�$&%�b��B�q��(�,-�����0��d�o:�y�`O�L7�j����a���X�b'����*띔v~̲�'������(q	B�K(Rl����1�_}��0r���5�l�o���"��	��F�o�uc�k���z�N�m%�Gus��ْ�����f�0vA�k8�8����z�����3zSG���Ce���=L�Б���4E��)Zk�"_]���(�k��1�t���0�h=]�����!"-h۔ �@��ʓ��l��h+S$:Y	���S}��k!��At\��b쭑@�H���7�lnL��ᩣwM��׆ͰlH~Hzz���MfjCnVb�w;Yu��y��[����h��y:VVi�v��7@���8L��jƈֶD�I��3Դ��铱x�L>�F���1�`��?���D��*t��$���j���#Ġ��ЭM[���Cv|"J2�P]X�.�mн�=ȱ���eQP��'^�nC�`�VmЭ�:WԠCY%ڕ����;w����0~�`L6�F��xL�܉�1�T,�6��Ϩ�Ϛ�%��͞4�Nn+,���QK�b��%X�h1A�R��`���b��ų�a���Ys	�a���m9��t�<,�9s�MÜ�S1k�̤�̘8Q�ߴz-��� ;m�̝/�]��`m�l^�[W���5k�s��Z�ڸ	��¾-ۅ�n�F~�R|	�� �녿�[�`���t�uB�V���e˰r�lݸ�6�ǎ-��-doƖ����n%����U�S��b�e�T��3f`35j���Á�㱳�vf��΢.��~0Ύ_�=�f`��9�5c֎��5C�P�s1n,X�����9�j�d4����!㱫�@ln�;����j �S��]i? �;���p��$0GM¦�ð��`L�9 cz��t^Rq�h,��*N��I��c
�u���G�1�g`�L���s�`��5X0c=A�6��۩<�o��e{�mA�v̝��f���y�l�V�]X�f7���͘=g���-؈9��c��X�l;6o9��.�ԙ�8|�2v�:��ۏcǎط�<��&��l�z7��5��z�^����\�������V��CWq��
�>Ξ{��`���t��X�v���c'����k8y�9��'���ٛ8w�~�x�.�"�6�_���W��ڕBW/ߧ�w�.^��+W����'���9��{�#�v[6���-�"4k�K.���B~n=z��O_���7x��-?z��/_����xt�>�"�x��7���Gx��	�?y�����;x|��;�ۇ���XP�s��0<c�~(��	�#��o �	���a�X���p.(Ddu
f,���+0emw�WĈ��]:�����v+T�#��!�¶�M��GVdt��#��f�dT���>cQ�kJ�AZ��H��Q5}��m���Chu/8f��*�������N�U��)�C�|~1<rK��>y�����Q��l���$��6㧡�ęHl����:���j`���1�O�B`EP��;%ex��������m��AI[��S�Ⱦ�`�ۿy���~��3��og�努ؠf���>��,��]:�^b,��.]���Q��\�����J��k�@j@\��a���(��P�������#��<�΃i\�x,jF�g�H�q(P���+p�L;ܸ�����{Cp��p����ة!8m���������vŀ���j� *�Ў+�vr%�*ŗ.<tk�VBd�3�\�g��t�Ǧ�6�zgT8�y�*�/G�F�k3nj�NDHi�|����
0	j,}��7',2��Pws�hƒ<�=�T����$��q��
��h���6ΩZ┬n�Zቪv��W�^�fH����ы�x�tT�`�{�fc��T��)X�EP���NZ�/ o�kf$ctp"�DO�*���J,Jn���iXB�2��>&,s�Ⰴz�s3[c^f	���`�s6�Fb�G,vx�c�{468�c��v�W;�`��?:��X��*�[1��C���~��уn�d��T�P�; �%��Q���@������� ��J���x��8W��m|b�8k?�������hʃa^q�#��\#��!#|�0�;C}c1"(	CC�0 0�C1��cd~���oj:GE�:0H�G#;�%�:6%�]���T��
U�ơ2.�S�ѷ8c��`b�ն
�	����F���*����V��-�t�;ap�2�(��W�
�rs�9;=�r�.)��A(�B��$t�����Щ��zyx��R�#�����7
�����@FWw�x��'�w�8��ٕB�=�u�t5��S\6Ɣw�jLg����-طv#��� �k���uX�`C�R�ذ]��zx�!�;v�N��χN�莃ؿy7oۏ�����8��(��9�����ޣ8��8.%��Ҿ�☓{�Ğ8�s�Щ=i�Q\9v�O���GN��S�|�����Ϝ��sq��%���".�:�+�~��y�st��gq��\��2�]���7����x���������3ܥ����č��q��\�tMl׺����?_����p��a_>�p�}�+j��<})�q������#<��X��W���?����<��g/�˫�����Їgo���3<�#i$�>~!������~��\���w��������%޾x���މ���c9^O(,���wq��-\<�3~>zg��8�[��=5�x����������������{�~H�>>��w�����gb����������������'��k
��xJ�O��5�zI�=�c^~�cH�?�Ӌw��7xI�~��9�xO�q�_�닏�����|y�_���(�o9.��W��ͫ���ˉ�B����wʧ"�(�^�ޭ�}�)�_'�~�o����wq��}��G��y�!��K<}�Z@ͫ� V�d��$~_��/����/���Wf�����򼸼���O�t�ZگǱ�������X�u��7�~`���G����y߾�A����ļpP����9�xj������ć���7�p�ӇvRF~�(����.�N���W��M2�-ǍW��R%����Ʉ���y�/��m۱:�-�7iX����S$F�.8��AЌ��{��wzg�zH;��q5��hh�.o�!��"��p$����=��{�:�B*u&���CQ�l�X����(�X��.�PݳJ�T"�*��*�G~�jd�m���D��#�&]�tD��ݐ�.��Qp���)�W��@DeG��=�>�e�l��C��`�(d�����pO)|�O ��66v�i(���F�ή�q)>�-�^�0�l}������U�{UL�D�W�^�[�ߛ�y?ϝ��6⣁���a�_� }��=vtœ�T<����CT^0�ݍ���J�ab���rx��@`��pj]��Rxf��SN[Xf��yZ��-�ʀ�"1Y�3����Atk��w.D�a�>;K��a�9UB��g�����J��W�]���b}9�MCf�Tķi���1bg��#�H��,���(��};��\�e��/��K*ZL= �v'w^j$�� �L��V����7u@c� ������¼��i�cD�U�Y��<x-԰WN�ܵP����8�P�)�P3�|�N ���4Q�9#\�0�U$�kKڗd�%�'b��Y\���1#�f�Wci�n��g(���m�F`K��X�mVu鏕��auׁ�2h����C�a�ةb��=3aפ��4z6N��-S�b5��W��]ԣ>2v���N�1{��sp�43���á3�{�d��3G�ž�#�n�,2�&LƼ�31s�t�6s'����k�6a�_�;Wmƪ�K���_�Uh��5ؼd�.� �z�R����`c7�/ۉ-Kw`���J������z�{��{l��^��7�-�I_�|Ǘl�J�\J���q|�&\X�7wǝCgq��A��ç��`������8��6���8�s�<��'�Q$H9K�r��i�:uQ���K�xv�:�ݻ�_�<������u�ڵ;V,�ٽ{D�����x|�
�_���7�7{����q\=q=��;7���E<�x'�o��y3�f��[��.����Dؿ<N�S����W\�ҭJ5��7$���)�l���� `�t�)^޸�OO^����z�Iw�_�������O����K��_�=��>㷷���w���z�1D��*u:���3�]�m	�������'�Am�o�~�g�˗�T�K�K�n��~?����k6֯\����D�/���ZIߎ�)>}+�𺑬O�1"�;���������ZQ�b�z:��ޓ����l�7�_��0�O|�G�J���~�D�s>�Ò���$�'�뚯�3�����?~�=/�fI��&<i���,N�N�s�|��].M��:�=%�%fi�.N_x�x�+~��쩌X���A|n.'>�˒ H�g]պ��dq���_�U��Β���K��&^'q���<�b��7�ϟ�у;�{� ��]�{��=zt���۸�������.�;���۸{���z��^�z%������t��a�3�c��}��ls$����_���l��F��$�#۟��{�Ļ�$�ڢv[�c�~�?&L
��z!R����#�ˁ|!����Z����^K\q�:�虮>�䜜�
Q�_�H��R*��?�*���ק�pt�t,L��P�sOĢ�4�LHD<u��bx��p(E�C>":q��T"<2Ґܵ
�CR�n�ꌐ���艸�Ð�c8rzE6��Y�!�CW�������C�ؼ;ֆb��@�_\�E��c������R0v~>�*�����1�+ה���V���=~��#g��'3>�m�SZ��|�����+�7h�&�C�шm���5��͇��:�)0NɁqFt�Jԗ��xө^$⳵�0q�]������3�W��6b��Xn��V��E��!��9Xne' o��n;ᓱ~�w�+s�4��C+<�ǹ��س�+�%`Jq�~ PL��a]R���}�w"��áA����>#�h8��U�$�&&��o5�Mj�� �$�!��5��f�U�H��Bu/t��a1|J(z��G���(�����(�Q���j�Ŧ�8!f))�LN�Y\*��a�	��"1���
ޅD��!e�pϠ#���h����Q8|
�[u��W4:���[ Z�zC�����H��C'G[xG4m�_�;u�M^CL�r@^;+a��!95o��c2j�/����猦	�+�ሼ6Ψᒺ1V+�#��\Z��oqkl_��wlžu�q{�<�{/O\��wS/�n@��7���޸!�^Sc��� jh�����+r'0�߿�x���3�у�o�x���Ro8ږ�����W[c���
�����a�B=�_>S��1������4�<c�h�pؤ_ߓ1���Y���|=7C��f7���/�q�\Z?�Tt�otq�2����k]4���'�/�?S�@�)�G��F���@���}ucq#�~�A�	ĩf�㾈en�;�)*O��}d���>s�dI�x� ֗OxE�˫Gwh�� ����<���A),��{��"����X�*W�l�)�q��SS_��+ŕ�����o��|�(foas�J�FAj��L��:��R765���k���|mt���5u�Oi�K=:���nloح����9�����Dߋ�	��+#=?���Y��᳑���8K�P�E�U��Ǉ���,n,��4�6��2�����=Jˌ�"�H7'����G��ׄ���{I>�8����#U<"ņ�+�1�,�����ϔ �@�m�������R�$a�>Q��|�H�K����!�@�t��4q��z���=�-� �{�X���b[�m��ݿ!t��-< ��������w��ܼuw�ݿE���˗O���|��R2�ũ�|�M��_��Ab�S�J�߹���~�-IՉ�Ð�|=�-�?�!	���� �\����눝X_�������;Zo^���]���yxK ��;�gh0��k�~���g�n�>�m�u-�~��'��_)O�L%g��~�����őSXL�M�'�������B�-:�	�p��IT,��B�
��p�&��Ƕ>U�H���e�
]�!��H�w�GVk$�템.C��m,�k�1cq��B�O;�>
�5x��->�*�>{=w��ǝ�=p�YW������ǃ��6�"۞��w9Vl�AX^�
j�WV��"x��Bh�6H����!�c'�d��̦�E0�́I|��2ī`)���a�<x �g���o<�㭩>��᭮>9�7;<���:%lճ|��І o�?�i]�/!����sf`��#���a��2�i�㹙>�8�H<S3ǯf޸I�w:�7z����
�[X�^�㉶c�B�����p��)}F"�� �U���h��N�N��Z��$D�xb�6�|������#��O��ݵ'b�J������~�Q0� ��SW����h5�Z�S�)Ca���x��&NiY��)�On+T#����[�*5�
"QJf��(<�z߾��ZC�;�(�yY7��P�z�!,��c�������U���jc��6+�Ⰶv�0�>eK�U��^��N���)�a{KClQ��lW1�^EC���#ekT�AT��q�¶5��km�|�^?���n0�1鮡��JX:�!�d_�qo�J�������๒d��
�mѰ�;W���ew�� ����]74���m6�F�*c���s]I������W�$i�T��{����^�|��Hu*Zj������G]q:�n�)�<%i�ƕ+��~%i�Pȟ������y&�x«�p%.����|I�O�Xs#��#���<��9�Jz�o������J�\ş$7���c��}I�!�Ci����Su�����'��t��D A3C��
�y?7PR�R�޷������K}�?�����:�H����������׿F�$F��a,a��e]��o�]�u�.	���u�ʆ�X7�uߏ�߾�����u���zx_���Hl��<jG�ѻI���x���{x��� =�7�Խ��(Z����|�G����c������|�������_[�0K;L߈�n12���G�o^��uO���6?��N)���8I�@� �(pI�%�5��e��I�|{�V�t�^�����93l2v��X,I�F��8d�%�y���R��q
�Qb9U��p��H�d����q�e=�w�Wa>��v@dE;�w���b��g����=��s�@<��oo��_���/��c5>|����x��/^���C��]_��ОTF)���+E(���$t邰�v,�@L�N���cV��=�;��4��eB.>	��Ʌ�bu�UK��֦}x�}���b`"^d��SM'�t���>S&����#KW�Q��w@�ˍlpc�
�d�p���`�6��;s<ݱT[�TpR_�m����N���\ߚ@OGlq8�W�f����X��"ӡ���PJʁun�KVU�V�����h3|�:�E`F22*|1oMn=�����(n��0�E� ���s��]���r$�m��6ň�*@lu92�vCLe[xf�9%~E%b��5� ^�����B�/��;=^ْCR�D٘���?�]z���\̻����.a������OOo��c��?��:ᰁ-v���Rs�����xlu�節���n�xls���8\�(��llu���I���L�H��h�Ա�my앷FLc5�䗀ײ|��1�`�.��KpC��],��~�(P�Kŕ&�հx��Wz�s]��0��Zw�:~?����㤪�`)>���̽5ֻ���{�&�=U�(@���W��>�� J��$���x��_H�,B-r�k}{��b?��H���Q#%��$���bc[ �  IZX�,������ⰿ͏�y�I��%/I�G!^��k�?�����$���$�?r��9�J��m��Wm��C}��JLn�M�~�T�.����ו�ppg���sP�DrDK�M��1߆-��+����?��)U�u'��\⚨��G�[�?QZ���+�(O�h�� P{}P�OH��ƒF�� �_�٠��W Ozz���u�S�Di|��jENl�Q�ӧ�ǲ�$�J0G�w���������k�߿/t����cȓ����!^�R����?Ɵ��C���O�%.�<�$���~�z��8)���x���|y���A�w�r��~���v�n�h�������8�f�#f^���9�^����,�%�A72���M��Q2/��� ��!�g�� m`_�X8%#GÇ@/���'�`Ғj,XS�U[K��`��-�Y8|.�:�)>�(yx�1�~.�Ɲ��8sV�`��b�zڙ���}�e�:�rL�z��oI{�&��.%��yЏN�ZD24�ҡCa��!�K(������!ql�^&h?G-�q"�غؾg�2���������W��$�3�~c,3����K��$߿7��Mwv�2u�TS�5#|�w�'S�շ%�㾒.^h�㽑�;ࡑ%��j�\����V�=+�1��z�!����D8�&��6�g`�ꍨ?U#:`��|l=����J�uO:�tDJ�3�b�������������"�����Im��J���G^�X��g�v�O�c�a�,֊Kh��ݺ�g�c'�p�h�WÌ�k�E��{�#)��h� S� dEa�a��'��☦9�)ia��6��҄�x<en�[��������^�sc�R�)x4v)�,\��K����u�8vn�����W���X���ʎ�*g�lU+L1��>�����'��o(�c�l��wi��6�_oz~��I_q3�5P����C*i�/U�_�Q��_~}'�}��|����x�I�(�%���J��J+)�89^R��>~�������J�ح6>Ti���HG�~$����_Hz���C�U�����7�%����T�H����,i�}/��}\���?�I������?��!Jd�����#i���<���?��s֕0|n�?j��v���+�Q�I]z��zJ�#]uEA�o��c��W�y�SW�*��r��O]���(�#q����;iX�pY|�:�&����j��5�����x~��(D稻�{(�*� y�)��������K�$��u�6n?���o	[��}�:#y���~���i�?�ݻd$��z?J����"��.ѷe�������>i�|�#�O����_+������מ�%�g|�1���ګ�v-���Cȓ��q��[���'�P={�p\���pT�
G�m�[�[Ll�50s��-5ᩉ0O��VD��`��
��(Q��< -�#�Q���& e�P��#�k��?�����c0zF_�Z�aS;���|t��{�S'Q
:���
�Y���� tX�a3{a�A8u}<%�7��K�۠��8g��4�FQ90�ɑ���
��\���#��y5�1p0Nlށ݋c��I���P`�R��)����58y,Y�����lB�n��x㱵����:&ثj�%���(.\cH��{��I/i�KnL��Eyc�̱HV	{TTq����m�^�/	p���X⹆	ިXዚ3��wz�8gl��!A�ֶ=�V�A^�
�d�41��h!��k��88`��o���}�nl母��k�t�ebϾ`l�]��[�`��6����ga¤<L����S�1tl%2������"xe�
J�_׼r1׎Sz>��uDɈ��0���O���r�o�� ������P*��T$R�u�L�8�0��t�N%=��Q�EC�P���\ܛ����°,l�n��Fa�)�1g6N^����`bV[��3O�ěM���Ug�L��^�po�v�쀓Z����ź�X4uQ�g/����B���?.��ߺ�?i���.��ެ��'����ʖ��p�V�R����>6�ǋ�ppl�oI�a�Wę���rI�Ϊ����*ٵ#c���w����<
)}+�~��(ά�J�;I�KU�Ȑ�i�������x�祖��2��Y�8�᫾��H#��&q�����q7�_-�}/�ܿR�t}�����_�u�wE����|U��`��O]��u$��y[Z6��G��@��^'����kYIU{��J��G��~�J���1}I�?�rdI�V��ڴ׭�	%qYr~|����ᱤ�=��cI�_z��e)�����uF*������ç�p��}��{��zx7��?B�D��/!�$�/�?B��RГt���<��M_�X�?�\���w~�,�o��Zѵ�q���ȓ'�SP���ZLi�P*���o�*��?�<<�{����tQr�iM{�T3�QEc���a#2��&kg,%f���2���d�e�)9&�P	�(k$�A>4�Q	b�|��x�B��A�2m�nۄ)+Vc%�|�F-]�Ҟ�X������x��#�n��N��4�,C�ðh�0�yՏ�u��k�H�QCK�E�C/� �t��l�'�ÿ�J�����=1�m��1��ħ�g�3��j �y��W�t�O�O����=y1��W_�� ����ݱ^�!��Ԍ�����%W�=�#��'.�Z:�F�]|~��S&`��;6*�a��.I�b�B��_t�N�����R���,�F��,�^�/u�q�"��#�+q��+����m;!���I	P��BC�`�s�C=GW���\x2�1p�����{!�y;��&��������K­k>x�2�n�jTu1CX�J{�ANϞ�IN�gI+d���ѡB�tBd�p+��]��QP
��v���vh0�c�����"1I���dl��1}'�V5���*8�HN|X��(�B���3bfم`��%N+�Cvd`m���<a)&U�Ǌ�^�\��}q+��8bB@2�MZ�_�m���\Pp�Φ��װĖ��D�/n,�������������Խ��=�B�n�%��X|Ëp�N�c��Տޫ�=������9����q�ؖ�������c�J�n����l((� K��W��ԕ�����n��U��M�/~Ć����x����"`�$m(���z����M����I��ۼd�?*�x�{I���n��nҲ���ç���AS7��K�%���m�����g������/�C#-��?g$w����s�����G�[��ѣG�Ǳ��	�6)ˏv�����}Px��Mz��?@�����K~tK������=#�1��/ʚ�1i��p��3�<w����׵�a�㎢��bH��Q*ş�<�h�l�$�&N�?�~é�ӱ�.	'U�qZǂ�N��qTN����U37p�E�h�Ĭ�tt��F|^&��2`����8%d��S��֊L�QR.s��UZ��N]�ճ7Z��c&�d�xd�o�Ac[�����K�}�Â�%�l��N��f�x�+�mv������lz.�~�d�c�����*1rWա����p'����p4�X�_�� ���]�ؕQ�?vţGqc�~<^�ǲk�������ZO�p��U�Z�[c���=��%}�<Qx����_^���)Xh�u�]^���):e��<-+y�4L	��� 荺%^�ZṒ9^�[���)�:�]0���`sq%�VT�kI��������A}� �s��f�'��5ękA8t�k7�c�No치���Sp�)��R����?���<�y]�~����sQ5b
���/e�sA1��J`E���ʍ�࣒�Y�p���DB/$��IMDvj:%$cTpV�a���(�ᢌ6.�iᔌ27V�y,��ŭ��q��4,��=+\��'��a�]8���������x=q5vX�a��+6���Hr!ތ]�����hV5V�8⪲=v+٠��n�Me�K���w�_����=d0�IGۤ ��y�\,�oI��ORH ��w��aJ�F�.���D�I^�'��K�GZX�l��^���BKTҔ�_>KFx��b���/x����<Uz_��+�}y$i>��P:T�o��G�|o��7�{�+q�q���ݹ��^9���f������OMݲ�����W�g��������|��P*��A�������{�N�u ������<������:�X7ܿ��z����L���� �wF�f�{��w���~p=�!�����Y8蜉�8�e����8�n��j8�b��Ƹ��W��ၼ+Ϊ�8bA[ϚR�m����H,�DH^+8%�4i	ЋM�V|4ⳠM𧛐!��3�ȂEF,R�a�]c^�<{�t'�,���i3?�!PK�Qz�C��~Ӳ��X%VLŐy�H��FfMZWv@��}�x�R�7k����%��s� � {�����}�qr�O���ʁ��K��k��m?�oهWG.������U���x�ۨ���چ�q�jS�����!�Q�_�����o�u�u�]Ե��<1�ǐG����=�4�5<ױ�cs�S6�ݖ�x�l�g�&x�e���x��+Aq8���5��_�H�τof:�`��zXv<�f�!�@�HNS[���\t����1vq!���A�ɹj��<�綇an+h$eA#*����BK�Hh�%�.�f���xx&%#9+չy����)����8�b��
&8�LG��R�B��tp��+Xc��7t�s��af@�ia=l�1�2�0��1O�m���q1��EbUzVt��c��XQ{,7��b}{���9-{�R1G��N�:"ni��#���{mu+���!�P��7���_A���p��Ň�J��Ҋ��*�Q7��"'������ٝ%�S �����#j|���?�C|��HÑ�_A��#�������<�ۏ���_H<bG�Y_��ǸR���Vn_�pzň&���K�ػ�x�����.�ے|���$�߿'���yB�����j���+I�����e���~���/�~Yߋ!�a��۷����|�:�� �B����Q]��We��g�\e��3�i�}y���	y�J�1��SÇPwz�B���	-_�4$�S�Y^FU�
'T��ݔ'�hi��n���QX����(�
EuR����i��X�����"���C5%-c��<*Z�Et�b ���0��aвV�}=k���rX<��B����腧�&%i3�uF>&�)��I�գ;�����8��o�����فð %/�,�U^Yg�p\ްw7��.X\��q
8|��,��������xs�%�/؈��e�l�_m���޻�v�a���.�ɐ��~P�l�������;�͝�^N�Tp����Q��Ⳟ�C�^�≖k㱖	j�ᮦ��y�T2�o�6x�`�'�f�F xH�����?3�0,5	�s�:� �E��9�+�$b�Ld�z�(�FQ�0��n�="ma���G�ZC=�
a��K�LP2Z��A9.j��bB���F�0$nD��Yň�*BVq)�33��2o���[4t�M=�nj�3M�p��6����=�3�99+\Vu�5'�����s��]gl�u�'o�o����c[�8�{{�`��fS����}�w�"/Y���X��9�x�_�ڶ�K����;��������]�}��3�������X:)���_A޻� e@���O��x�ߟ���ľ���!�߭a����8�@�.d�<�=~��?�`�b��f��0V]���<�D��4й�xN���~'��o>���$���y�g�E�i�4����
H�F�x���������߄x[Ȝ�q��]���_ȫ����w����������W�W�Gq���m���G�ޤ���31��}��GyZ7���ǆ�֤���s�HR������3u�2>�T�i��n��<��VA� O� �����쌥8P"��;�n��J�8E��O�Ψ�㴲)n��ᑅ?.;��[�9���>2�4���MD���,9Y,��gX?�3�Cـ�������!�U�Z�­�NEEp�/�cn&�b�&�=-Q��1�.)@|Mg$UvGveW�w�!V��7�
���aIn�&g�O<���u�Fg3���'�����x%��
\~H x�f�ǧ���׵w��c�}N�w������.#q�1_��������e��=�,XB7�ײ�����'-�/������m��j�dl������t��F�/u��T�O�%��H��[����TȖ7#{�mpA�g��qL�������p��;���#*��3�$=;�����ٍeز��&�F��ȩ	CV�`�T{·�V	V�Mw�m�'�"�Jo��$
ν8n�yp�JF@qb��UX��8d�E#�/�.^Ȱ�G��	�t����%����3p�	yc�V0��اb��g[X�rK'{����k�������qn�h���;O����ql��/�9��qx�4�9p֟Ğ1+pj�&��u��ce�����71BG��?xV��w]���˚op)�I��OI���� �G���ӏ��XK*ɾ�2���8Mw4w:��Ͱǐ����H+��R�<�m�Ö��}��7�G����I�=E����%>�6��n�%���y�y%F�8_��ݯ�B�� O �����ޓg1=��c$aH���H��;��p���^��q��n8�"�u ������S�0��������.�ԏ��;u��6�C��H�����:�a�����c ��������s��i���H���`�;Ȼ�J���ǐǟ��ǐ��7���
pR��lpV� ��q��1n�]�q�5� 1��GOt�5F��*�dU���|�u���6	)��k N�܄�[���-�8g)~�>&Mæ	�0{�0���}{�D�>�1d� >�F���ֽ;z�퇢ΝѪGTVנkY&u샱�ۡoN&Ʀ��Xv���e^i�⭎j;�(A��H��~ �d^���IPk�f,0f50|!0u%�|�{,�y��I��@y?������'�`��X�
��Di�f`&V[�o-�'�
y|K����#��`��V��`��.Z㣹~5p����:&yxN��b�{J��X�Ռ��O4-p�t]�
gTMp��濫���b3\�5�!���6�o�}v�8�3���g`<֏���q�6�5f�-Ì)�1��&V�����#g���9C0ht���}@��C0dꤑ�9k2͜�YC�kFM��!#��2�n����HTVE��:R����v��Xi�}�Δv�U��qe3S0ũ8�����gm�K���}�b�b�:[�˰�;�'����qi�\1�/��΃�, +��pf�L<X��:��K\�����6h��S�N�{G�h�H��Hob��7|k[����?�<�c�-�R#�_���~}W�?��FߥG
a�M������2�>�%w��}��7�R#m����~�?�`��G�,�w����go���'^u����B����	}M�HI�J�y���o).��FeГ�-A�}`�_��ƕS"ͧ�#�
��ϐW7ϸ�y�X\�u����?5?
������F:�'�AU]����l�n�'F�.��=~T��HG��L����.�wFZ/��?y|խ��-�a�<�Q����UpU���㺖��%�TH2f�Uj�#FV�M�!@^Ѧ�Q��.ǽ�;�j�A<#��;e5����]q���WauI��Ɣ�
L�n�)�;cy�AX5h$�O��c�7������:֯؁%fw�l7o�:���;*���E���"q�+�K �]�A�oupS��)��=q�����⥒^D�}"���O,n���O���&^x�i�'Z��d���A����t� <��������[���e��B��1�^�+�9s-�Z�N�FtmB���@�����⍮)Q�^i�㕦!�h��R5�#<V6�q�Y⮁�X���>e�;FrP�@h_-�lA�l�'&x��S��bg�..���.>�h�n�^�٣͚���W���Ux�k�oX��+����e�>on.Z�{�����x�r#�ۂ�k����XХ���0,���m��� ��*R�t�����fj(S��0-s2r�m=O�P�/���3�)YJK3�_eK�Ұ�!;����fn8�l��jָ蛎+���蟉���8�������X��\p��	Ǭ���C��]=W,W�Fk���w� TW��p�RW�v�s��I���I���a��U�"�/��*(�|��1p]qc[W�C����I;��<H+���4,o�ȓn�m���?m�R��<���?y�����K@�G����$�'�;rg�8(�7��kʃ��-�~����'�+�4-G"=�?�<�u%�<�����3���Ga��l�x���?n�5��|��៎��;���t���YS�*�^?�N���W ��>7x.����r �k��q�=E{��p�9�PI�['d�+#]N�2�xV�~AX3v"�n؆[����8�uv�ü�LLr��@�5�Ew���hgj��6.���n��ᕈ	~)X����5�qw�L����6����������C`���&� �)�4C��!&�8�O<��㥮�X��C	�ֶ�UK|�v�k;�Q��~0v�sG��ì��R���Lɿ���7��\��u$s����'6�)Tv[�� ���y<b�৏/qh�$�*��{oյ��Z��e����]��Zh�@�B����K�Nq�@�$H<��@p��@!.��ONR�������~嶺393s�ڶ�o�m��8⺇J\�����y�y�� �PeO`�G��^���Y: ׂ �\M��G��W	eȋ3�!�L�hW��uG���(|�kW�ܛ#�w��7����TU�Mu�1�B[,��`i�^G&�4�mڈks��܈���a�c�w}��� ���;v�;����F���e��� ��?��A��]�~��ϿAO�>y_��1�'�����fJ��Pb��ι6����K�Ǜ�!�D���Bk�p�=s\5��P.WU �"������0���{��L�ˬ�B�{U�^5�����߷�\���=�?Ʃ�/!O��
��]���k(�߁�'�]Y��7A��!(*-�>y^*^�;<�[\��b��K���P�x�{2�lV!�|�3����F�M���z~�.�c1�7ɲ���dO{���<ƃ�2�R�d�c�3��U�N"C�!��R���/�<�X����/C���f����N��	�F�%�,���2�y-��\��2!_����{�T>�*���Y\v���`�6/˟	xr�{ʠ�:E��p��?*��7��ۆ�8䱡|��36"ޣRm>m�U�m]��}�3-�a�_}t02C[K�[i�^�ٝ{!io
��A 2t<�4�[���j�1Q���l��`#j�kؠOk�3Qc���Zhѳ�-FR�<���5���ǆz���ŧ<ώE٥ȏ��mæ�3�ʷ5T�tƷ&��of�����A�,�k�lKw<$��7���3��܄ë�^�l�o�#���B�XiPh�L���Љ��	-]���E��J�k~��f�A�J�9z��c���X����o Oe���g����W5��,���ষ/�U�y
�]����[�Q;�3�%ǚ&8�2U�͒ӕ.��p�������������B��+n���5��8J 9G�G�*5Ы�	��f"&U~?b8b��D�)J�����H9�m�b�G,v��t�FZk����Ml��'[�1\�	N��޿5�|3�G�B�͸"�����`z�o�)%>{���P��k7+��L�Lq>���t�q�H����	��	�����-�p�څ��!�k�F�5�\Z�l�(#-�k��P]�ՔH6�!� ��_L��,�-ݰ����?���xX�'KE��P\�^��g����k(\z<ԕ=)���Z��8F��Xo=RX�T�����x�^�^�b��ׅʞJ�h�"�,N3���sE#�++�Uz&���PM�	K����7/������>��CVA�y�r�sd=,BN^��A��.��,6	 %a �# Υ7ČB���He �4���q��t�%1��VZ����d����"Ý,��P9?*����iUx��L��������?X7^��m\Xx��?��{sI2�*���>���ρ�@Ԅ���l�U}�b���I�uq�vc���Eo[[t6���5-�m�ص�'<:��cѸ��F��f�5�(�3�9�a��z�4����m�1̲\�K�t�7ՠ��C��N?b��5�1��%�P-�-�Cږ=z�l�qp�/�qCW�ő:G�U�7�f��7�Zt@�[3ܷpDf��
��J����1#��
 K��e�n(��D��J5>(�#��%�s�O��F���m<������0L�߄W �3K�8C�{^���u��Ó�MS�p�ӝ �A�+�m5(�s��q#�sF����P�e�e�=$���ظ�}�w�fa�c��Uz=O�s����� ث����m�,�]�ǲN=������;����?`���K͝�C;̬��c5F��b��z��� r��%�� ����5��kd��Vn����[|��_tî�3qa�^��!?.ň�-��5���F���
�mm����#̅
#%|��=��;�
�$-�M4b�7�{���E"=��!���a}7Ɣ^�u�l���m��9�S#����]�ǯN�20p�H�� � �*���J �gy����c�����\ѹI^<i^7��ַ� )7�T��<�M�mrCl(�
���"-YXO�L�iƯ,�wA�p��<=�>%��`��1=�yeb.�[���1�<��,�T>�-����t_~e�3�<yh��H��<kx,�!�0-Y8���=T��w���C���,�\ֹ�+j_P,���:0�ɫnSS_��[Yxh7??_�������T��lO�n�w ����C�o;\��"�s��Zp�~S���j%Z��o���)f��a��ڑ�x�/'M�چ_a����
g�����Mo��
s���b��� �#�f�z!���o�(0��r��ì�n��P#s�i�����ő)3Pv������Wb����(��la��t�`�z����uŮ#�ʹ(T�	�3�<�{���J�w/�D�I�^x��;���)�<� �K���Z{
��k_��o�[!�"�T�Jr�v%�����h�p�� Ν �%{��<'< a��W��,J��V���K��ID��Z/\�n�C������Q�=%���.��g0������A��k4�Q�皩1�L�!a�?0����3�q+�)T議EO�>
������ݎ2S���Tj(г���Ё@�C���賎8��j�>�S��bV�^��@�E#���ŷJ5�57n��H�z�:A�-�F�]2Ӌ�ü7����θh​�t�?#I0�!�L'��y^"���ැ�׷ΆEI[sP>��0�#^TÐ�ޯ?;01�1��խ�[�Ȑ'7�\�XO~/�1�	��xȖ=w,��z�*߃�:yW��N�h�"�3}����߳ࣿ�wr����x�-/���M
Ks�x~C��	�+�I�K�{)�Y�
��(rPڰ0��pb�}�m�'�-K��0LK��P�����˫,��P9?*��J�'y.^ea/��~8�e`�d�LIIy����g�y�/I���v�����/��>s)"�A�����
�}K<н�)�Y���5���qz�n<=w�Y�=F�g�&c�ll'`��1q�J���6B)�F�7R��pb�A
5������`��I��3�h1��������C�5�@_���I�)��%�0��]��`�����I�������(Qy#��O���l$O�,�哅٩2�<Vz�)�\���&x���)n'��8m��:_i3d�ė��o�!���9y�K!z���;�t�I���;H���s�d�+���ɀ'CK���D�W-��HȀw�^e�K#r���ѵ����+���]\�S�AH�JB��sx�h�?�;����3�������,g"g� [RF�O ��5z�X�W�`�\�v�jg�%�N����@��n�=c� q�\
8��s棛�ZV1�7T(���EGsS,�8 ܹ.Q�ܴ���q���Y:✉I5�p���M�Ď�I�]IeȻ`�ȿ[!��&�<\�!^���g�*�Xc���<�[�F���E��D=� ���A�>ٻ�������=�����m,�^��:�F���+T��h�"�?K�H�5����qr��ţ��(Ȑg���ow�[�� M���%(��1��g
�C���U
��c`�),Cv^�x-���mT�;2�IFV��+�GߓE֗�!�rz�W^���r�����
���վn��'�`�o֑��+�VY��޼ח��We�u�?yt�'��pj�����)�M���J7�n�n��~E���F����␸�Wlo�	?8��t[7�6{��C���̕���b�REl@ ���{�X+1��`�����;��3��B�'}_�1v:�Ҩ0��o����B��uEn�y��C��[�~Jw�$HT����	fѽ��n�"��(���3���<y��uõŶz6�R�y6@�OQ�qL�0sW��ג��=��CJ�߄�@g��8�=BĪ�8X�%N�y#T�L��xQ��E��E$�(O.��xb����i6��F��D�y��K{74��^�.�XL�6�R����@�[>p8
�〤��[�s�:`=��_u#���p���:��C�	ެ$�t��g���Z
��k�Bo[�2U`���B��gT(�J����}4�����z72#b�s�|t�sG˿�-��;*,\V����6�cᄫ�yoI5��bBq��ĹjJ�V��k�3����sF$5���W��>�յ��p�D� �q� �!�����E+�7�����ϕ`GZ�!�����N���{����ǿc�{�s�����5CyW�g���}������H �<dp�k���q^	�c�����<g�C���G|<��9������8�>��H�� <C����������C�����P�<�O�e}*��� �i���Hً��u�7�DY���(ǁ�m��^_�*_���s���{�������8�>_�ȳN��1�X��&*� ��sC��.�K�c�'=�ڹ	��B8m�{7���̨�v|����F��a���:a��;�;{a��7&9���rö<���7\E��:`��ޫ��Qc�ZE�g��fZ����; O�� Rbc��f�.���!��Xc��7R�~�|��k7�8wro��W���=V���g=��/m�B�!^bO^��>O�y⯒|D�^����pR�0{7\r��s�z���ZR��KLdГίu�Cg!ʅ!�-Ͻc�ss�.X:�*E�O�8�Ul5/�Z)c(��MAa�y��E��_��!VSB�|�ݍMѝ2��l����dC�jn+ ��ɇ��(����4�"���ך@�^ywAho3t��Fo�f|�G���Š`��7װ��U,�]��0����|pN���F��#��O���RMkh�@��CyN/8�-dx�e���).�PH�g���|Ji~��F��+��dXa�a`��svx�B�4���~*�;�ߢ�������]�]���p�4c�Y8�� 6��7����g�ڤ�����'e�/+��s��Iì�)-8����ϨN�+��~�߲ȋ1������'b���Š2��q���:3,
��� ��O�e}*����C�v���?_�8�NG9���^_�*_��B�;�~�����U�+R�c��FZ���\���M\�g(
". e�A���V:��LS�%�b\]��1��3�� j�͕n��TG/���Ǭ�0�n#̠���a�O!=�`��&8���y�	�F*y�A��c�z��h��8�s��ۺ���=����}�qױ죎L��s'�%��lj�#�x��D�%̐W�^=�&C)S����ٳ'���B��{������q!�֯�vZ������� ��PJT���%jwz<��cιJ�l�Fp'�C �>�2o�B��g�]�v�M[\u��*;,$�a�B����z �T$�xa���h�O���-�ִ�s&)�1њ2�B��&����Yx�v�� ��?�uzf?�M['����BObG�)=��)���}�p�^A/k��EtR�bJ�b������Wh�:�}���XXo^��wl}��'a�] �L6��%#[{�/dO�y���b�6��9�(�7�����}�'pl� y�YR%�����Nd�yb��;�'�ʋ,��!O>ە������]�]�e��g�.B�ǃA��ԑ��Heah�y|��~�Xx�x>C�<���{��
[Ơ��c�g�"�=��Ɠ�_YJ�>��R��{9]8�|�����o�Ѓ��^�%��i�Oe�1��>���6�c��mS8�8����:o_�*��s+���Aô�w��^_�*_��B�{�8?i�7�E�A�E�|ss1�}�O-��=���p���`�m<0��c�wZ�w�� ��׊��=0����6����х>����.�����^���������a����=0���Վok��t�	�:�!V�D��G�M#6]M����Ů(z��0޵&��c��'�[b6���z�S#�:w�)\��.SH���:)f!����O���x2��iP���<'�C�B�>)D����Z��5&Z���x6�눕#<߮X�!@O�͠W�r�]c�&�SU�]�r�k�E�������O
L�hџ@gj�6�޹%�.#j�<lj�1~��aR531�n�����1��c,5bhv������ҫ�:���х౛��)�zk��_GmÐ�>�x9��{��a�@7%���o���]�{(�;��e��_[߾���&�g�.�˺:wٌ�QQ"�zI�J$�q�W�ԉ�Rd�㕸b5.Ņf�U�[�ܱ������AО@E/!OZ� U����.d��2���ːWq�\��������:�ެ?�.��<f����* ���Iz	o��!�ŕ�B�հ�ť�Xd��!X�"C�Otw�%�*`�$��r9`]8��E���!�2���!T.O��������,�#�)!oo���'��d��)i���� �*Ky��җ�C4��U<�ƫqe{R�N�˥\�?��|�W�T��K�#�UR@@w7���� �$�������}���;��37E{����3�o t���Ӗ@�Sl�3�kl��7N���N�w�$�Z�U�1&��p��^.^�ѱ3VM���5k�� l�f��>�:w��:�0��c�kc��goL�ѽ�Y&�� ~��u�n�9ظax%}�-��.��ڮ#0���͈/�#~Pg5��wh$<yO^��rГ!� �^y�m�w�s��I+7첯�y�����+�'g�����铲��'70R��N��Z�h* �����L���ٓ�����l������沵#��C=�%(\E	2���衰D}��+�^���u[p��wXNߙfn��&J�Pb��[�
�`s��8�ױzW�s��x�:��ꊎv:t!��N￳w�^��'Th;+�0H팉v^D���
*0�F�y~���ڈ��=�]���nu�y�l�8�=#f���=�TS`��=2i�9X�kO�%��I��Y:�6A߭���Z���b����q��^u[���W�(�jj�K�Ո����l勯m�ؽk�=#j*�C�R>��Ѫ,4�
�DAN���C��4��ea�c//d`P��=�ݚ�>�]�gث�-�����F�U��G����N1�*`J��t��bh�~ëcʤU�,��W�ᫌ��=���4GN;�* �҄��\[zeo ��P�XD<HX�(�|n���X$�{�;NR���?�m�����P��A�/\�^'��`X&��)��知ߛ /=��)/W���
�BuEv�#����Ұ����J~~!2�g�n�=��g�"w�fR\��$=�BW�b��5a��~r��"��W_��l��H�L\o����q�{k�l��K��c��w�Y�C���fu�Q	(M��o�c��'�֐�C���LL1D�-U���� ��j���$=]�0�{_D�½۷�G���
R�RxJ�G�Y�J���;�`鈱�E����c<�0����v����F�L�s�hk-&��b���84r&p�w�Dc�ok�6|�V�!ժ�WGܪ�J�ੵ3��Z��y
Г�m������~y�ji����P�r�c��{4�8l�-���;���	��t��� A^ԆU���@Jt����⑭y�D�D�o��ZW���p� ���K%�K!�;H
Ϸ�"2���j5��̃q(=��Fc��/�b���7�f'�z��Bl��s�xU�8��{S��'\�C�4��_a������,l�~&�̙���FaF�.���/���j�F?Ki��p�3zԴ 9�~�R���j�����Z����ؖ�pb�\X�������L��ܮ
5�[�`Qx���*=��&�\P� ��)�������	����F�k}Ĺ��5��X�n�(S7ܵ���Z�`c��;%ȓ!C�<8��z��� ����޼'uD7|�?Ý��?�[�	�(������!У^���$�eFg~d�G���gy�ɶX|���TH7�^�w�Õy����'��� O�����7�"?�B��챓!O�;Y���^������3N�zg(��`X&���V�u�w��6Ȼ��@x��_ac8��_)�,��:UJ ���P�z7�B�	�X��}򄮲����!����{k`Р6�����[̲n�.5�Mu��ޟ��ir�g���ޟ�E��L�R�l���J-�;�a�wmL!H�ѵ!��#|�.<{����B����\��,��!��P)dݸ���[-|��Ǵ&M1��cUZ{#Ҽ�Q����cq���Xܼ=��]Ǔ�L��3A�F���p#�5��i�Q�� �m]_�<i%�K�c~�A�!O��ǐ���5�vCP\w۹ ��q�����ǙWQ+��B��	�ۼ���^�'4��ZK�<}]�m�c�w9����Q�=[\�mT��ؒ$;_laW(�A5�1���~Y�gӑ�b'v7�s���X�m��\�*���*��z��x`��?6��=���/&w脐͛�q#9�id [,"����?D����:!�5i��FV��7?tt/�ִA��Vb(�����l���CK|mろ#f���0�5}){�w�a^���VZs���3n���o���q]�!z��D�5kR��+3�#�8	\�a�S�}����6E�Ez��������o�CO�\��&4�F���Y�
1O�<>�B>т!�?7�U���Z��I��Q2�1�r'���C����"�I�o��R�CC�yyE��������r#^n��yw��<�O��K��Yĳ��?=�C�&���:��(����B�R�?l�Y�t=e=��J�ɰ�������Zޖ�2��\��_Y�����T�#��R� #=�)����{���R��܁C�������aΰH��Un���p�u�5#�3��!�B��=�gL�����}�wSi����!��9l����z�U�p�"���a�������S���;G'k��Nŋ�bJK��/�"���I"k�6�CIvv�X�6�������6�pG��x��8`���,u�`����c���~\Mqx��+wa����O�4����z!׳	��<��ór� <^`�õb�Z:�B�|A�īk��=���e���GF`ːw��	�������Q,�PD�
yRG�I!b����c��!=�	O^s@WEyO�^�<i�gI��^~���6��0yWl����2�c̬���Z�Cj�9<:��NC�M퇙\-�D�v�ȑ��Vc��h��qgLwo������s��]AJ|��`κ2j"S1,�y�xD�W�\:n�ݵWc� -�߸z�uu3���$�tC�t����bC�
+��V�K#�4l��mpf��#�^�m��DO[�R�۬u�Eg\6�ŵjv���q!/*��O�쒵� Q�W"�p,.m8�=_����sP�����DMs'����`�p�,�O'AU1a(��?dcSY����!�Q^	��*@�
��0
C�#�C�Yx��_c�P��Ya�?�H�5�w2�=�/��<���{��z&@������d�{>ONK���s�7O�[�������id(��@y$D�0*#��?�?]OY�� ?�˳\�_^�t�V�������A^FZ������[寕��,F``���E:A]z�m���$���}��'� �8����Üa�B��Im?�rJ/�L	��	������8'��.�x��0E�
���`^���8y�˷���1��3����*Z^�8Xm'�K��q�dG?|�G��n����[�Ь����x�÷8��3a�	�X�'E�i�T|��Ξ���+��k��7�B���L1�clU��b�E��� /$�=�c�-1����ⶣ?�����2k'	�l����E�g�Pgx����y/��P�Z��u�G��h��:\޶�"D�yCy�I������Eo[���`��
�j�4����!��ej/�����![<��B�)�!���`��kq����7W��q�i5����:b˨�(�|I�7�h��X_���%�Z�
ZƩ0Qm����Z��i���˹6��j��=�(�/��8ȍ(��WF
��xI�4�Y����+��)��Ճ��'��x�M���Z���=���M㍕#���C�i�l��7f�ֈ�6~P�#���(MxX����w��G�!{�.�n�Gju@��}�<|!�����>��˱Æ��IS?1r� ��#�DK.o8,��FQ��<����M�5���]"��v�~#C��0�|�+{����
 ���z��%=������ߒ��^�{D��e!\��s&~��$�;�c(����{��� ]YFY�,�+���p��G��x����^�:�n(�Y�!�2c(���	���W�K�"ɫw�=w��9�o��vxRJ�5F���FJ�e�T������,�-��Wi�K�=���r���ߡW���������b�7ڬS��T�eύ���ϿC�7�/���{/)wo�\Gj�-�;HIO���R{%��W�L���B�|�/�~�"nl$��2��R��RF�{����� ժ�&��<Q��!���v���t���((���`�W4��gJ;l�=e�qt�\����$#{���������=0�xc��=z�qv�.�!�7O)]���xQ%��v�VʟO�T{Q�>���71�Wo|\�3}��U����v<��Db��:L5�`hMLh��Q	��4,��;�Y9`L+�n�&ѡJ����g%�2E��	����T��O�*N�`�t�x�Y� ��+��ũn��nȓ	�"7���V-�Qㄝ�����- ��
�<��v"{���B��Jy�-C�q[��v�;btU1ﭷ_}�-[�'��>�]���}s����������c��#-���]�|���/Ʒ�
�"Ρ�P�휽2rc(
-g&U�ʠ'Þ�g��Ƕl�g|�cV��yzߙZ�c��Eߋ2���#F}�!�7��� Lk�	��i�����<й✊���g-�q�Ml=��3� �Ew\�1�;��)��H�Bq���3wB"qt�\D*��`U*����O$8����W�3C�6�5���x^y]y���	Г�4_z��7B���9�oIYNG�Ł˺��{Ա�z�"�/C��D*W����u�;�&���{��d�8�	�X���ϕ�[�}�]�'���"�e1�E��)���w�'��������7T����r
q��,���5��X����[1��.��J�R���ߡ�����ժ|�?�ud�D$]8�l�e�e���P\V�{�����y�:n�#��L���d �Q	�2T��Co�$V���Q�<���wC��?�e�t*{,�7
���;Ѭ���`�z�Ë'��C=�(;��/�4��1Ȣ:��!��^��KĲ��0��	c̴l�'O���Oи`��	�j�qp��{iCi��ʁyT^;C��T@�(�t�~xm��-�7&��z ���T�G�Z�i�9�}��ί�d� d�O����I�|�c��!������=��'ҋs��ڼ�<Y�x%�3�`������ۥuõ���HQy]x+��{Ae��a5�7C�F�3�����~��­!�	��ܐC	�K	"��&o��s�xqF��2-u�ia���X��M&�^�=�#?�I;��`�a��~��1ި&e�ZlN�y��x5&����zM�+uD�V8�a;�Y!��W��,RFr�^�����{T*�}�"|n�F/[GӺ���Rl�ҙ^�Y����Vx�s����Ӑz0k{��7�ͤ��zA��0DR�ϛ�q���?�9ۂqeCN/ۄ�#'p|�P�q�e��(����g��O#z�O���'���qD��=RY��H`'��x/=�W��[!���J�����mb�,֋^�^�<��'�@{�xȒ?��DXh����|����By�u����<ﭠ�L�-�OE�^y�q#��N]�!�3���,y�f��!	7N��� ���^Q��6��#u�rEϗ<3�Ε��c�;���g�˰��:(��P����y�&��Û5���+�Y)�	�p�<��2��>?��"����e}X�b��K-ţ�e(z&��T�%1�I���`�k0e�E�,���	H�g�a�2J��K��xF Ý}N#�K.�oJ�ߛz�',<O�!��ݫ��A���*�{�.R�Ӑ{'����|�G�����"��Cdf�ۭ�P4{(�?����Wa8dYPT�����g6��{�;WnW�#���xal���Z�z����/&�C)�u��y9�a�k�9������!�\8ҷ����$	i\�QeC	vƪ0��=-4��IGN
od����&�e����T�,�Qng�Q(}��=���&�� ����b^�{�M��`���mŢ�cf�K��.?�5�tS��`���8��DA�>xa�G���J�)���Z;�$�s&�s�s!��JT�|D�����qD�A$A�M��@���Csux�w�J�G6$
�W6C~H
��fZWdX��p�;_������	C�Y�����MAFH,����-��1]��X�5F�uF	���F�+0^��,O_�p�FOW,�3x��-(^<po����"���,��S��ra��I�l�
�w5�ݷhE�O�>�J!=�:�۠��5�R���&������v�$t5�BϪ&�Jd���K��O�y ���-p��W���[;�!=8���p���U�q���J�~Ȥ�ac��C=�6uBo��#GD�/�������g(��\)_V�W�7�@*?K�F�s\���/�Qqż<�<?�<�8��%(IF����!Y��P�,!����H�����)�b��v2�1,��b/��q%}./��å��Ʋ0<	��;'�$p"cJ����T���v�iZ�n\TI��b,��5^d����Cy����]�g*���<���y)�#|��3�9��n#����߾j8����e	 9@ƿ����dQ�beឥЍ���+������Ё���f�+�����r�
"&a��w�yv���=AN+)�Ľ��E�p%.�@��4 �D�����~@#啡b\/^�7�r�dy5\)����d���#�ŧ��|
���Pp%xD���9����y������� ĐT�n����´LJ���y	��N!v�~��q=.m=�G1��<�`��"E�z*��%�H�{C�W{�X�,�{�YH!��\����D�?�S�8ovOY�-�~B��yOE���b��t�4�ȶ���
�8���������.\H���=8z,[��Kqc�J������5p�.A4J�E[)�����^�ܷk��@�����æc��Ct�������y��0�~�k�ۤ�9����{Ӫ0�G�L��uW�fQ���1��[ً�Bۖ�����d{��l��m{�O�=��?��#5Ni��b�)VZy�-U��=����ֶ��Ž~R�`��7F���.�phD�V/�<^qːǀg8Tː�^>CAu�W!�n��G
�J���񢁒�,5�(>D�Ƶ��G�\��]q� �_}��"���:O1D����|�rOCi�.��r�}�R��a��tc�����s+��F��p���e�^�F�<E� ��Y؃7Qi'&>Np�BG"鞵!��qɀ�֎߼=��s[�w_�mqo�+��V�F�=>�b��:'q�mg����vb!�7fV�����S_$�:�c�`��z��H:L�#̵�C ŝ����
l���q���8�a4�f.��6�q�Z�s5-Cq�ԥ/�ĉ�qIS������Ǐ��s�ȍ�K� O�9��ׄP�����g<1�{:�� ��2�Ȇ��*ɓ���r�?��`H��/?I_^9�PcSJƿ��h鵤�z�yE���3	P�����3�Y0�G�L������*)/qg/ǝ�%��U�XqL-&3�G�/�ְ�u�)����7�~�K���S]���B*U��'���o�<F�cJ'�;���ʥ�~ē��R� �fы2�ҭ9�l�Yo�舸��iRoS��mH^D!�r����/��Σ����(���w�����@yD�׼��>��/�A�52�9��% Ň�-L������ʁ_��Yď���������s9YJK��</F^I.�m� WѰ�NO�P~�#��B��TdJ@��kx�Ω�e���ފBd)=[j�_��'yG���=8O����#�tZ���:�G������N#= ��/!3�n%��T�Άҝ��b�&-�9���m������&���V>r��4�W\�����Y�����N���\H���ͺ��O4��]������NKNSC��9���DIa�pIf>Rv�ƥY{q��j\���-Fl�_pa�F$-BQ�-��i��5��X(f��T�d�����w��sq�/襥�!�6�OMCZ�]܌I@��C�6m5.���=�p��8�f,.|6��g"��R��9���YRyq�N>� =E�3k��\���Ɣ��e��/�C��,d��@zVn������3qbW4��[��~���ӱ����ڼ?V7�5��`c���q�_��U{�����!��C\�y��g���LyS.��_���u��+��v�(��1X4��<w>�
¯�Wa��)89p ����j&�ذ��ƃk�E��Dݧ���(o��w�.N�S�����fS]�� t��_ơ~�1ױ� +>�`����Tk�%�a`k�#�:��Wa�^���N,�1*�,r��)�}�m��5��krL�:8�5��Z�ę�Sl�1�B������`�.5L�{��HR7a�GK̪��8��Q5��ɒ�ɽ�8)�Y��e,�c��#a�@	>&V�G?U��91o���^�,lp���-��ݩ6n�'�ߜ�@�Hi�byZHdK T�	۷"�Q�k�wE�_]`�����Zx����A���<yN�8���l	���q%�s�M�?6PDǘ�0�B���Ͱ����y(a=�0�2t���p��|<�I*�4?��m	�fv�{WɐP�+ݻ��=v�3�1؉yi�c�����8q�Z}�V���|A>�������Y�mTb/�E�"n����4���W|GT�E5S�|vR�1�E�nh�9�����������_�}$S<.(�8����C�t��.��D�u]�j���!Bw� 2��{Cy	w��4V�.�8�|D�tn��W'{��,pC�����o���w�y,���%H/�=��SVJo
L��|F)F���{R�� �����^S"0��,�����Bqy�A��;����<�6p�Jn��QJ
����C���sgU  ���A���Xm[	��-����3�
/�'��������t����xG~݆sE:�x7�*��ɘR�Q<+�s�!Ǖӎ�i��%�=WD�3Xp��Ȑ�k�<���><���g�=$	ER�q$P�6�WD���Cbp`�j����6�q|2}�"5n����"�y��\*��./��y/�q�A�"œ��tN�۹H�����p��l��v2N~3	�����_MǙo��xש83v1���.�D��W�3�B����$��DR�W��E��J.��ѱ+����r(v4ꍝ��aw�>���0��v���3�0%S�a���6�RI� ����0h����e���C�BZAT��ԶE��5b��Áƽ���p�t��ȡ����帿/E�Y"^����p�H1}c��rz�����0���9����8�m<���/g"��z$v��!�����	37#j�:DO_�CP|1�zB�ܦ���tJH�O�Ao���q�.Aݽ�p�A/+5i�"t�:��=�!��[����8��-���y׎8���?���+��� ��L=��qu�^�t|]��S�3�����9ٸM�y'�R�"%#7y˔�d%�ƉU����w��Nm�е=6��������)6x|����ng�l�+��=sH��1H���۷�p?#K�9g�Ł�����IO���_n�xK|�y�_�	3������q2[����c�p׎H�]02+lc�#w�$G��ݜ��u_ �������e�TtW7@/u��zű��e$fika��N�O���xbv�"�l���;D�K��� T�r[� ��z�3H�w51zx�S�k��{L��G��`йb�J/F��'V�fm�����yÍ�Ħ��M� ���Wϖ�z��2�����&o�\�t�ا�x��w=�a��
G�l�������d8�����8�g;v�i�Mjg콐S�9��5�s-?!e�^�@^!A/ʐ!rT.(���}]�W8b���(0�ѧY�W�� ���X@@5�"3^넱<_�]h�����9�/�_kK5v/Z,�6,��l��������φ�+���q;#]�c��Б���_[X����XY;X炞*-��jЅ�n7�'�a?�|3f{4B��������a&H+��e �i���oqnW ���Q��AF�H5wB��3�t=x&.
����p�N[�5�Zmy2N4� 2�1�H�$	l�Ps�L"����'_J/b9�E�Ʊ��s	�o���u��X�t��	ǂ�!9�"PO���6�½B�'&
�F���n,��+�
�щ!�q��J�y������q\D7)��EI�mdl���p��(D7�km'#��l<��r��D��.�Qy�ZJ֨\~�S����>����O��^R3�ƕ�Yx?On� ��%�n����T��p��"D��Drá�8c��RQv!bnPOZ�]��	r^P�R��+�ƈt�����Ҍ�Fl�B�9-�(ϊI_�$zy�!<{Or�p��X��`�.Z���q�� D���]'��롈u����3j��b��tiH�启TFDY�g	}��9y����Xon�qeO}��oј��sqH�|"�� V���mk\T�k��#V����Ow\�4)���q�3=�qOjt��P��?S�9OYw.��u!����H�M�"T�	"5��h�p���i�3ږs�u����}��|�Q�,,`p�ʃ�����@��̙��Fn��Q��~pŮ�۵�E�:�fv��[�Z"��5�~����q��<��~T*%ݸ.q��o
��B�W�U�%�	lC\�1�t�״��Y/ <	�'"�����+Aݩ\^�C�� ���o?W�o���T<����Vx���H���	�0K~i��]M��+wn"�~2/����q��q���UqP��V�pԶ>��f8���.���!�\?ǩZ��a2n/ڋ��[T0���y�����fee�9s� Hg'^zS;r7�_�Ni0�|3
S�>�@c'L�v�R�:�6��N�6�ka��[�?�&�O���XU��h�G�/���<L�Bfz�Xx"�vy����_�,���@`��H@5}y�%H�p��a�O?��ys�v��;{{�oĢ1}q�˗H��	�'�:�5�@Ѿ�;y	W�E'�;��_��T���d	ĳ��@:=����S� ��qa�qy;;����
��ɣv�y����|�����QBNH���B��� �:PQ�ߒ����.ʻ�q#9	��
O�$�zO,�3�1g3Ԏ�&&}����v��I������\��� �x�-o�R��<y�r��Im�T��^x�� �$�(�{
���\�_�<6�u<I�{(���d�Ԕ�8�a�u�?��U��gC<�n��zBJ�ة�͐e�˵q�CG<$�e�{B:�*�z+����`�6�U{���;���U;�@a��X;�<����	:{��#�srC7�=� �;�z��D����o���A��ˀ�ir�y�n߻���t��1-,��^!���RE��=lTbƷfJ�q'��q%"�mǢ����M���mj�a��[�N����u�����E��l�I\�8qf޸S�	7k�g�0�6��eD�Gʁ��1�m뢗gkD?'[�륒�嗇%aO�!�"j6	�����b���n\�%̝�c����r8a'`��5=d8���kב�s7x�'�vg����S�#+�^������301��|==�R��Ho����G�Po1��I��>���!��+Ī>F��s$���"�����Ɉ��q���9'$K]~�'��� >'��s�!�n� K^�Ͻ�L\
�E� ��0�����x�o�D⬝�����w!2�F���C�7a1����XjL(}JH9�!yUJ��� 'A{�^B���������Ĝ�ω^��n"n�8�k��"�Y��|��F�i(���� ٫+nyw��/����(��DAqnE>J2�R"t�0xS��o�A�Ӄ��Xҝ� }���1�S&�=�o?@��-��gL[�Qs\7n��up����#s����ܐ\���8ص��f}pu�A�=|$��X�>�Z��,�
���#{@9]�U��_q��حh�(u3�WuAb7$V���8W���]Q�Q5�b�yC,��;VL���{�νJʏR.p�?p��J:<����C8Ѹ�l?D���,}q��=οo���qE釨Fmp��ķ�3ޭpE�.{P�nr���Ev��
y����>���X*�H[֋�P����0�-���g�R��I�&�Z�W¼I��j�R�S�
�7������'d��b�GD�[������-@[�t,� i����0|r*�(/�����VwRpa�1&`r� �.��琭�*�଺"�up��G8(�k�Cc�;�p�vk: �ǬD>��i*���r-�įI;n?����r�@�W�J�f3��zi7�pr���z�x��ώ1�H��6�Xm熝j7��;w��{b�glt���ͱ٭~���?��7��e�<9���N�n�e����P^d�sW�9>(���ylݲkV�ů˗`��%X�b"OF���X:u0���q~.x������}$��N�CRx��p/��-��Ŕf��A^���'���.R]��p%qױ����v����聧o�U�٨1��Z�r�t<T܊ӆ˭0\ �D����~1��}�9&z�c��s����q�d[=f��#`��=x4�� ��y�k�⒓?��Ԯ�<��1��F��� �LC�b(�U�{�Y��b�:��:�箸0y�r�}��=TX�n�Hƾ5���g'��_��\���T��x�@���b�z(�xW���0���8!O�
<���b�<�`�i�~��}�pv�vl��Lmĸ��&S��a�!�xõZqqG[-ZS��'�|��Q|W��'Oē*)�����M�u��ii)X?o.�YZ�k���*���ϲ���L���ʻn�6��e��= �j7C�����V�ҔzF
��^x����7l�9�K6�^��H��ᲱWjꐤ�Ai����}x@�z�i0m16�4G�zmq�X���Rc'����5��1��/7L,r�����'�c��Wץs���U9t���&c�ޥ8�)֬��I#{a���ص~V���Ə���!T�JQVJ=K�Kƚ���b�c��뙜/�c��sl�{��e@%ap(xL�)�>>�O����{2�G�~���V�����bT��V�#��Q�n��v�s\�1ѻ��8sMx3�\�UTk��9}^����6�r��u�W!6cfw�����H����_�^�����E#�t""�N��nC���
c� ��$-ށj3���3jL���<�ٍܠ�}"%Ϩ�Lٓ'`� ����a�${�r�͐'���Ǔ�8n,�����D�a�܇އ ?49Aa�9��~6i?oƓ�<8���KW�<K���݅�f\ND��)͝do �*�+�C��V(�����b����,$�^�����i;Ę�q����8[���lq�H�h�L�[U�x�Z� �:Nq�ˑ��=��� ]��]�/"o���gB�'�A!.�?�]�z��Y������jV8�)��mp��B���p��!|{l����7X:z&����{��8p��{���A
���k.�-�ɘ'�j�h���\p��",<�%���@<��G|�~(�qM�W<���⼸7�v���M=���>p`�`��XԑR��cW ޯ+�!���f*DP�wܳ)B;���o�b}��h3A��㠢�)����!]+4��EVr
�g$��@Q)c7=U4T���/֍�G�V�o�S����s80r��j��*<[w��vf�����8n[������!R�%v<��@�cDxŸ|�؏���Ԗ������˔\*��XPA��^�#�n�x���B�ͻ��5�F`����i�!~��s�g���j�W[h��Z��*,׺b��/�:xc��/�Sۺó����>
i�	/�)���B�g����=0�
�鹸ؼq7�/Y�_~�	{wm�夳ؿ{=��^���wc���6�7���K>��*�x !dǂ�b�!DF��M��?ͧ'�1�{H����_�=�k�0����7qx�tq>,�j1J)�l�)[,��lЧ�99{"r/�2%�M�H�rc^�=|Sz����1��1dy����#>6��4���Iy4��U����c��S	@yJמ!c�tb�m���#̫��7�t\A��"����A��8��Ϧ��'Jz%��͏��!�=�#�s����!1�![{���zUy�x}���i</���~f2�w$���-��-6��A�"��](|ס�f�GT�x�!���+$�㍒򞑱�!�[kJ�eb��j'�h���#r�.l��3?0�3iG��jgy����`���P��=N��+"��W��2���<\˕�㛞�K�ӄ'�!o�E���_iU�TJ+k��v22'_t2Sc0%���[q>�����!�~il%v��F������.����V8��g������掸f�������
qt����@�&����W�bX����ŰƐǆ�!*7��r�PXDՋmKy�6,��;��+ѻ�:��-l[�Sǌ���1rd?,Z4;����fԍĔQ]0�_g�^�=���3N����w�ΝW)�%��)� i-{�$�_����eO��!/�1ACoe#p�X5p�zC����"���)[�l�Q�
�P"�\�hK5Ι�q��)������B1F�;�%m�`X6X�R3@��������$T��-��58>`n���3�; ܩ!�|��i?!v�8�MW���Q#�!t�t�M[���G!Χ#"|;����Lҍ҂���(<o�<zv��-���R�QR�߲�/I���m��v0��QC׺+����O:�@���������F"f�����;��c�2u�������8�G�P2tJ�ޓ0,��؛'C�!ǣ��8�/o>���qֶ��T7���t���Y#�Qg费�fZ�֤��j�(G�5� x';������ ���t���q�:���Ք��]���P�i���h?�L�a����8YE��5�p�j������f��K6R�0A�v+Wl��k��~	�NY�e�P��O��Oy��<��݄3��"éRM}W�	�
$�;	��j����A@�O��CjC��ל:A�p��/��/�j�;?mP)!�(/\zS�ϸ������;Ng��r s�>�i�I��H2�A��-�a�n8ۨ-��ö6T�:NƑ�ñϣ5�j��Ǩ�pj��m���@\�yw��tdfe�) \�^��r��@/�5�e?|���k��i3~����Mq��'-�Nh]�Sᄍf��g�3v���E��"����pE�_Q��q��).5���Pp�bN)Md�s������y�V�<^«hy8�����'حi�}�u�������Cy��Z��T�֙����f��[H�MzO�<O�t��}���ޥ�|�����)�{n�9�d�3��]�G�x�o��Hlܰ[6mƊ%?b��U��vgO²���O u�$4�X[ F�o����؞-�@ �mb"�Ŝ}�b�ȣ�0�>~1	C��Ы�6�\LC������7�V'F��*����d����R9� A�1���p-�d�ޝ^�!���9�C������M�|�Ny4U�*�a��t�c�։��Ǧ�s��n܇��-1���G[bٽKk�\}��/%�)��0�1��-�k�̖�OZ��
��=�z���Q*+'�ݰ۩.��=@qf��#R)�����<A��N��ǰS	����?�k��;o↛�~��R7�^�Ip�]�Ђ\�GO�����!/��ϵ�x���7?�z�}�D�m�Ah@0�mݏ�?����D"��J����<'o��F�}c�Ds[Y�Qd����*�Dy��Ű���ca���

�K���� �^&2xo"z�i�<4����I��k�P��-TzZ�С���[����z�7�>0��&����bG� "��j/�X:"�`��ʯ���e�Rt~�j�,�ݰ��m/\W�"A�EA�=�Z8����f�!<:����2�ia��c��"���/�#��ʐ�"��D�o�0�g'ܵ�̝�gMǔIC1e� ,[:;�`ߎ_�}�|��?��Ǭa����d���8��G�rpn\'���s�2�Ȑ�Pgy�g2(Ȑ���|���m��ؼ+�u����p���UԈ4� �zE�S�H�#�� �L��vH�t��u�ڈ�n�3��Fڏ�ȥ�m�hs��a��p/W��.1���%�8�����!��8n^�t�E���Թ��
���H�?.P�����P7@��?��#��L"Һδꎬ-��**  z*<8ba�0Bdrzqɐ�Gi�S����Tx��W�!{w8���y�Op������[�T(�J��x!���%<@笼qYW�������-�!�NGDv��xv剼4�<�_x�����������Z�a���2q��L�X��U�x3wD9࢑=��EմA��q�:����T#��qTg�)E����z8\��^�%��Eܹ�@�J�/�3+���_�H���	ĉ�	&�"����Bx[Ę�Q��5�e�ĩJ�(3�#�l�f����c��p��b1F��p�۞�����wO�B�a�׵�5e}\4q@tUK$Yh�F�"�H��5�pY�m���Ek�%�R�	�RcC��ٛ#n�;`<�L�lƻԓm�9��<�T�g��d$���8���|�%�\q�`�u��ס4\�#.nĎ�d7�BĒM�;
���"��A�@����K����Ӗ!#�u�y��R�p4����)"@z�E>$�IK
Cp���i�1B�#Le�(ل�
=��8b��vZ���qC�Λ�gI�p|�ͫ���m֤'�/�z�@�,*g{�~�֞���{�ef����$3��<�i6�′6vQZe���5X`b�V
�V��U<�i/5��U>�C ������ ̧��������x�](��Ch���]��,w�y^��]��{��"��2n(V/��1gq p7�DZ|p!���Ӛ�S�o⋒��qp�FlܵkV���A����9l3���Q�z�y���GM�X��Ы�/}3H"p^��\�����e<��U����b|gd��{D��,a؉!w<���W�BH]�
3R�7ۘ¢|̘4v� }��0��	��i݄W��N����m��\��Ryɿ��j�F7��#��`1�5�n� ��2�=��
�<��K>b��:<s��k��i�Vz�8��8u8�8�{7��R�.�2�I���
�Y�+��e
5(����#ݭ>�:�"`!H�Hg���$O�!�3+!�)&��)\�G�a�5��T���N&�ه*�ؖm	�"q����d�[٢����'p��b��=F:��A_�*�����*<���A�'�h��n(����<>�~A/Aފ	Ѡ��+m�E���_�COsk���T!�|���#H?�_�}��7�����SMT8���5�R�8_��,�^H���u+��h�@��յx`ဇV:ܪf�b��#Vn��U� /�
)]�'��(}.���#�|2x�p	����:��" �k�G���D̻[�|)�/]�-��bάј�`�/���~��58�c%�-�j�Y��b��سv9�p�h��؅Ғ��܆
ӅW�>���{|�=z«G���k��0�Mqr�d�5�7�3V#�\'��5�$�`�c;����Ʈ� ��Y]sD���㈔�	���A��>b��ӗ�!����=g�����q+B�Mp�����RMnQcr��5�޳��h�@��{�H|�׫���:$����<p[���uq~�x�^�N��TqJ�GO{�������,���xX��y��ô�)��@�M&=n�]�ĿX�b%.|���j\��
7�詜�>�ƅ�UH��7�s�u��fK�y���#QNdȓ�k9�!��%�q]�����"�O`�o���'DV��9!ٌ:25us�W-��̜#���M	�X"��S�Gl#��X��_A~�T�x�Gy	����W9���+D��98�h�sU=	�p�}s��OpW�'�a��3Eh���'���Hu�Y�����VK��yc�[�m��~ڊ�Gto��_\�X7�_���8:h"<>�{�p���#����DϽD |�
(Ճ��C֊��5f&v9��ԧ4j��6�q·7o���� I�<�D�㖢<=َp���^�:����!Y�)���W1�H�Pj�6~�I[wb��X��,���f����c������ +;�{6B�[+������	�}�����[���g����)J�%A^i^N/ۂu;#\��ZH�Qk=+����	;t�9#Pi�0A����(=	�%�w��H�8Me5u�j MZ9* Qy�{�M�k�$�!��jӳ�� �)g�gs�]��VʷU���:y�,�c��Aj+�w�u�Hv�=�ϥ½[��G���F��.�������R�+C}�x��;���8rx��c������[|�i��>N�}�GN����ظ��'	����p��_�
vl��͛�c�Vܼ~C���<R?�A6�������yc�']���M�ܴc��a�ى�	�x#�q�q�){���i�^� +�:5\��8���y,��%�q�7�k(l{Y8�i���A���}Lo�S�F�k0]�.����c��#�Q�:��ª����,�RM-�z�H�aa��w�} 7_��{�^:9y�V�<~�@��S��T�F���m%^Ryy	y�y<\��sB�6�'
h����;������Z����+5�]F��"ã1�R�I��@U�4�R�H�vD6A]��[,�( ��yyyy��w[��!*O|o��8%Qq��y3RD�d�Q�m5�ѝz<�	�xo�<H��0g7t�ĭ����յ/5��D]�Q�){a��Gƨ'�^�1����G�o
�WU���h��-��0A[�XQ���
�(s�����ab�9-��ţ�p�p0�Poz�_M�-�HGS%fPCuF�%��oU�����	����+Գ�f�$�']#��n�;���F�#[�Y8"���p��1�qB7�>|����Ky_j�����?��������p�y���|99������+B����.��)#��O3���W���k	!Z�[��e����aع����8�[�7G��'�]��dH��ȯ�"��:^,"���������8��G��c�xP�n��	Q*����u���%�$ �t��$s�����xἅNSڝ��i3�v%R�}[`C%Ë\�bx\��Ĝ=��V @�B`b���I�0�ſ�S��q�@4��<�o&�����P�rnVw&�"��	�L<������"��iQ9�P-=�˦蔔��:���Aa� =���9E((x�"J7�[��2�w����H��G�WI���_�'�R$` UU��U�8W�ฺ1B�����8���؞���tUx~8�7�ƒ��(�WON#1gQt,$����E�oFq	�.؉��"��J�c�{g'�N�
�I�	��jhN����頻v8c�s_��i�����6(���\�Y/��������xC��
�9<<{[Zt�i�?�]�#��ǌ8E��&]��duN�>'k��Nڮ
l�Fz���d���c�϶ыp71�y��U��W�1�44dEc�~bA�e*'�����
	d�/�m�L������s��N����0n�[��d?Ct�Hk�۶GL�f��	�-�$:9�
��r(��9�a�����%��5F��h+=�������Kpz�,��E���@�GZ�C�쟰��@y5�	�7����KunN�Q�}��X��q�n���b��=t\��P�����Mg�Ca�~X�`�/e]�L]p�lo���Z��[�	o�Q����{	��v�)�;���8���u?G��(��"�CLנgU<��S�Xg>���PZL�UT��x|:ە�˂`�����֘Gvc>�
K��hp��a!6N8���^j����}-1������-��P�8�E�������;n���ሕa���U�T��3�u&�{�b�Ϙ=e�vn���� �|8nf�D��c �����E�xnT��C�ƥ8�s5މ���b��u8�(�A�?�A��u�Ů$�V����N��[U7o�	rbbQp<Sk���TT��[�b���8�JN,�ۜu����Y�A�̣��p�/n�rM�p2�(񸈻ے��߱7p��Ep��
:�x`Q�1Il��[�M����Q;`$u {P'�N`0D�%�`Χ����Q���Bq�3*{O���5����9}W�u�S*O5����	�@��Y� ���:��¦To��41��.�ܾ�C�a}��XK��o�h�:H�l�����G�Bdz��O�{��}!�+nm��k+ Ͼ�ܚ!L���"�So�exzq�c�c]�#��Ra��#�Ubi�a�#��Lz�9�hk�#�wQ��jXd������8��dov�YnX��ۻ����U:�+ɓG�ׇ*j+l�?���H��Bg?��3Uܮ���)mG��t�Mj���R/�2U�˖B�Y:�a�J��W�1L!�K��G�E������r�#�!�z�4
�˦�%;���hs�II�8�oΆ���X��L?���qC����-?!>" ��O">|vo�������>���$ǝ��s�db��0����x����vz<����e}HX�Q�z8���ݓ�"`�B��z
�;oDPG�x��	B�.�H^�K��̜m�X����gp-]䭜.o
�qE��,!��L�E�{�k�b��+bu��]����\�9��ȐG��X�!I�Xj�"�pQ]�! 4s�ꩇS�z�Åe��ޏ����F���W��ի���O������y�]��"J?������a���M�y�����]�^ޙ���	fZDT�*�:I�YS�p#IN|񜥈�;!��)	�(�DCB��$�Feȓ>��<�MC^^!n����Z�v#���x�=@<���� #��k�q��g��(=	��j�}$��+�)S����)��ȣ�J�O�]��P����f8��
��y�/�`�;N�s��-B�q�����ԁ�Ki���kZ"�F�#��Ql�;��X�W�[�P�T�1C/�ኝ�� ��$�F�TM'e]�t�s*�V:�d*C&j\�9zdk���W�����f��g��+B� �l:S�-�]ϽVix�-�u�y\�y��Ҳ-��o�dۺb�L����ӵ�lS�̕��c��/NQ�&�lX�_��2[��^�&X�8�uE���� �m��D	�����iHM��zrV�)����%�GQ��j��|E���(��Sg�!o��=T�w�i`�:⠍^��	�㔃©����N����'�œ��Y������sߔ�z<��iI�	�R��w�,v|��u����fs-~$ݾ7Uc!�
=�C��!
{1��_�]��?���1�7�	��j�cCj�WBB���Ceѿybn2�.5���	ĺu�a�J�ܴ��,G��ߡπ���eY)Ta��ܐ����U �Q-<>�q!;���6�޻�vnE\T��>���G �YN֌��I�_���:88�J` ����K��A�j��S���f��c��=�ht��G#��m��M�JKv\β�r-.J�uQ�)d��ۖ�f�nhbf���`�������jG1��O���q�k{��i��->ƃ��Ԉ��&������o悩�^�D���(S�p�}�!�]Hp'A�X���!��%���K�<O� f�Ð�r7C,Q���?~O�Wk	��"	������q[��n*���:�.�G6n(R{�c�˧B�=�[�燈!@\b����������X\>����̦�c��+j4觰�@%�!��P�]l��H��_�`l��xF��%yc$��E��!W��,<��=�+b�-)$s��Q��k4z����ǻisO����(4b�x��-zj��p%p!�s��d���>�Dw=��Tc5�-���)�7�^<3=sIx�!�g�^e�KW��AK�m���H����(n��R@��=y9/��'-f��kY*�c��!8�7{���NFT�1DGǚ�?a�!�>c2�!���ȑ���=B ���W!��f$���;g�����<�U���n]�����R��#Ò!��yx� �_���^d(NM\(�<�pm���qh��8�D�A���=ك��M�'��/�Ҝ�����&���O��4"���pe~K0ԛ�>�O���RlN�9��[��ZM�����`������G�O�8�*�1G/�8A�fO?���S|���Y�z�t�����O?S�����P�,eOyˋ��I�'U(���,�nE��PL���{�6+W;��	_��{ ��	�ݽp���:�,^4Q"��%�U����ɐWz�@����1����j�hI��IuCjT�����PD�qc�'�?'��ob &@ٿ�E0��2FQF�F��<=���w�@{�TY��5T<y>\��3[y��}PvA(�~6�7�|sj�9�פ�g!y�,�6D��.T��dU+' =A�s��5�)��?��q�@�� 	&xa��N@���)Z�p­>N~�[{ME�Γ��bX�*�A�����y]��r�q}�
�ti-�s&WU�L��L��FdUk\$����N�qd�T�]�{�P��5�cE���,pVAq�ϑ5��S�C���]A��r�'�}q�z��?��)�O��œT�B�N��@�<c)6����>��ܱ����A����b�sC���"D�`'lwl����"%�<R3�#��}�X��k�Cz��b��I��q��U��a?"�w���n"������n ��]T���l��p�a��`��q�g}q��.�e�E��'�6f��q�g�,h�Q�����d�[�_�rp�n6��`�G���Z���Z�la��:,�vk#A�s��� [��������C6�8Lm�j_����}-�ƅ�C�?��8�6?lW�RҰj�fl_��7�����8vl7�oZ������pp�Z 9W�������1�� �NP�>�7#$,����������G �E�6�'L�j�A�������d�����0A�E���j'LT�0��#Ŷj��s��z�o��u܍���wƣ<^�MA*���p�%Q:r>s-�}I/^L�g�@��{�_��`��H[��\��o����)1��{��R2�t�Q,q!(����V�Q�/���Q�� Ε �OYl��=����
�{�<y��m̿��?�g��BȊ��ql�T"@�$*C^*A/��C�5�#R(R<l�C�����x	�+Pz�y�*o����]`�%�1%� �Zë�~݁�A����0�r���6�$����5����_�0COz^[2���jl��'��T�yx�
�y�
�W�p��p��+o�̇Z�/��5��>��ho��PGoT9���yd�.N�Daf�au[���=xq2
����P��@?jX�P�����dL�n\'c�"���B�k��^����7Ի"C#H_�ŋ.#����I�.�n�:�R�+*��"7:g��,���CX�z	zw퀖�bЀ���c��;`�Оۏ���8~r�߈S�[�����x^���EwQV�����p=9�����M�K��� �n�7)C�<�+ ����y��'���w�y�]k���jyȖ�f��a�s��2��V�A	�Y�@��h�Xc/�7댢�(R�+�� aHX?6�N�g�c�ɳسr3�݉���°ɸ:q��,��sq�i�ph��"�&�D��6q���w�.F��_�4d�|��C�#���k�Pǂ�	���D����c9T$��y��Nb�+]ˣ/q��E��u<m� �cw�/��3g�ތ���s8�X:
��j�.d�8�X�"�(#�����v�ܸ�Cܜ�dp�Dǈ����|d�F�뛀��Ex�]�y�g\�
OęH�P��:�,*C^���kZ��UNU��)j�OS]8C D�=M�FQH$њtZ�"�ܻ�;HO�m�*UC��x�bu���દ8��9��o)@O�>�j���~�kh��+�f�}� ;�F���`[�	8�3�G�E�ʁu�?b�9��oW��<$�g��q�:�W(�8].Z9!� <����8��-��G������#py�a��a�M����5#=�Q#r��6Z!e�/��,1����o�3�$B��J���9��~9ŗ:&�q�:8����.8�k���+�-�~ơ�#�{������^��6�*7�ڹᤇ?���g
o�_ĝ�YHM����{�ȸ'�!��y�r�#3�q��qq�N����/�'�1� �����&j�>B�0wzX+pT�*��Qԉ��j��Z!����I0\�_B=��WZ*m�ĝ\q�ZZ����@��m� ;(��t��va�����u�n��=��l4TOm�4�=��"�Y�P�D�|����~��[�w��!�I��$z}#������Ћ�S�~�N��C۷b׮�8pd+"�B�~�r�1 �;}��	T��j�լ������38s� ~X�+7�Ì���׍x��+҇4�]�?y�����Ђ����	�(룳���
._�è���#���%0bb�!6��w��TL pee�~b�,-0���q��Q�D����<����t��G�¯�C�"p�\,>�W���]=�1� o�Z%�F�)$Sm��0�l�3�g��`9gc�+)��g*�����#��7Kl���v��֞xj�, ��W��Q�,���޾�*�y���+�p�+ls�C^�#1Q�'�f#b�*�l�;	t�б{��k�9��-{���!�'��&�yn�=^�A
��
������!�^-Ĝ��V�ET>���=�����z"���L����2��b��Zl�ؗ2�7�dh{�+���	��WCS�m�B-�h��q\���_Bר�d��W؆q�(��r!'W�//�`v۲_����jZ/^wK;�4S��3ݬm1�t�`��p{,�2N�C��X]�V5�§@�*C�Q�Ab��׍�p�L��\'ʿj�%�����|y7��r�ʑ ���8`^[kq���ł��Ü�T�\D��=�a��,\�x	=�׮c��i�յZ�h���h��'����p�����}�wF� �N��+W�p�Z$��-�Ean:��#<-{D=�{�ʸ��|��1hs:ӫ�.,l4�@q���{A��<�{��������fa���8��ʃsd�ϙ�U�ˋ�Xx�(�x~W���`�q��qΈ����VݑK=�w��Ax�Hd�d�c�w:
k.��_����]�Z��?���v uG ~\��&�p��x�r����Uȝ����p�N䆜��I3��h9��}��8�X�QG�V�/X�/)^3�d�N��|=��7_�d�;�:��=�DƮ�H܏�n�I���'���p�x��?t�kŞO=���<�8-�Qǃ����7�g�G�.N� Md�2�Wҋt���sWy�����8AfMk�#�D�<CO޹<G���FyglK���i��Y3N� �����?���:w$8����2�� Ғ�<,��[�E�1�~b��!/��B�Y#�:�J:��<~bd' o��]d,�8@�� �O���޸���+��J(��u��.�ƺW��;1�����h+��2/�H @����T�P���[|�[�ƭas�[]	��b��/D;��I��pg�J<�z��O���+p'�*g�^<ڑw/G�.D�k+�Z��Is'7����5C��pkO��o���spv�l�^�����d��vq�b���Y'�tA��_p-6��R��y/���/�\������Ian�FX�o���x�N�jq���	������(����U����2��:�4�c�{��!��H	
㇈�%�Mw�*y�/�`�#��G@��f��X����+��m��-��e톃Ԙ�r�1��C*��� �'}�Pz���ZV���c�_kĬ܊��R'��\�^�9.a�����G�΍t��w���`�.�ٿA��p6:��8����Y����O����5�q�vs�0��G���I�oѴ��X��<)O���Y��׉�_�SD-݌�-1��}-��f�ǉ5���)�-uvF��0U儁���)�F�[a��z+���tP��8�i�R��Ϡt�<B��e�ӳ��)��n]������G7LiԐ�~;Q�`����]0�F��V6bd>��ٌcç�Rv�b��XaN�up�0[,�NY��/⹅���=�8�1{�(�y>)��l��[I�� �7��x`�n�����GZ�� '��HP���l����'6tLOEn�C��-����~���b����fM�Oe�PgoĻ�C�kc���ᶝn�y�9�N�أ���K@{�u��ʴ�tS<rk�T�ڨ1��c	��!*ȩe�0ӽ6F�0�ԉݮ-�b��~}ݍ-ѭ��X ��V翼�:֭Gi�#I^)I������ƈ���z����ld����i�s�
6.�_�y���5�����Đׇ�[��!�	�O�GF4l�V !w�/���U�1���Z���Q:w�ѹ��ʮ�QdȻeưgG��R�uS�*<�JrO�LE}2�����D~Pτ� ��z,<��aOx�(��T6</����; �?l�6�?��m?����G�Ѥnةl��� _|վ&N���6��R��QT���(/�3q�bΞ>I�G���ܳ,w���R$d��O�r�W�9qN���ۧN��ysĖ=��]
���A�!�/��Al�O�oI࠰G��I��Hl���DP��k���+�R^a��ڄ�X��aB�n��E�`�p���8��kl�0��bq�}�w���yr�Wc�'ߊ��6{~��>c��~~�k���=�8���yO�/�RzV��|��+��z�b�!���	Ķ���q?�Ļ��*2 �������<��G��	����e�c��c|=.���3z���k& �\Y*���9o�B�|'����y���!��'B'/��!/��B,\a�#Cg5�g)�è�� �	w���/{ ���aO�����+�'p!�W�m�6M3D[P��@����,Tb�Z�>c,=�����1�у5�h��vֻ�c-�j�5�z���Z���+��4�d�7�%��� s�f��jK�:�Ly�D`y�lA��#.�9o����)��H0r�1�@��i�p�O����$Q�O������f�����{�9YI/� tfO��QH�+�!�4���� ��# ���-]p���Mp�M7�4��>�z�V���si�݆#�����$������:�p��ވ�~	.G�!�4'��l+Cw��K&��1��|Y��-:��xsy��J�4l'����
;x�V�J��G(�zJ7Q�ʯ!Rad�ݚ�p��H�z@*,t���Ӥ�&���%Ý��hGS��v��g�1����Nvk��=6Q�m7%��v�Q��kg���c�`ǀw�7�%	ֺ�a�`3���#�_����-����˛T�4��&��d_�
Jq��m���ElT4N?$:���p(d7�w!$,�G�#��Y8��ϪW���{S��\M���Ӱ	ܼ|ѸQs�ش��
��xh��1��ڃ���0Ӽ6����Y���u'���ir
�4j�n5�4W��8��>�Be��3�������#�����߹y`n/�h�݆�(��H ��_���"�?�Õ�Dܸ��~��U�*�xza��������1Vc��Z=F������|�cM,��o�0�ɧ��D�bb��r+_�Vyc��}P�߳�}}@Wϩ>�Z>����Z:��%6���[!�V�
�;A�PC�c��Tmޓ7�^SAa�<eOϯ�s,�����!�6�B@Æd�4b�j�k]�sm��ܢ��fy��*�Zk|P�#أ�eZo�p��2�F8O��R�)*�(O,i������Hl�����ãjg1w������b�ަV��耶Z[����K�0q�P������<1�ZXX���"<�]�<�J�I�+�� ��I,=� �M�Ţ�Qn~�LƜ������a�"��_�wFzh<
��G�WC���m��62��j�X�ð�Գv�enREg��M���4�@�����z���V5��^]y��ΈL�!O��!<=����� ��U�#s@���k>�p��)����捚�ݧ��M���h^����,�W���#t�*�l���`��1�a�2��h	�L��q�&a��I�0~�-]%Ns �!Ov�W���xr���<���Cp�I�Ocl�9;��!7/DW�x�da �'�}��^x��!�'�y�z�W,�q�qg�e�ܜ�1T���q��܅�<�{>+}���N�-Ξ80~��&��}����	�q����Q+�B�v��� ��p��i��>���e���ðR^�b��G��-��YcJ1��,���Y�
�5��TO~�4���A��8�ր:V>Hv���_����#t����sUlq���B����F�8I��١��6��3�����a��^�/[N.�������釈��C��_�k{	ȩN�
y�4�j�c���nf�����5�:����hzX	(���3�r��@j�9yϳ
pe�FlQ5{����T_C�sN�r�3ȯ�(q�:k�g����^G�r�5Ҕ���Ŷֽpm�y�_�	|�����}�J�!w�i�����q��.�$�#��+�/)(��^$Yڋ!�d�/�������y�:җ��}��S�1;���SWH[����w��8��U�������NKŭ�ױ�<�s�g-���qʌa��Fx�*/d�#Cɾ���:_��{C�*�p��E�DL����n��ôybn^ƫ���{�� ��
ȣki�"p��n�T��<>](���-����R#K�:PK�G:�t;�pAu�+\q@I��r�Q��S{���_��9��9v��&򢼂�B�������z
��3�v#Sxv����&��'o;���5u������b'�pؚ ��s��{�]e�V������1�5r$��K�Q��B/��BE�g@)���S���z��+�����عd	N݋���ڂ_7.��u+s0 ��[�Ԣ�V� �a�[�������+t���wm��ݾD���R١g�n�c����va�����FQ�����t�,�H���Wm�H�&�ЈM�y�B��k�Y��,�ja!�r��v�
=1��W�׳��ydÿ1���A�&��M�a�nt��1��U�0���[c��c���`��k�P��pz�Z��c<��=�:a����8|*1��5p��	�M�\_K ^����sD�� ������ ��|��E�G����C��! ϭ.A�'}Fv ��6��D��{C��ǅ�W�1��)A��ɓ!oo�z�Qଣ;���r\�➲6n��"MWG,��aˠ'�u{d�\�qg��'��)�#pj��l��-�Z�0�����`�_Pr>���p�6QH�<�V�0�2�6=���kZ����:P��9���l��+>�� 	���U27._�͛7E�L�y��pt���� ?��jZ�#��2�a�b��n6qF-2S�7<d���}SP����7aw��0��=)�{a|3l�r@�{]��F25f졓=y/�x�B�uSG\�i���6�QE���!P�!{�oWx�9��x
d �C�/v��t��3�y����	���Ъ��|�:�m	ۚ��{���?����	,�0�4ҩ����AMF�q���ޥ'���
Ga�ρ$��!� ��b�7�P'��7{~�=|�洕!��y_3�[v��1ވ �X)�F�͜qŤ��A֑PI�w�V��-8=�"\N��5�Wb��qf�l��	��?��o����}�X��|Z‱	C��ކ�83j��@��Ee<S�w(OO�I�>�p�l� "�	/��Ӝ/"���e��}�����s���t\YL��zB�kQ\ME�H�c��!y+����IG�U!���F�CK	�o�gD�]4H���W!�S�;�����v7A���ȷ�d.�8	P�U	�b�jS��$���ۋE&�zaO���w�:;O)�b������{s 5�����|q��fecDY���{��K�a�0*cg�Y�u(xN ���y'�a���>Pcg55��4Sွ/�4h���¥e{)⒇�7�/^���/��y+���+9��C�z FU�l�Sg$�PY�i-m�B���Ae�=v�2Ѥ#g����"�=��_]ĸ��	��1i9p/��yob�(Iu�fe�fj����7�g�,y�B�U�õ��5;�Kz>�!����8gb�(��ٰp�Z���	R}Z!IO���Db�V��a�OZ��	�wW������<a�SR^]e���(C��|�h�[v�v^�G_<A/����#ja.5�ۜ�qX�N�VdswQG<�ґ�%0=��M���%p?%i)�HM�#�a����_ܕ_�y����!v�A��-�����ս+�3������*l��'q?Ջ]�X��%�c�;�$�S9ስ�k: ȭy�q�u�R�����jAi	�df�t|<�<�5�b �QkƎArX0N{�m߷�A�ڶ
���ښyF�Z�R��¾5���/�a�|l\� gO�'�k��<��2�^��Ə�9b��}�u�DuqF�vȾv��?��/�`�hS��3O�+O+6I�c�&S�4EE��:��8`��A,�������nZ�:A�Z�����1�0���x��t&�DP;�R�i��u.A�8IG�T��@���Ȯ���L��{9xv*	�{��JeC� ;7Qi�	t�y��m-<wl"��1�=ֻ�X�"+�r'���csG<#�����	4Y��LS�JH�R��8�!��U<�Ğ<�pR���� %"�"�ׄ�rss��&��JT�˞�Ң,DoZ����������U/�Z"צ6�[z���w^$�I��J*��T���^��4'�@�BJ�R����3�f�z�'�uMSj1���|��Ǡ0�Vt�ULŘ;��@�����
��D��ԓ��E7�z�{�k��O��Ru,����]?j�1ݻc��1X8f"f�Q��7^����u���9x���@J��6�o��hb�q{ө u$2��� <���ĩ��1��C��7�PX��������zܣ�w�O���5n�(ce�yy��w���M��B�'�������ZϏq,J�ϓ)���z"u��{�I�JY��~X�/mCuʰahۨ>�|���m�)û���	�1ux�l��j{�e]��sA�Z�����x��b��X4g"6�]���pm޽��Е�2��=�X�N6L�~_�(��<l�����F�7�g���ӱߙz�3�掉yy���.��a�D>n/�1@�6*kx#��wxD��7U�WByC(��*�-ip�%^����pt�f�nڄ���qsK ��Í%�q��/���	�F����gpkI|*.M���v��D�����M��� �@m^�çDp�H�"��=s��X)���Yx=C4��MAX�gn������1s*?լ�B�3C��ʲ�m����Np��rk!<D���#�*q�-��ذ�x��Hě!O�L�N	+j�O��^�O�[9H�:A5�Ī]�;�C�&�԰%$�ϗ���
�(%H�B@��
���f�(; T��ϿE��K�W<\�Ï��	�UI�ʁ?_�)E�����ͼq����B�,����W��� >��U��${���+���V�Y�JL�g�;T�3�j��~�4���WT�r'����˚ye�q�Qw���>�𒅽���ӍO�B�kjE��C_��%;o*�����up��cd�\#����{Kq�;�ʾ��۷o�ν�H���T���c�!س��A�arF�b.'o_�H�ǝ.^���w� +�:�B�܅\t��d�8��	�� +:� ��)�z�$`ʐFH7�]�|�E$��:yS0"(͒��q��(s���ǩ-��:�$�U�,�#�S��v%�d��xqC 5�t�8��CN���W8��V1��R�� ����~��������v`C�6��E���j�1����[`��/֐G���O6mO9��J[1t�����}�m\q���\#��u�Sa#O/d��z)C�\7_�N>�B�E��4Vw��b�},���������H�=��gph�6�nX���~x^�*`T��po�"ڼ;��cߑM<H���	<���\�������)0�Q9��hr?����Ы�)������fv�Z��"^���X����������t�C��0��3�s�+Z'R�򼽱To�x��8{�qp�hGIF�	�u��&;{c<u�|�-�0��d�B�y��*���3�jc��9��ǩ7��GH��{|�b��FZ�0��ޫ�Cf(�t~����1ݛ�*��X;���nݟ{����������V����������Wwoiqw$!!!!!�BpB�#!<�yfg�@��߹���Wɞwd��Z3����o�u쇶�<o#M|����3,[Sh�%�4@+����"���i���M���1���R�FZ ϚF:ys�'a�=��P�H B��$���!��a֔I���b++_Ѽ
*vy����N[�PT�rk=��F`Oz�`���8�˱����w�X�����G����[<��Ǽ|q?���t`������D�>Ѥ�@����8@�u��8wo%�ptBgW$�u��H6�H6�x�l���1���G���=]=�&����Oz�q]��r��x��`�3u�{p�i�6�/���?�X�N����p��팇X���Α���e���XƭyC����O�� ��%]b��u�lӈ2
��)"w!�k������<�_ɏP}��}�9�|�E���]���=���y�;�}���|�_��_>{��4>|�I|������W1�0���d�w�5�k�Z8���Gm�� ,���5�ϊm��}�A~b�.|?����ʐ$|x�$|y�5�ۑ��L�|���nF�ZB� ���V1E��S �/��i"*We�{���Ry*��*����Tw��
1�矱n�<�}�S|9�.�{���m
��������������;��x&~���~����	F�B�0r<��B��������f� �EP>�Z2��9�|�|S e5�u����t��f6>���b6�o|Ĝ"S��	�/��_Fկ�X��]C�.M�<�t��9����2ǎ��Տ���=�����5y�A��S�Q��@ގ#(��,�� �@Ȼ�ݴ��I@�����٢��ʅ����W��v�+	��W�"�#�F\�S�D:ڌ}G�b�?uU5����+�^���¿{"���5x;K�����%|����b�j�o>����%���oĖ~�=䩊ڊ}��V���k�q~)X?��	���_���D=xE]��y%]Q�9�D�s:��B��
�C��]�ntn�#7��amP?�?��9�OK:.VG����ǰ��u��h:�kמr�ݲ��~�鐯#x�v�@���;��Fm�QB=�<���L�Y���A��QO�,+7����� x(��{��PUM��O���䵬�!���o�aC��(r��l�ё�+�B�4��vqu����	�RE�Xv�����"f~-����=0����v:��r�	�Qr~�ڊ O�#�����ڟ�`\N���~M�}��i�L�O1=�m�b�I���u�6/��h�Ұ�r�jk��������8}��,!�m�����N��l��o�N�g~��%���N���k~I���OO>Eƚ5ؒ�͋Eq��H^B^����EL��|��'�vƧ�6�d%�Y=i9��+�#'�|�[��~ AW�Y��)��Yօ��3�`�
�*jF�w?��~��x��^��1g�?K�x���Q���{��TG��&�s������D{���D��g�	4c���e��7<���5��S�GϺ:�Q��x���\3���{�����X�}2>v�����x������GW�$�ii��p��k��	�Z�d�.���ǈ�;�����}�ԃ�]�1}ry{�,d��/\��e=X��Ui^�~��z��"�RVpDK$��<b����]N�&]�V��fV�N�=$֓n���@��p�^(�{�3�
�=��JD�G^��Oy��]���PB�-�Q��Gx��7���oz�].�9����'=͚��8H���G6��^�&9�CAa���~�_�	���v� ���6��=�~&�{��'�vt3�i�C �߉�G���;�;���h�1O	
��O��>�C3V"y�<����㿮4�C��ەx��+mrp�2.k����Q$�\��z�e�|PF�m"y�nyGy�]��q�⑨�ذ:״�ԝ��S�O[�3k�[�����>]�jj��v5��k�E���X1�������;�c�r62V�CƲ�H��=���~Ś��"y�oX�r:�����e��3ߛ�x6�W��-%s���Sӯ΂�D}�i��eG�����͜'9}�m�>�N�v%��.&dC��^+�!�P����׬�Қ������;	G�f����u�	�l�+..��?��̅ː��[�5�����/��M_|������ZMg9�<<G����ðɣ7��["�o�z��+�!�����q��δ��m5�4�\x:�N���4���kv�
	���O�<�Yڷ��٨�P��O(��G|�y��uE�G?]�h�DV���uXp9A���G��c�n(l����X6ɏ�������<�"ȶ���K�ڐ�?�),k��0���L�Ruzm�"���`���l������N`_�o�oL��C
VOV}I�,䙯oB����;�~�u�G�|L�s=�\�U���r%��
'����,	�N�%�Ӆ��bz�܂0/(K{���������H���EU�V��=lȫ�l>G\�b�$��i�g֚Z�<:��!��~]L�z�C�Y����f��E�i�|��B7�g��a�#��rVB;�/TG�Z����:�HyQ�`�����=X�ڿ�,�72t��.��{i�Pl�Hq�#d� ��UӴ�O��:���A��!��#��wS@�9ѣ`�C��(���z:���Ϯq��R�<�ME?7�7�&��s�3�t��uq�'w|����O����9��'�E��M�<A�6;,���P�"��O���/C����~_G���F���z�8'`-����.�&&�F������5�e!tj:�F_�Ŵ����t���c�<��;�s fDD�̉�WM��.5.u����¹��;��q fv	2'�L��0�;� �K��s�z��
�>}��i�������BQ��[X2�|�!�����o��j�Nԛ>m��t�?�d�j�U_��=nES��X���:8��v�����eh��F�<�?��]�q��oW�%�ً�����w���t6��S�2���8�m��l�	�w��c�9���g�O:���޽���������sG<5b
�ϧބ�)(�~r���.�4<�����C�{>М\Q����E��9y�42�AC;qyg"z`/�b�+�;���Y>�3�e�ͺX��@�u�*͋@��n���3�%n�AsD���b�kS�B�p� ������z%'�5l�fz.��r�^�1~���Ӟ�8��턽Oؠ����H�{!�/�w�S�",��q<ۑ�Cc��z-��������u"�;���
���u���Fy� �´��a$��GJ֔�|����]]�qg箸�K'�^'�#uv6�����J%f��gp$��*��[�GN!x쿮�4�4���Wa����+;�����io�Ⱥ����O�X�G��������8�g<�G�� {�F��ZD�y)ȓ�-�Mk���6ؤ��a��_1g�oX�x���	?|�!>��-̞�����ŋ�c��XC�[�b֧��O?er)�HY�����I���ؐ�k��h�Y;�i���`K[�3�y�4�w���5���􅅓n��;@�k���MWYPg���;x�Ӵ�v ��':E5J]���Ä<��?V=���b�<w���F�C�cAh?�9�5ס�׹�7c�LxK�l��a�y�]�DDjWz�CQ2�Z4�������t���3G��Ko.��;Q��6j2�=I�kh6��T����ԮDW������5H��8�f/ï�߄_|���o(N�^��W?C�w���fr0
�v�怬���<����Eƺg������Dg��@�j�,�Ħ���Q����1[�2E��(*�s�כ��F�c0V�=��#�5�J-G݀��������� ��Ù��o !)%���Sd*��S��^�4��DS����͢xM�-�
Ƽ�x,�;�O6�⨱���EU�V���Ƃ���3���OX2���U��鴋"1;��(ung_x�]��A��q	A�b� �^_x�!3x�<�o3un��yu�����#�sZ'ȳ�倉��؃��{���gX�Y��\��f� l���R�.��\��6P�i�l���k���n�<e:P�?yFg�/��Z����'�
���q(t
�F����H�þȍ �������h��,��f�yKX�f�� o�_"f��i_�a2g��E��i[@���/e�et̎�?���>7 �9����:�	��t���N�&� OI�:@Y��N�X���l�5�X��Ž�bߒTS���Qu�g!��s��!%�V�z��"����;��X��E��3�z཈����p�3�a����:\���8���(\<����o_~�y?|�Mkҭ�ſ����c���/q�Ǎ84����Y�{��wv$�u%@��ѷ�xJ��7�X�����u��W:�u� �ź}�N�?o�F���@Hz�m�3omy��S�z�\�Z�"APk�vp�kށx���+�{'<��[/��  ��IDAT�'݈���8�����L��VFL��]b� ��;;:���'���5����^���<�̶mym�@^�٢MZ���dv�6�wǾ��d?�.�]��	yg?���ygC��'����~�L��4�`l�FSdT{Fb��N� ��S�����C�!���t�E����;�1J���S�q��K2g�}��S���O����Ͻ�ڢh޼�n�\錻��*<G@z��w��#�r"�y9�W�����=*y�^�������s�����l�;�q;�����;�thGtb����$��q���捓q(k�2�q��0'��$�?Do�B�͗u���TE�ѨvK��,���+�|[;_���:"���(�w>��|��Nn�<ov��2�h<3�)4n��qk�4�DCAQ�ܚ�f#z�q��DH ���{�bٺ��m�,���7�]��V�Ǜo���?�����Ҕ��i���h6~$.X�?�Z��g��_��֭E��<l�)F����^��c'ʹ��M=����k�ڊz���-��z�D�z�Tnn��ɷ���+�5\&
t�%6�i
��^k�
؇��M� :�c��;Q�[��/�ex�	p�i�3غe;�W�ǖ�%(�b.�o|k�w�"{c�G?r�W���d,}�z�3�k�J�>�Rz+(�}���gbf�Q�w�@�_7���A*�c8�3UA����:�$����f#����7��u�lGM������)����Q����9s>ҿ�G� �&�z]�u�y���������GWd���<�D0r��yY���݇؁�P�Xg����3��b8�K�~�$��O|��G�h�/�jN-QRk�ȳ��m�ѡ��lO�7K�J�j�f�f�o��cٸ�[!�N��c�5gP��|�?�]b��//���iܐ�^�S~y��1���D���,�`��Hª��`�շ�~1SVv��\v��b_-�m�3�k��Q��'X8[�b�~0T}Q�����՜�L�Q�k�Z�[*K�K��<��W�=���F #�?v?����Tm��v�
�(�9E��!�-	vl���me����H�b��������-�C�u�4JV�w�	<Y����,I^�_0C��$`�� ls?����={[�4;_�n�0���R?3g!�W#���1`�����=�{z�.H��:�k\"��=�u��[ R]XN�@>b��ym OG���;��OGE9���<E6�	��\�V�ӹ�ǪOp�7�B�n�7�ai�Xd�v�z�y��7�ut�g�����7�p��1�����V����]�s]|1�E����~�8~�_{'�
��z�]V�_:C*�u���B��� �ZW�����.=�ɌN��@<���h+g�������f������?�^��!�Ƚ~�<� f=�<~��>|q��X�%�_���O#� D@���.��0�w$�ZԸ$�!�/J�9���h_5[w���şF݅�Kכh�xn�0��сl�?x��3�$�|���#c�et�����,�{�m��C�LW��
�`y��/���u��'O�q\����m���^=���-l�,�,l��:�#��!�څet��#Wuļ��p�#���lc�}A����<��9�υ=}֒B�]���GA�����rUAb/��g3<C�k�\���~ȳ:K[�����X�o�I��F��Մt#��&�ܔ��9Ȝ��v���Oj8�Nv�G]� ���dwEAN��NyǢ�?ќ�;�����(�Ԁnx��8�x�#�l��֬�����S����w{�ݾqw�c�]���w<��a"{:��aW<��wv�̎ q���	���0��v�<��Oz�����ȟ��/xE��[�¾z+����������JO<I�t;�T�o�g*m<	GU�0�%��5x�e����J?T���B�D�WF/�-�u6k����<��J�h��Jȋ��-/8Z5�mx�ؐW�p���܆�z���"Z�/o3%y��f�v�������Ǟ��OLŴ�>ƪi3��d96�KGnV&
�~}:�W�������OH~�sL��E|Mc>���M�ކI��� g)��s�ڶ?��L�(dt����@�}a	�9��t4� {j��Y�AiyZ�'��K�X��
bP2�Vߐk�u�L��]�<cP���
�d�r�I/A�?!��G�❈d�8���^��2��k��%�����E��b�_���o����z҃f��'��J4��G�0�1Ht�����D7��m�#��攁<ExՄuM�H�҄�X���}F#��W�����z�]�p�2ۅ`K���Ξ*U$��d]F�x�7�q̭~�U�m��6� �n��ug�OUئ�:�#y7<���	�J�S.L"d���zJ{ڝbvNk�&AO���>Xα�A���1X4z�5]����Ǧ\�gP��lyYq(���l���yʏ'��憴�X������ʓ�2�'V�E�n��O�PS=�^v��b_-�U�����c�(~�]�&�mw�6�Aѻ|�B�͚���(�~�����T��/ֹ�<B�O=�M�Ի���f������)�V��8l��)Ǜ���%Мy����mA�۟a}�P����������M��kZym�ˤ����,9�$o0Q<A��|�R4�m
�ެ8�O9�������GQ�?;:�w��z���ٗܰ��8�5¤vYK�N�re�NeP�\��L[��Fs����a�����y6����t�ׂ�}{�֋]>��"���ܛ�7K�:.��K��E�Sֲ/'�<�=�cOs �IzL۠��˕ƅ�+���" \���͊�	�f�n�{�f��b�v��_�<^�iNl܎���<�>X@9�}W����ޘ��9�>X���ʮ8J�]\�/���ª�p|�_���{����&`ه��y�6�_Bu��׾��I�s��$&lR�uY<J{}���,/�%⽑�ph�R*�F햭�~��x."S�����ex�x������k.^x��i]�˴�/���n_f��������ǾD`����o��򙳁����b��a5r'���!���.�x�5/������]v�D�I&e�)�1������B��Vl��0��X�<B�2'��D:�˂�XX��U�\�$�Y�~�&�ʆ>��������||�5(GqP;j;c���1{��Z7^�f��D��=u]�QM���J������1�0��� �_��v��� ���?^t
���ј�0s�~u�H�4>���������p�?.��Wu�����<ͼ�D	?�A%��jͽ?@��!� ��x���c0�:����"=����N&߫��c�{�����d�譯�5�h��A���/n`'y��#�tw�&� �AɌw��V
������U�8�! :�aoG�vӣ����ѮK��������#T�G]c��~(�2��3�Γ�<j����5�g�gkδ�s���.xlO�Dm�����O�����澧0�ڛ�q��l�x�7h>�=�q�|����G�"�����Gx�����1�p1Ӄ�bn�h��1�E{�ƫ�����
c�/!h�w
�0�J6�!�;xc�sϣ�7��x&�^���ɢmȆ<����N�Ⱥ�s��h��ʴL3����}����XA~��,ĳ�k�V���ϿG��3���H,��G�4�h�tG�[��b{�h�%\�����8 �C�;9�����Ů���IG)�	�h����G-�V�U=ضZ��
y��'	O���f�M��is�Ŏe�XM�u�v3�]CQ5���c4��D ���1zzTNA�l��uڅ-Z4�I'd�o�}g**M]��l[w���S,�bX��W�aNz
K��N�fa��N0�7�L�6�KH�#�wT8k�X�K0r�c���c���hH��c�B��
�f�;�&p68'��J_�h|)��y.��g�P�4��y�ԅ��ݶ:�'����C'c��3M$��e�����:�I�|�8�zi~}��Â<�]����M�WB�)��ϣ�� ֹ"�3����y���:��Т���Z/���Q��	'O�n�Ā� O�k���ľC�~�Sl���"L��P��sJ�q�y�S��vڔ�mR��Иe������~!�@^���Q�h-8|Q�D	��˶Gr��p
�Vl�����Է?vҙ��%�D���ϊ�`aGs�66h^l6�g�S0�����H��Gj@$ք����b��U8Vy�+�P�h��c&O����͞J�%��x�Ґ]kґ<d
V�$a�UH��P~��Y+	�&1��k]CLo���O��H� o���-rv�J3z_�\��W ����v�>d�����N�C3�}i�6��zb��+���`�ڒ�;� ��_a�l�{ '<+�`a�H,��#�Ǌ���	2]AS����j�������m
N��7A��18��͇���U���x�`�w#&��ׅ�a��&�,I�Ϗ��W^�g�z�q�ȝ�肇/�g9�_b�x�c��^E��\�@�s�?:�A���~�-$�r;r��	($wp!��^��c�����ax�}�i�P<��_\�������W,N{D��)Ȭɫ��5����n�6�;�s3�V��<��;�%�ݕt��q�-
I�!��\jw�� V��<:�[� O�k�yΝ���A�#$���Q(��}�1���r��t	3iT��N�fy5�8Ju�Pu�9��(�"z����m=���^����镎x�����g<�tD|}�èX�8x��3��ѧ�)���f�l�H�/�������/t� �y��=�B6hg>�+ל����:��~x����+;�)�0L��욽 ʴ]�4������eGz��0��,�mW������q�OO[
z��/v*�I��2oTu&����И)Ŋ�Q����$�pK�J�h<��S�t�ή�@�!�D�8@yGid�	y�ʚs��Y�U+�ɩf��������,����q}0�� �ڭ/~f��q��"�X�Ne�O�9#o����Xǎ��o��	�X�r���;p����O``֐Qԇ�VI�bb~����7j
6�Ec%��GA�/`�N븴vKP���%6��x�)ۼ6����DT�N7Ӝ���wW�ِ'�����łi��?���aQx,VttF�2���4%�1���¶���K؏E�����C�Y����Pt�]�u=�晗XQ�΁<���.ۓ��%�Yӵ-��� O@�u�J�F�N�8���ߝ��>8xy0*x?��L��#���D��t��`O�zm�?J聮��e��2`}�`���+ϩ?Ua�j�iC��_��g��]��M��^�� ��f:Hm#y�C�;�:(�^0ֳ�_���!�0�X�J�����g���:�5a�3�}� d�ě]��A@[ȣC���z�U�f]�Z:oi�ܕyn�@L�^(�~.-�)S�s�b�Q�z:����8\���^F&�=4�e�Q[��y�t^-�+�5y'��Mɇm��U"d���H���bU@�?�	�e��'-��i�Q)R섾�M�j�űc�L�2�ϑ>�Nh�I���N�.�<���6�R44��4&�Կ�����M^�{>!��j��ّ��Y�L䶐��ڐ�{�=��@+N��r횾3zL���ށ� ����:��}g�.��XA�j� S_�(t�zY4�YnZ3���h��8g]w7�'g��k��PK'L�_�����ح������R�{R=z�S�Z@���]��zKg�jg�y�騮$8��.�>P��%l��(3];��(l^�ܤN�i���S�k({�"��w0'd(~����eRdq%�P����]���HkW�낃�h���\�wt���XN�&r R"�c��I���;���_�_B��F���c�;�6A�*���ʝ��f�Q���v����p�C'�B`z�v�ɸA�剷q(�8����ٸ��6���?��C&�Y:�����G��^�d�������^��w���sϣX��Wؾx9��w���ye��?�����'��^x�5����>K����_��$�bШiZ���|P�5МhaC�v���6�g�_����D�yG���^X��4��9�&�'����� ����	�6��!���y#�������TH���J8��"���k������Q7B�k�un-���������kSJ�z~^���<u
F)���<7RY}rYg���ϐX_p�Ň�}1{�]���l�4$��y�||~��x,8ʜi�T;w�́�+)��+����<�NGG�z�>��S�ʁ�ʋTLO��O�R���n�����ʬ@�f4}1{ny��z�%N�x��;$�=���r@l#�c����w����b�{�T>����K�~.��S�cA�"z��*���-���{c���L�<!�#��W�hZ]�WE�t�����y��ZЯȊ��&��4�(�w7܆��i����2?(K�aQh�֭���J��o��n �0������(�'|m`=gy&!eЍ8�b�b�im��"y�m��Z[a��[�7c�z��G\��7L�"� �kV����eD��$�.�(��Hp`:�"����Twh���/[IJ�2��2r��?}�	J��ހ��˴�O0�6̹����P�"����NQ[�;�}�ɉFN�d���B+l��iJԖ�l������K
�y����:m�z����v�&�SH)��������X�45�Vb ��8Q�C`�ݒ)A���͏��,p�%ZA��w��j�T���{��h�T�8'��(W��l��zI��~4����zZ[%��V2�:���T�ơ�P��lm@i5n�]�|m.}�ĄNޛA�e ҺD G	�y_�]O������t�e*E������
:��k��پ1�C�5��p̼�NZ��rY���Ko���s�K�W�}76������'���dN�(v���Bg�����-<�γ]�r�d���tm.��f�H�䥅>�9� �O�1��Nlط�.�r�	�����Q��(��}���Qt^y<�,S�1�}&��ӱ���Y�<:e�~� �d��S��R�-��-Ƿ?҇߁�Kֶ���i��L;A�-fL6Y�DV�=���/��n��=Q�!%��U!�QD��Lgb�]����ثl�A�6�h�Vk�2=�id%�Ώ��1�c�bk���L�ޟ�lQ��dv�N����&Is&����l�E���է�Y%gVdO˔1=���Ʉ�n�XJ�[�8���Hԍ����ٺ���ͥ_�	U��Z�֗�)j |~��y~a�Hv����Z�f��Q�ǝ�p�����pȡ#������y~HO{{A���_G΁�C���[�T%NA����?��j��IorB|d�E�.x䪫h�]�8��I�x<����������܏f�zm1�#ki#��m��ei�6k1�~���~�Ͼ�ߞ~��xٟ��i�q4c#mP9PA�&������_�S�C����m�P������`_ӉS��	s��&�n��I��������>���cC�sj���|RG�M��hߴ���Ϳ�Z6^����p윉������5l#:�B��g������/Aު��0��K}�1<;d��b��-��g� o';���VOI�)'�I)�J5�I� 4�Y����S��#NC*�ZBSe`<V;�೫1�JG<A%��s,�rM��=�a��/a��d4l��B�6�o/�v���]M�ͯ?�L�sqǫ|���h���Ae*)�qV��!	�e��8�,�6�i[��H���?�2��:��z�*��:���+�4��Nn�!�UpOt��B�!B\[9B��ǃ����g��yTto����W瞄��qx:��Ј�����6hJϊ�hp�Bީӭ���j�<��3�>����������`NX,ևE"-2񋛷پ��`-�'�|�enȻ2 ��57�4z�ܴNT��f�C�{2�hR������_�<��1����JB:˼�o���n7�g ��Wp���A^qG�р�@����Z��Ģ$s��_*�-v��_Y�9�~��_U��/�' $�3i���S��aԎ<����N��Xl�/�ؖ�<�3�vI7�j6�W�p�Dl[���������,,��L��~�&�m�S�Ӯ�"aI)��d3�����L����a�NĪW�C�I��F��7T�#,[�C�t��HwL��.����Pg�NR�I�QTVmlEa	)�T�~3X��D��Y���:y����Y(_�KMoC^���1�k �9D�i�t��.<A^;�E O�.��ە�Ȥ^���q�o~�xv�_�Afʤ˔ɾ����ˬr	�Nmۍ����&�^��IP#�v�B	ǣy��k�xک_�%k��Y4Q�p���6�~Aȳ7Z�ux y��O����:[���(������9(�8�vt.��V�x;�V��$��@o���B!��?���Χ��ۖ�`W�^�*�0�'�ԎZEM�KcQc��e��c�y��K�����&��Z`t�C V��͢�^�:L'h*��#��Pl�-�*Ꮠ��o^Hl>��-��x	��@m�^6�I�������2��@i��n�����i�V���xJ����'��k��Сf�=	��*�,��-�����ǐ��GOb�G����X��u��"�ŵ�XC���NA����t�j������G��G��V��{"�6za\?����4��?�<9�����p4r"�����!�h1�N�:AΨ
�7�ׯ�;♿�ǃ�;�I:�ϹF�e���1c�A�k���"�կP>;5�;Ѽ� s� �w�TF'{� %���24nڊ��|���^�
�S^��w�W��ڱ7���{�Ef����x���0�
'��zڢ � ��3��2�c�l�sQ4OӲ!8��Sl�ӎ��]����<��t*�s=���{`pv���?��~.�s���@����C�N��膴�(� ���q�d[9�!��kyun�9�P#
]�:S<­S0<	I�Q8��ʀ�Ř�$G�b����Wu�#�(T�*��닏�����7a��zn2�e�
ky:2��	k>��>�󞝊�����膻"�qgD^63�>��>�y��.w+)��<���	������}�B�*j���4���K�_y��sBOv�o�W{�<�൅����Α}�4�x�S ���1�ٱ8���� /�!O��<��� %��hp��j�;�pW�@%HEp�d�A��5�gA���Vݽߍ�C�P��̘8����Wn����4xJh*�r�36\Ie��ǂ��O���-�e��� y�b��[���4�\;3�L���� O/r�����E���]�R�mQ9R2,�:����ؗ�>�Ĝ��L���X&���q�:3A��N5�y��y:Մ�.d�Yȓ�f�$jK��=B� ݆<;G��O���A�׶����墐��SՓDu�:�%,h�f�e�f�u�o��^����g!OI�UΣ�֚���(�Q"�;k��� �^Wiꆯχ�,� �cy��c�_"��9�뭴6�?��v�]�Rmi-�5ț�=��%�����t!УS�6�iW��]�)�d���Wz �
~���!ݐ<b2��� �L��ec�]���i[���:�Ի��M��l�nf��f�%L���:Uʓw!�[|�U��(��1��)f��ky�΃<���GP[]�:k@���	A�QzU������K���rw�<ll�m"��A�6^�S�9GG1y�b�oo���ۓ��1[�����@�ʩK�h�Ɔ:�tT�ǎVbݻ�a���Q�4���̚�Ml����s+��g]��nA澊�	�6��h�6���y�z!s�M�;���E�����q�ҥo�?��9E�[w��]���:uA{�%�-�Ѱ�'`-��X���|}�)���G�t����x�,����ݰ��~�$�?�lLIw9�<y��@^U��(r��Cݼ4�'�1�b�"��h�'�d�+�;P�m���ʰ	������������f�  �i�e��]��,�R��g�"�_,����{�I�<l ~�y-���6<�
�~���A���pjV*j��B��Q��(y�=�>��9�c���n��I@�����0(z��s^`�z�N��jf�����i3���f� ������wE�s�.�]���jDG�v�Ύ�)u���)T�i�;8!-�6�C��%���'#So ���3 3��b��R��
��V�ų!o�k�����*�]=&M�j�VbM݆�W$��"��*v����8��@�_#(	G�����]�E��u�śN��� ��C4���_GOA��ob��ѐ�grv�i�}�~C�Yy���Y3�}�,T���3}��`x"� U�3���o�v�#X>�v��k�$�σ]��0=���/S���(�cY	�'ؠUT*�#5-{aȳ@�@�"�h��x��9H�/�+g���ڳ��ǃ�a�Lך�ej#^�C�"�Uu��:>7;n��B~�����\�	_;*��k��^QID�"���cWw���o��
�F�-���Y�<Ev9�4҄<��������a=��k.���7�($ ���כnƬ���"�`3��@ކı8���}j�0���Va��'[�*O���)z�5~��I3��3�-(���:Y�k=�x�|�(�� oK���{��ʑue�c��T:�8Zv���	0�B��i�(JgĪ#���q�/�d��B�a]`�K��kX!��TF/�ɮHZ.A���J蜿���ǆ�	,W�YOy�t�wz��·�L�g�/�eO�M0�W�Ȃ<3xs�Qu�GFN��!oϛ���r�C6�B�'� �JObC�������;za�[y�+��I]�뮽�<����-��=��^v=�_DB������⛧"é�;����M.MG9�(&$\�^�|�3��Km���?���{��D�:e!��ϱ!|8
�4m��.�#:Ҳ���Y���Z��A���L���"<P���"�p������A�E9��L��L9*,��ig��sJc�֭��(�Qy� 6�\���öc�O�S$QK$J��°���,�g�G�I��݈�<�F��s /'0�w�<�_����?�bf�2G�Eg����L}1��3�pl.d_��j-^VXw�k�+�OA�)-��� �\�GP��GX:i^ݰ�*o��`���@^AgG�p�`����%�����Gй������=�폾��Q�pƱ�8XY8�hOt�B9@�g6"�hws���;�U�����ov��.�dB�G���/#�㇄����x|�4�t�����ȑ�"l>������|����B��1's��3W8�8b^;lu�Bc`7��
n���N�� O�T�8V�bn1��h>Fi��.��C��$g�Z��G�G��<�e?M�f��|W�w�rҿ���F�ص���J�p��f�*�#���V^�Ҩ�t�n*)�Ҭ��|�|z{�o�$��#q�+�p�?h?��CZl��P7;"za�Wާ����2�B~�7
O�߾�A�o�n�-�:��4
�yŏ|������o� �7 ��@v9����sP��r�{�kTL�ŷ>��a����1�������r?�/���ߝ�I;?��wǁ�&�w�1�0U����"����Pw�ذ��%Z�g��~6�ignE� f=Wx׳;R���ɰظ,���FM�6�D%є���՝�ѓ�8Q�iZ�]��%VDJ�������i�����`�['G�bVbẅ��R���!ǁ��Y40���4�N�(�A��j�����~7���Ts�1��T�m0m�M��H�G�������Kfݠ�n
�(��bC�V*F{���o
�F!+a4��:����VA�/�^����`���8��0�}3����{��Is���+�x_{�[�Y�`�hQ�9��Q�}6�GƳ/'���+�N�g�{�k��/y���?;ƣ�K0��%Z|����������vBJl��%E�*�kZ/����,�@���Q����KvEb_�K|BK!o���m��m�Q4E�to�+�9~��hc���r�:�US��}L$o���&Z�w�����}�R�j�L�V�c�ߚ��l�D�Ϸ�\M��WBf{���v:��ɬ�[D%��rg3F�D�@�{0k�����t*�M�.v��6���M�t��^�P���I�V�U[YLbum��J%A^NE���g ���;���<:�9�Q��w����ٗ��v�
�l��蠁:�Β��4�U{���ؘ8�fN�(���9�:�|�[��rTwZ��M�t�@s���{����B� ��k oϺ��z�m�h��u��]ػo7v����8����āfm���*���+P�9���_��)-P'��Y�l O�]y�J�<�f����C�B�شן�l�ۿ.�߁�>t��ByaW3U�����_��C��M�3;i	Y�EY�@�±���5���.�X7�[�
ym����.u�7��+��6#���ܿ?R�{`9�b!!E'(��@�*�ⵄ��!���W��E##l 6�Ī�aH�S����<:�[z�1�qڡ7m`T+�ղ�װ�N���4u��^h��-���ܿ~��x�'���9����G]C�,?�1/u���x�5�:����7�c�:��u�X��e�.?ñ����x�2w|�?]M�����	�LǛY�:3�6�`��ϩ��Oχ�&�H49��w"�M�q8�NXt&̹����m��ݵ��s��X[���E�X�R��u.�i��L!X��E�GOTcO�v���3��?���k+x��/܂�ۍ0��;�+s�vV�N��҉lq��3�����i^[<�������8�>!��&�x4G�NR���/:�c���X'�.E�V�%h��>t��G�������`Z��1g��X<�!,�0�y 3�ފ�zO�7!}�#=��I՟r �N��5O�Q']<~U���0�"�/	�>�8FϠ�
D�`j�u�d��6Y�Yȓ���o��C��}T���z�����1O��C��u�귅<����R�ʏWS���@��NW`E��3L��`����݌�_�5�t��������Ȝ8	�#ƚ�:S�/5i�Բ�v��m4���M]��wNDf�Iؿ,����Y�g@πɟ����y�d��7F�Ċ��ú�4C��6<E�H�A^�c�y���s�>�/%�^����u&��#CFc��b�6����z>*�|�ֆ���g�����y��w%�#�������u��v��E�3xs)��X�� ��!�*�t&Jɡ��|=
��лO���Ǚ�,�"f����Y(n������w��k:�m�i�݅<�k�{$tj�y�K�A�"y��<%�^1�:�.� O�_�*��҂=�_]��g�<Mզw��7�Ge��x�;����eW�:��f~D"��p'�N����,���6��`��� ��Ҭ����}�GdG�B�w�9-g�B9�v��N.yZ'��!91�=#��!;v��%p��&lG��>к��J�r�����C���<����}��pe�.WY,�St��ٞ�����<�n��3 )��X��g6$YǇ�A��{�mE�Y��Ge��/��<�[QQ�mʰgaoU&�N��~�fgmQ��w2��8Ec�5�27y��k�<E��ZB�_���"���w���y�~���X����"Ӎ����Iw���T;k����q�J��
��v�.f�_M�x)��:��j���Xkm}z�>����ݶ(�C����&j�� ��0���dї��c]������錐tT�cM��|�k�Y�����5�z	�w!��Wq,r"��D�CM�j��I��a:��q�Pj��98����#�'ځS�<�1�d'W<Վ���j#
�<O��"�N�x�}��+��2K���/�����?ұS$5�1ǃc��~�2��(�Zz�v�.Z8</yg�{θ�Ygن�Dc@<"�tm��B^to���G�E���-^�
�x����W�I���`�QT<��K���O����^�1����<q�?� ��[F������{�C+���<)'k}�6�6�a�����ʑlu��n�X���Q��F�a�#��	�	Iġ�D{J����{W9���	G����	�N�x��OҨ=I�Yv�Y��_���/���씹��^� <���:]刅���ޑ��aEk���TR�U9D9De���!h��q��{���%J%#�����>F�|�K(�.��(�v�y%`�s4����
y���AIXQ;E�8�ϴ0�f��,��T�Y����d���R���O��%�Gbi�aHe�ө�ͧ$Ú��Ƃ�]=(�v��ӫ�.��$d���G�yWOA~pl��O<�E�=����~y�Fl���y&Eǅ �I�[e�����|z��+�"�jCދ�'a���zE:�8x7�.�3Ti%,ȳv?J�]�g���{�2n���T��Na��k�@_�y���v�;�:��t�iQG�s!OPGP���=��Ț�K���ƜbБ0����ݍFe��t5���S}�nZ/=m}�a����^2�NB^,6{�c���Y�eÝ�i��&O�ݵ��]�<yt$�vƂ<EN$���'�B^F+s[�3ɑ)�	xz�﮼��,�_���a�X{��ʦ-n���]*�y��BY�엦�j�p�YX{56{'`K;O� ]��5Ɗ�7nyJ1�i�t��\o:l�<�z!�+��̊��O} �0����}�!�	�v�l�;yVBd����,d����H����D>
������)T�_�Tu��jWo�[��y~��0����ᷡta2ʔd�6F��mOr>��w�<n�[��]��m�z�2�V,q�D���pI�>t1�z��+]�ʛNkP��<�!ϤO�ZA���h����QSpPKc�<���y�_� ���KS���M�q�˾Ŷbۭ���=�����hsY2��*~��5�!���Y$5��@���ĥQ}������q�s�u.t�h��[��gv�*� O�!�6^��Z'��F��t�D��3������6�џ���K���C(z�MTF\����sQ8B��6j�^��6�ℓ?�u��I��z�mެ	J@S�a���m��(�E&���̢������z�#��ԓ����|pYW���f��kSL9b3�}�'
aI�^�7a�<r�����DӪ�5�JgE��L�������v�6�F�1(�
�?��N�T�)�g��q�G���;�
y:�liXw�[�ªË\�l��#yZ�z��Q3 ���ŮŘ����ʋ���T,2s\�p0<�\�̀��)pkyT@���ᮌ��mTV:d[p��-��No?�#�����M{� ��Y�G`4��Ⱦ8�[<���]����_x���up�S���/����N�\yϱ���	������%�陎�x�]'<Bo��vx�J_�����w���Hh"�b��|QC�_���[�w�}v!���6��������@Ok�9z�Nm �)��H�y�H�\�������a��U)���3��M���^���C��[���c�������sj/�IV���Z ~>��c)rN��s O���$�TY��5�<���݅���Ha��z�a,|�i,����Z��x<��ܷO����@^�H�|&��"R�m�.��kJD��O#�X�Ƈ���gXOe��)�����eN��t���'ȲD�eE��Py�8�M����E�y���[��GDo&ڴ@�"�,ț�;�+%(m�̘c쩌�<-��m�b�vJj��6:��%�܎ƼR֗�
**K 0e� ��/��oI�ם>�vV/�tI
�܁�J��y��U�g�i�GǄ-��y�S>ױt��!J?�M}��HȻ���XkǱy�	�ѥ.�1�j�텯1ǻ?r<䭧n�!O	}mȳ%���y�A�K.s�N�H�ǜPB��)X0�>익�xX�^.p��6���^K$φ������m`v����6�Տ ��H��G�S}��iN�(�
Dixև��������枺�=�)ю[A� OS��:�t��6i�|3�F�9�h����m�&��J:�&�!�L��R�)�\�KV��������쉔��a�f�v��k��s O�H^�U6���o�^lY����݆�NQ�;�f3�J��S2����=Ae�w82����l�S�hCH�JA�@䎹�J��K}Z���ں��(�֥�9Ո]�V#��$��ņ�!���[�Ny=����c�h�D�.N}K��&�q�F*�l�K�I<\��4��8���ݏ��՜���fb����fw�j�mY�D0v#乳L�H�!�����7����p�s;�!�'i�=LB���c��߬{�j���X�K��$��Op<~2N��k�� 'T{�bmܴ$�ڱ����z�8u�f�� �5�Ơ10����큣��P��,ڕ4�H�O�#�S�$!/0~(�AUXNGtG�_$�-�@\}	q~8C��Ⱥjp�1�ʞ�XP9�qBiS�z3;k[ φ<=��������I/��j���ʉg��E"y�=�-��4A�TKF�/����_�hj���GDy�.k���[�1�O��k�b�/�b�=�Ữ�(I0k�t^b�Ov�v���kʖ�z+^�WƊ1Ӹ$�rv�=�1����RƆ)������;�wuj�^���(�s�~�(����!����|��iZd+Z����ɻ�|�6�˄��.w������[�^S���/�u�>#��L㢃ܷQ����>@DO4�F��x��Q#У�=�u&�ٰ��\ص��]�Aۈ"}U4�=��U��v���N]��n��L���>Z|�HZĶ������19���"�%�H�d /3 �D�ys�)CGb���H��6�c���ms�A���Yї�N�;A�A�rd�K��cc��8�<��d�5�5�'h�!�Rj{��{�y3&݃L|*�֒GE�k/�)��k:���xAv�δfI�o��+u�5�fJ���D>
�F ��XTL���ěT%�ԧD�i+����yz�u��~�=�*�zy�1"��U�L�g��R$����L��ޜ�����&I	��D�:�X���	yGO�J�X��ϭv�˧�7ѷ�������nע����>V�6R�NP'���l�M��Q9��xv_K��Kq���Q7�v}.�
��P��?�<�V��)Ysm�V�d[v� l���h'��D~8fTޢ)����xj�B����T�1�u�#���%!y䭨_�q��4;�yW���I���q��\�LP��}�#�=���9:-ZO��FA�$��`�`k�l����ɬO�[B�v)a?u�$̻�l�y>+���/*��l��T�j{A�޷BJ�(�U7l���4�`E�s�悒+���49N�&⣼j)ԥ:�l���Y��9���l���p������B`��b�=��(� :@ſ����~V%�BZ�`ld_)���B�6K����-%,�up�<�)��ʶ��Y��V�,�	F�_,V��p�M"fٙ����$�������u�f�MX�ov���ò���� �h�4:�?�]���<����r���Q��W�g46Q��'�0f(�&?���B�Xcf����.�A�W�(�e9�'݌"�J^�Ps�v����j�J�;����^�F{�)]-QT3e�>f�J
AfAto}?���6ҫf�ٝ�B�����'Oc�糐9���ay�@,�Ӭ��>QБo؏��㱞�掮�����M��;��:��]����^X��5=�!��Z�/��3�����Qly�sK��&�~�r��Q� s�26��1��P�s ����S_�RC�����$ ��9\A�j5����7G��H��`����8�M!=���!�q��w: 
�d�f�P�d�;[��D�t'�:W�Vi�>hbWJ=ڀgC��� ���5�Q��4��9��Sn��� ��[[��Oy��ݬ�K�w�#L��1=�o�*V�����Z�`?y�$�>�D��,�;P�=[���O���b��/c��7c�Wv�r���bzF%�,[�awP1����w/�>��>�P��kQ��=� �,��3v�2�p�^OQ���R���#�	��3O>�������k�Yyq�Ow��O�n�@�����}��-�9�������v�YT:�<H�,�W�Y�RJ/�0�T˲��OQq��ï��jv"��-��1RՉ�F�I��4={̉@G��#����w��W���W�Ȳ��Ԉ��]���й�g({XYC��>%��,�B���`{M�*_�̑�#/�'��.����z�`�ȱ�?|��ߔ�wGds�o�'U�6�!���U�(Y� g�S/����+3�i�XSǼ�1��Y`�VY��Ӽ���'���'�;��� �u/<��kJV[��BD�Y������g�'VDGBk����6�@:ǡ��580}+��f����������k�~�� �<��9����qD��@S�4yo�`Xu��)�(�,�c]d3�
<f`J;?/y���+���oy��@��h�B����#Ǭ��P�N0XG�Yt�d�o�d
�Y���ιXN#�R,҂��WM�V䏺Y�b�m��*ݰՁa�r�����/�^	봈�`#��2����;�"ſ[�eY����$�~W�s/�_�Jt���7��b����&�nC7�$A�g��;�V�s3��]���+��n��Xt���={�_���zS�ڐW��H���I�q���eh�I�۱�x�_��PY��N�XW�R@G�JWB���{�0m�{�����J�R�{��l����1Aޮ��Q��i}���XGG@I���37;�����~��'��f:{c��]]�f�W�E���V���(}�HB���VdNk��Y�.5��5;͋ �d�~�}�){h�>�.N�7CnF�g6Љ�!O��)b6�m����;y�C���+��%{�"Dl���������!�t��&ۂ�X-c��Qp�q��B�c��+�?�u�y����,ܟ���X�լ����J:�ȝ"g�~�`Mqk�6��ߤ��-��o�6�<e@��UF�S]�q�K�מF�W��5	Q	rs��VR/�#)At6�Y6!/��`sGgڷέ�w¡+�9�"���aA�qj�(�����0�V/���\���8	�>�9��݌fB�q�TQoc_�=��9����BbL�`e����S�'�Z�3]��:��Y&��U�������~�@}�ȝ-6�ـg�`g�)�]��-��ِ��4�D�g��M��@h�wWDOiSyڢ�������%�[�rdX��(ֆ<u�׻��	�������c�W����i�V��{k�|�1���nLy��ANP,���+({}��mg��IE�����31��^�
���滄�}^Q&�ge���`��n�Nk+;��CRDo�G0�y�=�H)�̓���{x�:R:I�=��nhJD�1�7�z�)� a�hpTQj���!�/��������Q��c.���Ý��<�O��������w�{6�〖��j+��)}��D���>M�瀫��*�Z?z�x�����/һ�_.��X8*�p���6�i��3J�{
ǚ���(.��� ?��Y)��< ���#��"�i�N4|�(Q"S�|*!;T�2X�H�v��(x'��fE�3����L?�L6�ّ ]��4�y�����ȍ���8,��A�}�i:��@�Im�o��5u��,�`�D�Z Ke*L8
{M�A�PiY�h�݅Du�G�G�������_�o|f"�;�>�����~�N��΋��y�Z��i%=>�{�����i��%�6ܷ��ʵ��c���h��^�Z�犨	��c�L�����-��[!�.+�t�s�DY6��̥��/yZ��d�W$�pԽ�u�7N�fحT���:P�s3��CA`1�F΢"�r�\���K�xȢ���� �A��J	Z�d*�M�.p���8��׾"��2��1�2��k��;�X���vJ/s�R8���%{G`����蚻Q1��רVj�ns�W�����z�s����ݱ��UgM���)[:(�����p���ԑ��G����1��#�
��	.CPvˋ��)dZi�ο���ځ��ZD��<l�E+���ߌ�S_Ar�@p0Ҩw7��y���D��ɶ]�쁥�<ǥ��f1�r7�VR���EF0��1��u�2T�4;{uF�N�P?A�|z<᳒4�.)��sJ�z������H�o�=0���LW�<��|��z�Xo��ΠC��+�D�2C�!��p,�}��̖�f�?��'m����Rd��H��r��;����J�����F�f�E��d8� �)��aX�b 0�z.�c'�9˻��v����������F.ui��3*�z2",țþ�k`��őӒ������r�J;Y�'�����NnHu�6g�
�2����o�ofؑΎ��x�����g>���� ��8�mv��ӵ���Z�clדd����(ۭscu��I�]jj�;uʖ	��f��hKtEMw��C��>�V�3�:��~~)i������@V4��o�{5�˱�٦�m��`[�ZSǂ�C���C���/\��U__o O�H��	���b��6�-��C|u�͘5tr����$�Xa�z�x�
�J��R�TRyJ��?VFX	=�Y���l8M��rߩ�v0I[ȓ�٠�i�͞4�-^4��
���b�g �{���;Ҝ�]p�B���e�N��C��|��R3׭E��HA`\U�y�cy���G��P�:�8�<u޹�g��� O@���D���6�U;i����y��ov���x%j$
W�v�Q0�A+��T�ni�Z�N��ūj��&��/؆�c&�UFW�����3�Z�5�,�U�ncGWle�ۑ<x�f��3�.�w����C���ԍ�,�<+�q�Z(EM*�6��VyM�*1��'�= k�@�<�82^x�dd�z	E�4���6XX@eA��R� v	6��6;��;q�O��4�����Z��r)�S
��S�ā��2SN�]X7E�����.Z[4ulI��/���շ=�DS��6	n�v�=�v����l}��3^�k���zy���䙲)�����<M�kݗۦ:E�C�kt�ϩfӖ�:0Չ"���ڰ�p-�Y�S��lG��������-'�mc ��U��ԏJ8��h�S1k���i�H�G�Pe��&����e�,��H��<�ş��j������g���]����7�σ<�4��N�O�s�����5=�c��[�������Ur11���R\�W����~�u�q�;�l�*�qЩm��v���ơE����i�����5k��@o�0c� p�Lz��7^����&�V%���5k��ڷ��U\���=�ա�Y/!�<w�sv7��jg/,vp��^�C��-������e��<TA�Z�Pl醜�7�Pr�����Z�:>�=҆�l�3�V��C풦���e��S��'����)�R�(w��Ξ�NGT�Q�E�^XB@�Qa�n�&'�ҁi�u!/5�'2��m'�f���S�y��w~��1����I�3R�^p����n��z�pA3Q4�H���sc��9��T�F��U=�Fټ�#��<�l��qt���4� /;l��aqP"���cqp$ۈNǣ��L���:ڣ���5���FNt� /��Ӥ\�����~Wc����@V���U��x��C��Z��(ȋm�<넬�!OS�u�3� M�v�v��u��Z�)�P�cŨ���t��xAύ�7��	�g:������ OS�����J[��h��a˲��8�/if�$Z�w�������ar�Ѿi#��o$?I���yM�����k lO�@�^zp�a��=�m���w���b�����06�E�TD"�������;M.���I�C�s8�7�����b�o��V��$ڕ[N����"᭐�G�� ���V�R*zd�lУ�,��3
�Tr�>�h��3�=M��q�Ht�Z��?{�D�p�����U��ɜ�Q7P	T��ᨓ3���}�`cM�Z�g�	�/9�X" �m�t�1v��-��S�!�$=8��3g�R))���(��7�F�x9!�A9��dN����y۩Y���H�up��H��o���7�����鲴�x3�6�V�pt�Z��.�z����2B�vXA��@�E5E�ͥ���f<`u5�c��g!�5��[!�
�Ek�w��x���Y�������KXH%,���<�[G�)�d�{��k5]��_�'��LeP�1��x5�|;�R"y�?�Ce�!����ệ�"㑩X���.��L���"�2��mT>,��� �|�K��q��)��RDS���X���ƈ>�w�R6�&�Թ!��I�&�Bh�N�e�"��k;���Z3��2k�]�y��{cm�0,�p:��Vˊ0�>����!�~Z
�R&��u욢����(t'
yr��y;�l�Q��bǼ�N�DmL1}���lk����Ң�u��ȸ�.@Q��YW��[�����]�2�RO�Uc���a�ww�<XN��u�:77�0�>�e+�3y��[���J��}���k�{ce�s�Bٗs���*���Kݿe�=y5M({���? �����v9��h$ԎA�NtPz��l;�� țE��k\C���'��#7h0�N����m����Ҵm]mW5@�sW����-�q�CH�\G�$�t��T��*�#��SOk��t��l��R��*�Ps��R�]�$A=ڜ�)�'��MAeJ�� Ӗ$���[�������8z��9�Cɓ�V���yE�u;���"�J��C����v��&Xi=��g����c��;V��+9&�Iy�6�.��#+܊�ȫg�"�I��v��֯�";�&�u�fNJ�����X
����t�L�\6m�&E$ݢ��I�c��)��1)�+_�ʀ�t�t���|.]����r�5a��3Q|=J��	�|]i6�h3B�,��������[�����߀��@�Ng�Wp}(����?������o��T����/��Ǳ���1~
ah�v�ɛ+hST��v������'QDO1nu���
3R�b"w=M�6��O��X�zn�ΈIcB9����D�'4,�wΑx���@����Lp6�v^b�G��Tsn?9��<�g�9�6��ő�$��/g��S]�t��#��Yy-���� O�6�-�P��lĪo?������q�6"[��^��x�Ā=��� �����ԠQ���7߆�T<դ��>:�"�����F,�=򔖥-�iZ����l��^Q(�bQ���5���z��?��	�~���8�l�o%��#PE9�c�8LCT����v��#_�qymO�{ȳ�	����<A��~�y���z=A��x�������÷��z⭈�(]�i���Τ��uӂ��xM�����g�g��'/h1"w+� O�EZR��VN�	�y�"Q��;.sE�UJ���!�T��ⱜ�Rt�G�cO����;�3S�|nC�ּ]
�ǜ�F�/��=�[������""��`;�r�+�!��Hou�6'h-��+�B^�hl���ogX��yy���;���wc���]��un�'A��LST��B�y�jy��>m��ӵ��������em�w��2�ys'BE���mAώ�	�$v��t�:�h����p+�M�AQ2]�T?���� �4�Y}�*%{݌b�Dy�7��E�	yT`�~7Q<7��E��P������]���cD;��o��ȗ55�����JD�1�ʅ/�KsP։:�{�W,��X+�I��L�w0�ن��5z��\�Y��^k����7��{�[�o2v~�>V�Z%s����gE�Na�ԏ����n����m��(�Զ)a���]����T0CpE�R�5y��4���7�7��u`�>ޥ冗�ԧzz���,/Ge�f3.ׄ�5�=2��>�=��ct�V:xbu���eߛ�~�ė��C8�h�~JH46E&� ,	�ὐ7���C����T[^�R_��=Ոʓ'���YZ�7�3��k<GW|�F�;y �����4�m7���Lg/t��",sw�*�uʍ�M~�(��&�MqCQxӣ8��Ȫ��y���(74���_���ft톜v>H�����)lKm �t{�$�3�D����N��J�}̡���k����Y�g�c�I������sz�;~^����(lO�s��*�@\��) ��q��̦��n�fޙ���@^u���rfCD"6$`}�q(��;"�P�@��j�����ݵ[}Mq���PO୦��l����`� ��zg!OiT̮V�A����i[�PO��)'�:E�%�c�@pԴ�a���Ц�m??Cp����ڊ�7�<�YH�s~m � �O��DG=j	�����<+����Y�̟�������Ğ�H#w����h� �6{J"��;րW5�k�苦#̺�3Z3Ge��$�2����|{{�0���bO����^��j�D�	��{ģ�`Y�N�� ��'��60��1������=Ŏ�J;��ţ�#�$\<@�TIG5���Wɲ���hA�ٞM�XIc��$g!ς�V�s�@O�괁�d���?�<�@����:�^I&=��aCP�x�(�/A�=ܬ�g��c�6,j�<�v�BX^M _s��ȼ��ŕ\��<����I���S��
��̲�ӵ�Ƌf���oU�6��r�M,����(���'0c�}���fv>��0�~+����z�E�a�cXıL40�?��A��}P�61��A��v��������4V+�u���$m���f9l�QDʔ���i�2|w��Xq�]XK�P�Lpc���e��ByoM���<#��A^�C�[�\�t��`C��j;��,#lDF�� /��dy۝#�}%eTfZ�G���k����ɓ��Ҋ�uRJ�x����t+C�kM����چ*�]�6���'��"�ۍ���(���r+'f8-�F川���Hӟv�ii�ɾ_,#L1y����[?�N`�v��$՗��USy�����s�x>�D�E�g7lw h�D�a�S@A'�x5u��*�i/�1��z!P�h�ڨ�H�1K�OA����e�S=�=��_ ��:�:�ZS�%.�v��+�5��"y��i���9�{�ڄ��^��}��Ԑ�(�]`�ޥ����>����o0;^�.Ǒ���;�~�Zwk�ܕu��l�-�ST1�NV2��N~���Y�1��?+"�:,��Q���=�%�?
���;ȻT	��D�Qc�T5���Xu�TBG_t���Ɋ��(��}0��������K�(��X��I��C�wJ��QJ�(4E��Q�4%�<���ͺ%o(�I���?�4J��~յ�y��t�D�����TK�r�b������iw��eSXM}��Vi}`�o���)���b���%+M��J��2�{K.UD}��ۛ��� �Kw�uR�cm�	��m�����5�vy+X�l O��H^mS^P8rc�c#a0�����������,���.U��\�ϥ[Q��T4ƌ�z��9�rQ�LH3�q�vA��z���H4-�<u��)b'+����o
�'$�[ E��AOb�l�-G�G;l3f5f����x1��1��ă�G9M5G�)�e�]�F��Y	�AgҼ�璖�<xW���^��o,����iw�O�y<��f��p(���i�kR��������?��8Ru��D�o_!m��X�鍲PB�>�@G�b%����	Qg|XH���M��$4�@�(A�H�x�1k�t�����l m���F���h7�6h(]���ղ\-�c�ِw����^-�r�eQ#[� ���*T��c��5�@�#�Q(�h�Ҕ�||u�[��T�W��Zow������Ŝ����<]5���EӴZO`O���o��q!���3�G�dg�:=M�v!�y$��)oS�.H3#Y�0�5����	�z�w�v��CJ+�eo1��M���Υý׆�c��Ϡ����b���eO�y|�����ir3u.Qԅвӵ7
�ߊ#k6�ro:���M�K��b�����k�@�/��u��1�#�����y��hd��;֙ J@'��Fyl�VȣˍfA�mC�UWgm1�Y~�.S9U�������K�͔�AY���� �^��LS����7)�SMQ"��9�� ���*���c��tmF��(r��dE˔z(��Lis���z�I��W�,�֧�{Ӽ�	�-��~��#�5`���Y�L�̥�����;�"��V�,�mգ{$vr�j��6W	��S�ݍ�ct�)�����<rN��`{4��X�gA�=S�_g!��b)�%܀"��ޟzD�V��Q�'��ԭ��/��'6Б�h�L뗖�`]�d���U�n��yV;]J�Ū�����y����!�q�?��g�;�X�9s:YGՕ�o)����%ϡY��2�����X�e4�+C�a냯���6����S�����P)����� $"�}i�날��f��ev�Nt�g�Y�il�y�;���h�E$bca?��F��Yo;���)�}e�������g�X㢥����������wtM�W�NE��\��]=���|����k}Y�-A���WBȋL¦�A(��Tg�4�y�M/~Yc�������ֿ�)��\c"y�tl
hK�<����	,Z�6(k�c���L����d�Fa�A:0y�1���0KW���5��
v|���������R���m�(��Vw��N�f��*C|C`!/	�#�`cDw��W"b���?L���.���\�kSB_�Ҟ��7şg��sv���|���yS��~������f��)B�����v�
��(�u�k�7�PE�lf�m���Lu�5@p��=I��)EW�� C�k�;����=A��)����֌�}$���!��S��w�A�i�>��Md���2���k/��>b�`X7�kyW�Iȳw1)�m��>v�L�@�i/J~�'����m��8����D4��ֳ$��!�H��|<��+LS�����T���l#l���h�A@K �E�0+� +Ay񴓷�C��*5-�<�ʖ����#(��6p�F|j�����Hў�E��Ȝ�߮�����qz5'98�j�p� jI�ڹs�޼Y�I���<%E��G��3A�\0�����i�5���*�mT������pc��8x� AI��������O?�EA��8z0v(?ᩞJG�d�ܰ7W�5ѸZmz����FWv	f�Ƅ��wk:mCHd�� 2o���������͉;�{L<Q�r��h���[1kк$b�;M���*�� O�/TF�Wk�u7��4�Ӕ�E��C��b�#�� ,�n2��r;�"z�)=mPD̞��������T3%��e]�	C���_Y�KJQI��(љ�{��ޓ"5g8���3olF����|ҝH�|r����5�L7
N
h��Nд�����M�����moNѦ���Na4*���Г��h����Ɩ$Ҫ
7���X(�j������G��!��$lp�3GZ�R�(O��I9%��i��Nޭ lKAGw��	mt�s�B�}ɍw��t�٧d �`l۶F�Ű��R����G���d�}�ڱN��a�X�r���gE���%�������,�6^lg�w�E!����������c��ќ�q@ �"��&"H��t�K�_��ٜG�[���ix�M_i���wSgkW�҂l���I��
8v3u<�{Nb+G^h_��1ˆ߄cӗi0��ѿӆ�7���}y�+���wQ4��m$ө9H㵟�l����sܱ�kÌv#�fQg�����c˨#�s�#7�/�B���ޗP[T�a��r���[�yjP�� ��mļQ�"˿/�'Y�/F��v1P�M����_z��0��vGNX/���Ga����X����1��rW����Sdo��r���og�YeS9�ņw>B��6�l%�n��'w��B�2�H$��!+<��ӝE{PDGvgdo�l����	!���Px�3-����~�z�D��R��7���)���UX����P�7
:
N���d����$�N����X��)�����#�R�B�/�p���Zd?d�Eʐ��{�9�ʤ����#*�*�T�}���;Pv�K(�jv�j�x5�;-�2����'	ٴ�%1}�#"��\������;����,sn��H��F��q(��{S.u�KA�9�Z��a�Mt�r����hN�w�6Q�iCB�/� �9B��N��#8n)SMӤ
�
�,�ڠ�h|	[�+P��uu���{|_<An��6oR������C��[�5��ϼ�?7�i�����!(�<*��6�H4��<x�iSA��`�+��gXJǠ)��b7Y)��('4k��S���MFc���Vݞw�ɳw1>x UU�ԥ֡.�'*P<�Sd��4w7�
GUd"�I�u�|$y*�(Q�ڊy�m�1����ZD�v0�k��Fz�F�I�I�$TSj	���JN��ص�PQ�A�<Ї�O��`64O�ܩ�M�������E���:>�l��}�(>�h�2����ֳc�o)��@ŧ�j	E��]<�=��1�+�B�T�k1h��4���N�'�V��0�#�Ӊ�����������Q�Rk�KlM|4]�u
a�R��[�N�hچby�w٦�E�C�aް�X6v�ڕ��
w�쇲�4Є��Nz�䅢½%j各m��>�[!�.�%!O6�����r���a=�l⍘=��Dպ-0�V�5A�"T���Cì<�&-�Y���.�Ly}k݆����I'��g>^S�c'�΅<���F��A�'��	�bŸ)�o6�XPhR��;yZ�GG���F'��X��M��J�OO��:*"b�]иW�tC���׽/y���!�{�W=?�&)}���a-�fy�ԍu��c�W�:	�t
�ڊ6c�̅t*1���K�	y7܎��[�Jux�6��2�zj�l��)nw<�E��Ea�$v펽�0s�d;��������ZPEQ�S���DF(�-�b��)8�H� O�r�?]�ҧ�z��VO[��ݯA�{4�O �?��[ 6S/���b���T�&º���ٗ�E4l�4�6f(�	?+o}��X.6k颢v���=�����sw�L#J��=UN�&9�ᮡ8Ⱦs�mT���8�cE�[�	4s�z>���}�XVLdF'a%��QQ���8�����Mߺإ�$�!O"Xo��F=��Y�o����/�&r�f���O��h��L� |�a�X����5b���ָ�(�J��썥�:�]�j�}͟�<�a<����F��� 7q��v��+l���ry!��r���Y��6<	9�t�	v�ui�J���4(�D�v�=7GƖI�6��ǿ����sS��^�XY̳���~�����&�J�U�X�1��9؜7��}(R��FZ�VL���Kn� D�F�|Nx:���!h���	{�Z�'�K:��@�>��������5�<b�N����+*]>��}Q9;�FQ����n"y:ڬ�����w�}P��ZB{ol<�����(��OB�T��՘0N!�~}�>�,���D#�"	7�ӧ#��m�V�n�z4�E��T �ΰm�k	Ǭ֫u�E#�B[1'\D�>�[�#�/�M?���&�u*<Q8o��r:� c�&8��PK�Ak��bx���h���(�3���t� �� a�	קY����n4���'�I��f�����@�!��q�E�[K�,��i�#]7p8��������u�ّ<A�ɚ-���y�䥏e[����5D�@]hI5�"
�4li�D�B�gEӼf�W���K$��`�Y�Z��Ӭ��3R��AцF�	l	N�w	q�$q#*�g7RD�ڪlB���z*&s,
a��3� G $�IVn3��Fp�
"���XWwupC�����\���@�~j]�	��=CM�:g+��~�m�*�����{����u���Z�D� <���-���u��عb��x�Z$k͝��`� #m.u ����dY��4%;}c��K���aƐ>X8v0��C̦������زa��W�=�����3�����F�~b���W����G��j�(_�O�w>a6���P�:g*��r�mn����X ��(j�_PS�v����ȋ����[�<�7��%u����FTUך"�5r���UX�¿�ٰ����)-����M� ���t4�$�Ry�q�k$���<EAw*:��S���p� +ȊC���sAO�����*�'Q�� �?���f}�V�H+�������s��B \�@8'�Tt
�#�0����ڕ\��,�X��x���@�ّj*�"8i{��yo	N���[�y�C���2�(94��P�2Iv�,�g]��9m��e�A�Z�\�d��N���ZYQ;�n�z<5�%.�3]�6?��b�K�͞�<��� *��n�8�/���b�m!�H���=��ikWuj��(7������^�����i�<Uoq1Qy�v��6r�disD���խ?�\��D�(T�I9␀�Nq���6��!�Ä+EEubC�w4�}�M���a�ȍf�a5�pjl_l~�e*(Aف��;��R�k���-��c�DX�U�e�0�-oq��&B�N����:�J>�C'p%��<�,�G��N:2l���A(�臲��Icw ~8v��ۊ�kS��x��.tY�$�G���ji��`�ț��Ģ�=�c�u%�����U�GC�!�/�cz���p�&�(�;��q,�
M��^(���7=�%C��!���.�^���%n�8�Q�B)'�}_��V�ޭ#�e���AcQ�{6��r���0��>��I�dyK#��0�/�߄���8����,�)u\���OR�B>�L>ң��~F`{�P���t�v��Gy�����o���ǜ��7���;�_�]����`�{Z��?�e.����wU����n���L>�j���w�z�@���Q?lj�^����0��s���h��<�Z4���A�@��"z-�<��F�f����Q�ql��8>f<�_ÿ��s�G_��#���!W��б�5��>2h�]3
�&�Ɖ��P}����7���&�čw����Q�����q�Q;�&�_{#���o�}nC݄�Pͭ�{3j�LBͨP3z"N���F���L�\�ڑ�q�����끱7b7Aq���F6���=�aW�T5_�I:�$��iM���U���y[g����7���%�L�Z�gCTN�Ǣ10�	r�_�m����cD("q��[ Ϗ��f�n�a�Ib�~ֿ�hA���J�1����s��+C����p_��3!	&#�ʩH��T�v��LP��tP;�]$�9��Ӕ��n��&���N�&��=8`L���C���w0P�{)���(���/A�����M����:��	�N�د��1�Dlh6�It٠g����d�ͥf�� &țIX��vT[��O@.���1ȸq6���*'��A�ߔ"Dy��xZЧ��:jN���C�^/�~�ٕv1�;?�wAȫ>��w<�ͽ��r�8,f�Ͼ�Nz�Z��YHІ#��@J+��><BE{*�ȡ���Pc=�O��JR��ci�UjD��1p,���͋�Ǳ꩷�f� ̧��ľ�AZǵ�;�lD�4�@ꀫ��#ๅ����v�%<��\^8H0�r��n*Ғ��$��ʹ�ͺ�n��!�,�@z����َt޻����@��Z�~T5��j�㊮�O�I\xtG�m��C�[!OP�{�=���6/u	�1>U��7<a�����3�8��Ò�֗-�	.��c�s9�t�6p�h�����X5h"����!���˰�~Z���)���ǫq��߰:h�{���l�{S�uɨ�c���:�b;u��PY��!��kQ<�z,J��;G�o��~�Bde�7�ii���j��%��;ξټ���7[=���9����k9%a�k��ŚS~��Y=�ɾfN��GM�.�æ�$M2��)�"����p��;��5iH.�6�B�g�B]�j���{Ȧ>��Bǉ�C�t˓Gg��#�$`^C���+˨�7�Ķ�('Jv��1jg\?��q5v^� �.'������s!O�S]�[&�G�L�!��8ᓄ������T{ap
�$$�B��1�5|"
�Eq�B�pE�AI�/�/�u�m7?��4B��Ŵ�*���.q�8r$���P������V:�p�y4�����Ե	}���H9�#& o�(1�#ơ��Q2p8����}�O8-���	w���5�F��$
��a���u%������[ͲE�s�\�����l��(�9�D��v$t�A_o�����H�ޘ(�F��M���Zl5�|��������8�>yO���Dè[�������0��jB8����Ј�w�4�	�����a�PA8+<��B�����w�X��	8t�$&|�0o��wދ�{B���Qu�m�?nvkD���eW��N�{�Lā�&���bߔ��w�$���s��8x��8���8���8t��6z��ހ�Xrp�-�3v���m,���Wck��M]�<����F�����G{®�C�w�0��3;�z�:�b�a=�U��`n�q���.t��k9ZF�.��V�Ʀz/6���7�d��	��1}QO��TR_4��@S,a��g��J3�q}���&�V�D�4b�Ss��C���~���|�s=���P6zD��eԅE�!:�1q8�0jt"#�pF������h&6�#z�:���TO�%�X^J#�+Q��ɗ����~	8@��K2��0p#aH����P���D�b-�ܺ"q�CM�	���|�u��>�;hNQ��W��),'	�'��Z�ҺԄzc�cw�(��0�
�S���<I�H��Z����d�F|�g$�����tv%"�?�Q���&��x���<*>�}�w	�Q�`!�d�j�s���.�8�0 �<�ڌ"+�Y[E�S��@�~d󋈁�cXu�8�s�����߀c}�|*�]�q�Py��ۈ���p4�RK*]�Q�j`��@��F�@�Xl��_��[���7�c���N�G]&U�>���Z�d^�G���c����@^p �8:a��?o��!F'��B�s$w�2�6���hWo��*�H��mA������I�8��:t���.y�|�OJCC#*=k{M@�ww��qo�?���k �I��g9wue{:z�<�����|	Z,���Ia�H�z�Dd��(P���tOޔ��4��kr$�3�c/�ړ(w퍓G�86����O�_w��r�u�>����[j�t�T�}>(��EA`0�*%I����fM^����F��ڠ痯ͥ��(�w�
���BF� �Ck~u��rjz{��>�TZ��x�������&ހr��C'"��h����~�#R~�����j�����jGK\z��#U�}��(�dT�����5�Jꪃt��D�Hp�t��n(���Ñ�w42�Dv��(�C���1	��3;�K�_z�E%ؽ�z}�>�dX�p.t�~��R�L������fc��[�_�'uVqt
	��ԟ��1(�3kgWG��ʄ�X�s
�����4�=ht{���n����m� ��'qxm�Y�|x��D5eA��&Yeյw�l��)������=G`o/��#P����!k�d��~;��} ŷއ�7b��x�M�2f2��r?��$�>;x'�JY���Ic�e�]�R;����'�Wf��a�P��p�Ƙ��>|�	p�܎����)�!��������6�y=�$��%tl��6������TLB�=�֚���<��S.z������2��UԌ~�=ǘ5u���k�܇m�?�mw�1��q��� ��z+����8u���^O����r���q��(�� J���� G�)x���N�D�Os1������8���5���1=���k8��@Q�a�H��e���Rڇ��l)�-���o���縷3�"z���rAZ$�G
���=!��`�#�d�̱���Tm��g^��8�GY�Г��HZ|J7�$�<���I��g��(��t�"�E�������?�΅�`�����r���A�jEK��{Z3Z��!1�Lv8?܃��� ����I����� �bC���c8YW����s���>���P�V��A��1h0�T&�z3�@�<�ے���q�����^�Z�o������%ř����A���}��Lϫ*�3�����3�}�a�4὇G�@=��G�ߌz�H��}Ơi�5�57�nn��0w��}ާy %����L�*q��l��TP���o��|���|'�L_�\���Є,� �N��g��F\�F�F�oy���ױ\���סn�p��;����p�=�D*���⇤84_�zB7�Ņ��@�־hʷ1����	E#���0*]vAl/̉������n�O�V{��/u��QM�=F}��{B;�P�Ox�'HQihW� O�kz�
5��S�Wu��|e�M���=$�4�$ʸ��	�0�`g���Z�"8�C�Q�G����x�5[͏����㐎�i��1�L H����Qb�� ��h=6��%��|��y�{pй��22��p�e�O�q�{As[@����|�̚�J:&�Y޺؁��L"P$� a$
���Uo�&:sO��C�[���~���2{���˾z�J�**G"(tx�PAV���!*�
�}1�8�C�qF��	\����D����4�}iT������3��R>���i����5��׮�����S�Ơ��*q �$����8�������q�
���P����p�J�*�'6��a[7����N��M�?��@�,���\��]��\*�@�N��K�#;�Z��w�9�'1J�2i ���z@U��8�k ��7��ɓPq�M(����>l�x/Rz��|�9|���lS��ӆ*_���3�w�$N� Gn��D/�8�D�`�>�}����(�!9Lxj��j��t-v��l`%g�]s#
�N@��aX?p�Ӊ+d[�+4��j�F'H\�·<E�M$�T�~��=�ݏ
�ü��ؐ��L3v�Ml�l�x�^ðl�H,0���O��17c��Q<p46S?n~#v<�:��m��Ʋ=��6��T�s6�m¶߼p%v?�6p��80�T���c�E�xB�~����d>�<v��v��6
y[y�yǧ���7>����Į�F�K��h�iKwK�L����)�m�ly5�nũw�c���M&��k����{�$d�}?�}�{ﾇ���F���!繗���3ȹ��L���nF��`��.�c#�T�<���䒗
Xӄ��,E�u�a�����g,R�^���M����F��!��7��ʛȞ�"�<� �D��T���x��`O��)�`ۣ�Rw�����D��/a�u�0�F7���j}WE5�{��7��E��0m�=X�0i1���t(ؖ�Ӊ]��~Q���?�D�%K���g��O[�k�	f��M�}%{V.�5�Ut�V�QY�hֱj�fZ��\Ϳ�.�;�hW�����uat���2"z�3ZZ�B{��+���u�J�'5�;��	���ZÝA8[��͠�F�A^T��)�c~tߖ�=̚L��+�B͙�[	��!�fM�v��ԗ�tD��M��"�Y5�뒐�#d9����P��;l�a
����u�a荽	PN��+f�1�۩���S9s�K�&�2�%qݍ��z��4��%�0R��-�@C�v*�]�Fa[ϡ(��+�`ޗ'�%i���-��}����(�R��7E�a3�6*�m����:���n¡GÖ��D��[PJ��<z�	��k������¤�(�=��J��uq���L�Zw�3�:�f�6���Tr9ۼ�Ì�X:d4v�����;����7`;�n���:z�	�;��ǞQ
�^��CGa��1(2�Y�����g�F���[��c&!9f>��m��5�Qt�VȻȥ ڗ1l*݁��<��G�b�(�Hb}�x��p=�k2��e��}z�,1����g?���ۻ�Ůn}��@���$�LzG2�t�	E�����H�eS�룺���WѼb	�%$!'8�q������}PNC,)�1�ѭ�)���^�ڣ7v�8��Z�Oz��,f�pO�U�:EL�_�^E��E�w���&��8�z��������a�����8Lx/8{'܂�'�b/!���7���oa�8r۽�{�&���	Ѹl|�C��&Zr��G�gç]~��jc	6���F߄]��c+۴d(e���w�]�;�-b�5�`���Q6�`@�d'��A�L��z�б�N��������oHDխ����2�:�/=m�R/^��m�8��G����Cơx ��D��¾�Q�gJ���f��n���Q��{�`���(�)���A�#��r3J�މ��^B��ͼ���Ku$Co��ٶ��%��R����֗���k�;�3c���p�E}�"t��X>S�������F>����a�{���ב?���1����7Y	t[�����΃<��{~[��������";~6�2;ysz�z�º�$䲏o����r������B����x܍X��6��ی�`��o����,ymA���R߲���\�f9O5 ��XJ 9�'~��/!a��3��O�ρ!�1 ?����t���??������g9�a���k��6=�:�v��	���0����O�껖��P�U����#����b��ܨ$s��Jҙ4�3���,�
��y�ݏi�܊�ߍ��ށ5�B*���ފ�g�����&-�5��<ÿ́m��a��v��x ��F�7�n�A`�IP�G����|��c�/�ǞįO<��ϼ�EO�����������+���!�1릻Q�,��BK�qf�w[��:q�8�~�3���+��d�b!!c&�d��o`ſ?¼�>Ŵw�ǜ����އQ��]\q~7�h̟p'~��̦s�p�}��zPI-�F�P��m�����R\�A^SU=rޞ�Y�Ă�1X���=V�X�`r�#�\Ñ�f���A�։!J*��%�E��K�݂�\��aH�wLnBW�GI�
G�G�7�I��Z��|�k����%��#��	49�ߣ������j/�� %����Cj`��5~�X���n�H	��6��r�@,���
$��>a��
����k}}yod�� ;0����!8ya����y�57݄}��8Nv�z�i<�ޮ
�>P��J�}��:i,Jx�
R�N�6,�K�&�D�XW�g2XX[R�Y)�!X�*)�|�E��V�Z���[e�Yy�R�����1��5$���D>��u�Y�����I����.��X����AFx�`﹤G�s������c.�z����%����X���	X��E^�X���`�RK�*�7��=# 3BI�݆`u�� =0?"�Y�y������#�L���F�O��_|1#0sX�y~a���.����cszX�f'�F��!6?������Ү4��#���I���TM�$
"�OY4�$�h�(1�Ċ$D*.�$&A6YB �cy �����D\�訠1ə���S��cմ����^�������n��`�=��,Bw�az�������0z�%7�ui ��X��K����*�?�\�c�C�����2YG�'�����]+�`��;H���#�"i��A[p���+$��"vb!y4�kFd8Y� � ��$y��?B��*m\�H%y>v'2,-YW*eȼ����Y&wg�|b!�m��a9I���n�@to�@A�B���=����p��(~z�]}�q>�O� >|0��_\�D�U��F��
 g\}���g�G��/N�����O��'���QNa"�C��ܼW�榏p��QK�x��i�Z�O�G�'�MG�tN]��y���+�)���S�I�+�ח�a�4��j��P�j�ٶ���]iϲ��%�Q`ɞKՁ+��r�u�($O�%���=e����?�n� ��vY�G�7�d���G���Z�*}��j6���C�����PL� A��}���XD)�N��J�P�����9�3���*O�Ս�<=�	�!n_���8�o1g�L��Nb�r��P=��Ϝa�ԙ��.s�^�*J(�R-�b�ڈ-��X�ֆ�ef���]i7R�O��|J�I�ԳL��J���5_�� ����?T���O�������
�:lL�E�h6	����Au0IK�&���_��ˑ���w���._�A�~�7DOڷ.I����<�UڜT�;�q,.��Y�9�'�ۣRa'���
>10ç&��rvŞŋ;�1�{i�t��]=�����F����������4��$m_x�чc(K<���H1tA��3��XX#��,M5_N�@�+$�_��E}���ñ�d�ވ�Uo"��s��B$Ql$�ؗ��Cg{�����{>�'�I�nD2/*���0}!���`7c�n3kl7R!�eoTDǠ9���|����H������@�A!��&�HF�^	A
�N��h/����Zq#�؎��$�5٧T�����alǞȴt�>�������֒Bhj+PU^MZ�b�M�����ό��9^���������C��匯ɓ�������Wǋ+���̒�u%U"?p+�[0
l}Ql�cn�tb�s��2k��k�Xճ�1F�A��	�s%I�����Y�k��U��v[���Q���GA���P���y^(�w����Oy}j��M�Y����:�Ũ_����,�#|���F��"���v	��9�/?��*�ϥ~h\�AˠY��e���C]�?��/C�kAh^��k���F0N��dhډsa����58�6=�������B��� ���J��#y�oh`��14د��]�4����
���iGWv.��b��h��gd|q��G\0�F/	P�<	��1ΙZ�,�<\����t:Ȕ��5��XYDx��m"�����㤱-ژW��vǺ����h�*�c�W���A��>�-z�8>�,��
��z�Jy֞<�A>#j��$�/Z*h֛��ɼ����Af�w�f2|t�S�O��c�j�=����6HV��E9�W�3kL�0xﵼoA��)*��AM&�&V�s�Q	A����4��IH�ꊾ�$y�F��-��;Nĳ�\�w��];сx�e(��F��2gg1��z�'a�է�&�*C�j#�hs���T=U����jE�B{�7�$�6[�
���[ӄ�~�K�	���c�.��R|���;�b�r��zo_��S��� ��Z	l��N�0��2kӷf��XG�R�U�f"
���k4�S\P�
=Y�Z(�WW���2)azt���	���ý�.�h�`[9B'��R,2P!������C����X_`��I�8�Ŋ�m�2})+I���V��h�V��M�D�q�l�E�dTM�>�{��Q~`��ٞt��6(��*���渏a�B�_!�Y/S4X(�P ��a"�r��6y^Cr�I�t%Fed��EY�͊v�]0��	�J�r�1����JB6!n�,V�BUg��)�L@�43�M1F�����P��m8YT��<?lf�4
�LC���|��,e�=�2���g(xV���KȴP�tĚ�#�}8�-����6�Y��h�)H�<�ӌ�����L�=��� 9� VOR�����gp�X5
c��Q�V�kBO�ҸMe�w�|K�R�}�k�I�tS01T �$T��#3�7��]���[��:*�#�{�R�;9�p�V�L@��8th�py��B�&
�k׮attT���OF��)����M�ۏh�}�f3?kD[[�cslUMG��[f�a��Y�D���j&v,Z��$,kג�xa��'�� �7 �|P�7{�� ��s��h#&�ھI�R��	Ʈ���]q$���s������h�=���mbf[�3{+D��Cz�:t��>/�{w�P�{���>��ـ�!!���2|�
?�Ơ,	�@���ځ?�}ĳ�RN�c�wQ�yI�>���o!nE�C�B������� kgΨ�pFS���B���!��h����ooF�|���ۑ�)r��=�'᥃�Ok��r��[�n�xE��E!q�:�)�o� icD�Gma��O�B�y\=s
h��I����h�2�����x�b�D��]�v�>4���;�A�ԡRQJ�ϛ��b���N�>R���T��%�))�)ђ����D�LND;_ӡ���y�� A�t�Nt>�gs2p./�������ᰂn���ED��q���#\�(Fo��*}����G�'���T��F5.��@s�[t�`���Z0�ڨ�J{�����z�#?t��N+��s
��:q��w��x<���q���R?~ �lel�~r�T$}B�Z1    IEND�B`�PK   ���XL���kB  WW  /   images/e3ae6286-4af8-4c7d-b449-b4e8e59fa08a.png�PS��>��Kh"���HK��D�B(�Бދ4Q)JW�:�@� ��wD@A)Jѻ~��9�s���s��;s����{������Yj�CC�N�h.�j�@`K௖���~i�4$�A�5��oy�������	,� ��^��2܈�o V�~[�X�����;Z����^AR.-�@�: ��R20�(�.'*!��"���������:���?�{x �=�1h�4���s�/�a������	y���>q8��rl��w�Dڻz`<}��HuG$��U�c���vvG:�n��;;:{�Q�/w��6�k���UGx�9c=bwGq4����Gz����8����W,�h膳���;���WG9b܁��3B�a"�~�������Nb�pO�9ȟ`��@yy��1�������B�=��D���pW$�P��+�� � �(G'����=�F3޲���H��� �/���x�lz&DeÁ~�)���}���ꙓ%C��gW(��+ay'	�|�d�P�t�D!1:H4��:�%W�#�x��qw�{:;��X��-g404yI�W����l'��,&-� j/#���#��piRTVJs��KK��0ǭ�8�4�q��9^K�K(`�<�o�KȉI�o:*���%�u� J�b��V��3��|<�n'��*����'T�������rG��y QǓ�|<)?��ώ{��rG�
���?�n��+vٹ����u�oә�7�a
-��)R�n�4.d����N*�_U����]�ЮeQ�KƗ4��P��}AN�9׭�֑ Nȧ)�?��Q��e�J ����=b�=a+E�CZ��ΰ򅙓�C�� �0��\b"0}�WO�����~�Hlv6����B�n�LM
�z����d��I�����|�#�ɪ���D�z�^B#0�X��>�qA9FԌ�O�L܁��5F�{;#�0~(/�11#����{/�?�:�Pn	)(�_@Q(B%$���-��0(�q-
�Y�c�2wB�{ˠbّC(��h���_v*M8�p�3�_����{(���&0X��m,�h��ϩ�����t �>Q�2*�RNUo��Cwؙ�q�H�,D�e4^���<��Gą���T��Rf��l�z��S��=���T��4�N�����2}nDs������$�]�U��.�[�0)��I�6�}�<Ѭ1	����m~�T��<��k�N_���o@J^�Jzz�c�����6#K�:�p>*�j���Ā�_������K!�{�r�Ŝ��N�ndW.޸��˞Ƴ�rBm�Z���F
u��_@.Q�3�2��f/�Zǜ��������\�l1D�$�HL-#���
��Jt�	1y0�@�,	�������2
a20))91	44�`�K����mED����eIDEB�/^ Yx�O^,���ٓ�<1�^H^O'g^=`����&�3�����:������ۀ=�����D��SjM��)�j�{5� J�7Ba]�E�(1�ۮp/O'�NG�md��I8!+	��JAe���0yI��f���t����i�'���kD`0�0T*�W
����%��gSPB�HX��!�o�I���A� �sƣ�øh�ֿ97qćx8i��	]����D�{)�W~� 2����}w��9��&�����ڜY�rS�Mhx�*�M#��L����W�.�W1�~�S3�=��R���l��U?���P�d<r�C���c�y��,s��u�#[�����ϔ�]NE�SO��N�H��V�0�ߟ�Հ+�1��g?#��y���Ց����{��W^[�!�|�W�<Tr�f6�����k�3��q:���__l]U�L97��Z2<{�!�����f�"���)H͸"]�<#��<L�0ob	=_~�W�dݑݙu�	����o��Y?`^��o)����7d�@c�����Kx�*��J�"k�GWleʔ��ID��p^6��e����{{��хsJ��E��X������9^��7�%�܋�A�^[�Z�&��6,�L����3,��7��4+������ou1<�	7r��FN�������Ձ���
Ib>�y��y[W~)9sΟ&�=k<=�Ǘ�������Us�| �a$��!���?��Y�W_\F�¿C��yH`���@��c#ཚ�:$���`�#� r!��G F�?�?!��p�Z��F�J+]�OHx)
���٧!*��1���ޡ?~p}K9�MOHO|�a��
���O���L�H�ԯ�l_ڹZC;���Ǎ������|��lsw�~��v�F�����[eI$fCKi32��_g�$�R񏟛���x�݄�4�����r�y�$FĪK��x48���[�̀|��"��J/F����JG��̖`�n���]�&���ߕ������Ee��������փ�=�/��8{ �b��E�uO�|ku�ql�
j��Xp�3��]��1$ed�S����G���,�38ln=�n��f��&��4�nm���C�Q٧��!Kw�"�T��3���7�����E�~�E"���#:���?�������{/ܻX.����p���[�����ڣ���^]�xT��H�R��B�{�~ߟC�f.�jT��S��e���M^lmv�fX�����|� �t����qV�ţ��,�(:>�6�:z�j)"L�pC�R,��Dd<��Rxc���%f�|�a`v�<�� �I�����(�d�?`�@�O@D*��{>�\ԙ�d  ��_�?8J�ÿ�'�z�<i����'9��	b^�@���KU���p	f�Z� ������IWg`�	����0w�����+
z�P1	�AO��1AO\bl��)*�����r�hI�I�3��S�8�]M��=O�uoFƿ����?�[�y��)ѩ�9E�MнД��3e9�r�=[u�� ���V��&��)2E�����_1|V��;/{TK�����2EF�oo�D��F�}�o7�Mu�A������ۯɇ
<<<Q����o��z����������U�"T�)��?$�Μ�!���Sg��n���͡͜fr�l��I'^Zc�5�G����ִ&~Qam�$<���fZ7{>��ν�"�o�����A�}���Z�7k&�5@=?�j�|$;�zY-y���Z�Rn����6�t��ɽ5��C���U��Kʓ��a}W/���3\ȸ}�Ӛ��X��ƕ��R^�����Iy�|�qC��k-��������f���Uⱽg_��k�_?D䒧k~G�F�Q�������1�}|��qKK�g��~��qϬ黂�=�3d����huH���	�d?� ә\����L��Ǵ�ߜ����T��"��N��Fq-��9K�Z,Q%���(�t��GO�	��~�5F|l�M�2gg�7����6&�yΞ�&����!��(sZYh�$���Ta���:�D�a��-"01����l�t�Hb" \CC�Ȩ����`�\7(�>��:B����{��w!���LPO������������p�,�,@� �)�(�/�2l,Ю�4���J'ČTR���� �P���ms�RRnu#4 vaD_~�/)wv�(w2U�e�����G_Ŀ��4�����3�Ҋ��E���gJ���� b�#�kd�N�U^c]u@Z�8�"�=�Xg�#����K*��t%�`Pٿ@���P��I'���	�������Ah����<�jr`���@p�8�A&'� �苔^�A��z�i�i���b�BS����:�z����͏��s��V��!��)�c���Ⱥ��Q@0��q����*N���)��R�-B(�)Q��� #s��s�?7˟Q��y�U?R�C����W�-ޤ�n�Q'�´��0���U��Y_��'�`�5��Ͻu�@�#���G�f����H�^ϓ��s55ՏQ#����XD��U����cE�gKP�����V98����.y���+��Aa� ��� �u�z�'�z��Y������Oԕ�S��wAw	m�Čq���~K{z!U�$nO�e���ba{M�t�Wa\ǖ��C���bx\��K�,kjR�w�ޘ�"-:�K>0^����9��{:����LE6c/���^q[O�B�oK��%p8<O�/���
��yK�a�?鯍�a|`������y�Ҝ_��W���P� ec,1\�sde��~$y�pB|<E�q�ޱ���J�G���r:�Q��T��L�qW��\����kD����G��f�rPd?z ��F��yl~Sԅ#�﬜��5"=�:˖>>#�-��]�K��Ц���T�qQ/r�+ITÆ��0��n����-KkX�J3��P�jvLv;$a.^j��κQ�{�Rڛ�BKQ����&1��M��|���,F},��6�xW�����q�f6mڳ�_4n��Z�lҰ�(�0]1o׃��f��-��K��[˼ʽf���gj$zN���M�y�
��7���I���]�I>���n�� !R
��ߡ�\F���I��N��y�7-�=��k��E�! ��-��	,��=�;�Y <���y�@t��#��%����@Q�H��J8�_���(i�K�-�]�:K��5Y�0�Z��P�`��c�\ܛ��yZL6Oc�9�~ˌ���ɦ���H}�#�����D�G�U[��!w�Yg�&��Y��؄U4�?]S�1}�|^tm���k����@hx������hm����z�T��~���s��{W"쫌�z����٦m�L���в|j�63��w�O9~��G�><��ꓡ�z���y���Z޽�ހ���L����$���"���#�8c��TA���gI�L��a�����j.j"B��Ђg�+�1T��fT��:�z<�B׽�ܙE����<�_�R��<��yh��^��t�����E���SN�ve���s͛��^kL����z;�W�%C�'m���}��g��5�I3.]ݾ�M�~�����Ͽ]�}%�`�7���S����7��~�Le�8�ge���+ާ��(Z���r���i�Sā6����g�*����ܔޟ����l��Q�σh#L6�W��oBO5jgW{��uy���+�KlX�f���?����O��<�6�fm�7+樺\�^�Ig�o�#��� ����Ƹ@��7F������0Ց:���T�*@�rer��$�w���JP� �+�<��^��r�ӘǱ���3���7�t]�^�"t��C�B��й�-���m�����k�~�Y)�c_ͩTL�U=;.E�s��BӷL	`���)Ϊ:>G��+��ӴY��ya��-�=w�x�(����hԽƬ�,U��篼�-�
�+�W�7��|��9�f����>^0L��� G��s-�3�v��o?}bUDu�g�=!w9���Y�{Y{WK�-��N��������3�O.��qH�r�\�BdT t߸X���݃>y��_gE�U]
����k�2���j��Mq�*|�.Y�r�7z�僜G�3�a���o�^�A{��:���|�����j�������+[�6�cA_���D�E�Mb�����d�������k�ls:h���P��֑9ϡ~�:^A(
��+���^��)VeGIG�:�������H��f$fIb7A}֭?�A���΍o"�5�	ES�fIw���{�D�'d��Vxi�P\���2#-פ�{����H�!,�p�j@7@}�_�����(���P�N/�a4��s���<#�����#M��A`�Pv(HN������R����q穂��JP T���H`�$��)��R�ߧ�[�6NOr%h'��� =)?�&/
Be��]vzz
�6�� �_&��b�{A��O��Ӧ���QE�W�y�	a�X чD�M�Z��/$��mq��e�]~�u�>�	�;��Qɀ	Nm�����қʼ����C�i�7�x�x�}?�NYͩA���{����������^���{����ӵk]ቄ��)�[������Q`�o����2�~�����G	FnG��:�$ۅ4�)��8���ܔ�M�M6�T�m���ZmH����ݬ�(�S�2�����ٟWI��o�9��^���L\3Ln��=' Mg$MwvE�՗��C?P���/����.|P9-��ٝ��1�S�����bN~z�^'�]���!���w�Yl���F�?9{�Ѫ�{Os��d�[*m;OM#��/)�_��;�e>ń��7%�����O SA��5� ��������l�@��KZ�&�������T��/��m�ܜc��~RF���"�f��6fOܖ:w�	�\�@��8��?�Kwu�7Cۃ�b�C����}q��ɽ>:��z'ճ�iCa�Nm��_�oG���A΋S����#*������s�!L!�)���ι�ie��-�>�W��~Y�Z`[�=���z�g���Uk�A�W�Nw��~Ѕ#",�o��O�
=-(���f�o}k_��c�S�T[�o�F�=?l�#W��'�dǿ�w�:�8��|��Է�4�2 ��|X�� ��<�õ_9L!�1�)�D2|,q�/�$��,Te��	��"%�~�Z3���<W'�*s�ʽ���%��]�Tl�Pl��p�;T��k�OFR���;Ȏ��{�Z�A� �8����^��p��&��xi�/M����k��L����5Ƽݚ�Ή��5���'���?���0����� Dwv��h��ӻ��K�b|֭)��m�ζ
��W~x��a�a\
Vɬ�+��U�Π�K;��v��*�����4����"ٔ����U-��
�55�6OὢU�c|�ן�&_����g�V����5��_�oٍ%ZQ��𙀂�}�%4E��&��?�"c������H��Q������A��������65ن���ƭeb9j>�W�
\���A�8�!����j�d"	��/��x�&%��(�dW"�$�X7< s�u�N]�dl�e=�o]��H���z��ۋbB�.�R���潰��!)F\�7R�c�۩P���t��M����!�^�q�Q������Z4D`�D�������J��I'��	(���.ħ�k@Q�Lu��Om��_�e�L, 7��f�;{��_�i}��J���Ѐ��������nuoU�
�;���P�tn	t�h7�J�=�P�1���K�vc�%Q�m���m`�0wM�G��xz�{G�.�+1X����ڑ��&n)W2k��X�齆'��kQq�����(ռ�"��4u	l�#V���q^j��#Ϥ���wK����+�zɣJxz��`����%��l������&����&b�HIE��VV�G�&���K$!�:��.^�p���{�)ع�Fr:���h;����fu�������yV��\���&]��ѹ�'X12[�n�Iq�:��k��J��`�*%�cfM��f�Q1�e[��7f�b��_�[jV/�]*A�o?���2��kM�9G��Ƕ�}��qaTQf��t��_���~��Ѿ&ؕ_h�)�Jl������/����գ������7�#K��֚��i�d�%��^����W�mr��D�_FZZl�828F�-��5��#cg�*��m\fҰu�r6դ錆_�z nb(��_�zu�XrcY�2n������+�e�EL�zW#����on+uTqs;s|��u]?��|���Ʀ���MEZT%�S�TfVS+n�G��������V����0*�E��k'��u�0�����e�M6:K���E�ٷ
�r���4;K"9Xٺ{7�$�!��c^6-�<5h��x���*���$Q���T��A�QúGoX�}1��ť��N۞�Y�B�X[
�� {���G��Ϝ��yR�� (�H.�b�3�-��R���֩ddb拑�F����r?�|�W|M�/�3dF4aM�H�V�寈h�#r�~�9}�iȐ�
x���1��yi3�7%J���5�C,�>��q�_�.��$D���l������ŕ�s�
	��>.,zp5����T�ǘr5HV�-~�;-��S�B��y�(W�v����Bb��`���%�ܲ��|�Y+|��AҾF��{\�Ȃm4�B_Uk��Vj������ĵP�$ъ~��@)��gV��_dB3&��υ���_������ w�&܆:hcހ���͖�Z�Z�|)2�ehu��'�kK,hdaH�F����,��j�q8Nx�kPP���B�U�<b,?��3��Ρ��9�oOn3͔�%p�u��nyǗí�,PI������j������n�q����@v
�55L�O1a�SD�ڊ��uⶵ��o@V1�>D��ӥ02��c�����M�A{���J��T���ۗ�p\�4c�1S���������w~<Lg"6�#��}ç+�x�6,A�N�}��J~�����a#��uO�	/�*���������M��Z� �ƾm̤���ǁ$��P��[С|�,����*D���������{�-�ӭ��n�d�5QՔw���_��ow��>��A&Rֿը�ׄ�;��ע�4��h��I�xS|g6g�Ӑ��A�f4���G�Ő��)7?2�=(���G��`�9�H�Q"�W4k)�;�+n�=
W�̳%0csG�͛�>)����;������b�d�Ά��*�o��{�6��ԩW�#9����*���L!����N�cpK�B�z��/�ςm��f������(S���'�*�=�	����z�4>6F����z9x���T��L���)5��iC&�+Fo8ڵ��QjXMa���J�����p�	3�Lt�����'�����.n���ڗ�(?ѷz�{g��,��	7�k�A!VU��n���
�Z�؂��s].��	����#Ӡ*mEmC6��N6��̥=�+x@�s�h��(JG$˨�|���6n'&b�c|&}���n�]��~�\��loz�U����e�
Z"�)��⦽\@��zKPڎ�))�nT���w��LQ��~䰾ޭ� W��I����꯻)�HH9�{+�3ou��ӷy?�LU�	 [��1��[��ǲVe��n�n�2��7]%ƋE&ɶ:t��d�2\���9��?��0(�g^e_g�%Cڎ1?�2w+\)A'nZ}��N��.m��Z�4p��Π�uN4�l���ج�+}���n��%w���[c�T�+drr��c�*�-�E��n��P~V�B�2�UF4�]�K4�r���
��}-�Ky�9#�����K �Q�Y���r�T>�2Z
=+{O���&@��{kX����t/�.鵪%���j����l�� �	��A�����c��$���C�
�u��k���3e�I��5+b�g���=-��  mr*�t��O'ޝ�}f�4b�N� jap%�L|�}"SjS�@U  ���1-�#��T3�Y� ��_��,s%q�E�p�	�� �*K4�����κ�HN��*��T���H]P7)�?���e� ���v=⡂[:H+�db�v|-�Z��|L�9�����鶑��:��rQ���9I�Z�%��`rT�9�Ё�鵸���:�j���M� *��C��N��N/^����_�?�쩯��ퟲ���-ΐ���'Yj���p�������Kz�s�}x�|l�a�r���0���`9_T�	4�`z'<�N�N��H�G�#T�rq��^r����H��m��Ǣ_��l�:�v@��$J�$�� Fr�"�'G�6�@ܩ�u]�ȷ��U�E��� ��uk쓏��.g2��Ӹ`e0�7���c���M�y���=��v���	u0�|1I�zaY�S���X�,�,v:Y�腰�֠��C��RDK��.3���@e�d�'3�� @Y#�u ����d�sV�[BD@���α���r���I�;��5|����]څ��wl�+� �����6���M�����̋yzkՄ"�u~��}(�@���S��h�%��7�d�R�k;�@l׬�Xk��с
x��[���XG��;K �?�/���l�O�#h�ٽ����V��֨���i��GЗږ]� ����A&[�j g��CK���U� Z��[�ަ��e�!��G��-�bq��G���m���"t���'����*R�w�]![�Ƴ5�u���E4��A7C�F�AQ�,�U�+� lO��j6����]6��l����"�Z7rK���p_�U`�&ߠ�-y(���n��D�A]�lU�0�#�]�N��@��1��~�d�r���i�������3���qH�T�(�-�Qڡ'���a ��ӌ���A���ɕ�Di&�y�W���!)1�Q���򹬻�\i�Hh_����ۖIM��}������o�A&9l�S��D�G'�jR�6�$V��S5�����.�hb��	�af5!�r������ZIF���m�m���CD}-�J@l��
 �ڤ^�ߙ$Л�����^wJۖ�Z��ԉ�Dt�?�Ot!�@[~?�}p�����i=���lo�|FX	���v7}�cVEj�N��B���2��W5����9(r��nF�_ +��Eѷrn�=��J� i��)h�r��
�N+M�|�	$m��c���<6����,�����1'�r$ȸ2Z�q���y�(?E���d�g��9{���d���y�`���������$磉1�����<�����/���;;l�;G���(������6�����A������@��>����Q�M0�8�"t=�7޲J���^L��-dOa���݅�&6�y�Rؕv���Vx���gW��O�>x�;�h!޷C٠�15"H�6�QSI��(��<7_Ժn$�i�7�с,>o�w��q���Wj���J>*E�>d�
S�y��nG6ϥ�-u�|Ʒֹ���c@�DDmP���'�ml�H�K��.��#3{(ڼ�e�6�ň}4�f�����J�F�;�w���~�$�.C�AH��S��/���Z0������]1a(V��:ǌg0\H���uW�_Q����㭗
N�`��>B!��]��O�{&�,�^�Z�w� ��\��W�)����I��5w-��E�	1I]
�2&=Ŷ�e�~�[v�L�{_�(][�Rڪ�V�b��=ſ��	��.��փ����O*?U���Sc��[������[�"�+}TKvc������d��j�	�3�F��Z�z��#yj�"����!ɛ@���ӈ�n 7�?.��+ @���mm��db[>W�K*] �+Ϲ�'A���)u�(	��ٖ=��t�~��҆GO��$�pp'��Q>t:�~���{~n�T�iF3��⼴kM��P�?�a.^g�@�]"8b���-��]��V��F�\%+LS��lF��ܤ����0_[W�6�W|���]p��i�+;b���5��QFv�D���	��_�%���m p���䆋���y[*AC� 	��P�,j�L��}d������O3S�	pj:f!��\q�&N�� *�i��Ր�6\�����m_S���.֚��#a�G�x �m�BQ�1�c��x�Nߋ��WjU� �P��Vz��p}	�$u[�ӯ�g�c
)c��
��h�m��Ĳ�8�:3E9kG�J����e�L�ɯ=~g���D�`�[`
�e��?) 6nkA��$Q%� `{6���l�?Zo2��p�=Q�޹c�n��-q;
���O��Ȕֲu]��o��gmaS0g��!��Z��RQ2�ju������X
dJ�4)L��:w4SOm�1�V��ss�Ϋ�����5�1�4�L��1gJ�:w�U?P���M��h8�����ζe�)�A�p.9g��^֎N��-e�����=�e���Hz�1�Zj׮'� H�WZ��5cu�{�'�r��>v��5͈�Gc�mb�/u�� .<̲)�8���N�|�2�˼*0����3�s�2�eR�١��:q�wG��l��Tܝ7l�q7R��tﻉ<`h�ѣ��.]���v{X ݅�IW9�0�ziȣ�p�jUQ&���
EQ?V����<�NnP��1G�-ch���4�n�'�]4۱	�<ě��o���L�'�L�;�$�XtQ�id`V�%H3U�e�`�ֺD��,"S��݀�7sR�I��~��H��\�(G&�wJo�ͳN��~�xB�4A���$���.2~]Ƙ�ܬ��PE�͛Z���pE0��~�ԈC��"��N��hA{�9�[^�7�,j=&V7_V;(*�ukM/}+&J?��7�tt�;��Vj�j"G��}�9�5�]ơ,2�#_D���k*~ƕD�ymÎ��~Oe�X�(�";NP!�\�V�P��m��PR��]�VG똯�iL2��S�)��/f�t龢V���C��1�iT�����x���35�F�Щ�S�D4犇M\7{9ρ���v����ώ���h�:�] �<�fL���v�g1�{$k���P�����3D!1 �/Ц`��ṈM̮��>Y[�jpXt#o}�Vf_���ސ�
ه�T�T߉/c�/���j�|<��;Ф�s8E�)KȀP�-���h������7;t߻��G�o&ެ�L�FA&������:֌6tJ��l�v�w�K��.b��S�5�ؘ�o�w�dܽ�b�p�3�ox�jp��y3h.G ����x�d���X7&�4�X���P�z٦lLsZ�{�_���������'�ӷbZ�Kڬ�9����U"��8N�=z?0a�f��n�K/���x��p�@������Q�wB!���k�^V�o�>��S��K$v�`�0���פ��Y1�"c?B���]�L�P�w�P�'��	�q!�e
�V"��ZԬwi�5���E��D+�#��PS�h-�QY�g
JGO�����
7?���ݷ��:n_)0a�|Q"���@ �EEn0,�%>`15�ʍ̚SP�᪛�|
�g�^j��A�B�g��ˬ,�:���f�@�+����Iʡq���Cq��sU����i������-�u΂=����Ϥ��O�3�}-z�\�G�'��d�* 1~ ����@�O6w���xݺ0���@��$sL��nnzv�~Zn�����r홥m��VA&�`Ǉ
?�E�jۆd_��ǜ�}�Sb��/�0Jcv@���MrGȄ�{]@l��[�^��K���=���q~Q��o��Q�2�EX �T�4AO5�I�;�o�!����փG��^ f�m)��}��b]�pj|M3�8k�^-��PܒJ�$߶�uq��G�5�:v˷�v�(urHY��~�";���Чƒo	�,ӿ�/ދ��{��2�f'g�uz��� �q��K���JG?ě�������ՑϻL��S�8���K�B,��&���$��BZ�z.��(��6s��f����z#� t�>Z�8�hc�3R��! t��96�m�@�T� �1����.�$h�&����>y
v: gG:!�G��/��dmf�9��-A�hl�����X#/:���9((|��o�]2C VnQ��CV��˶���5���b:#��.�k��@Z7��:�d �@������=&^�X`Yk�F�G�ٺ� >t�R�6�JP��,��h�v��N+tL7�ݛ���9�BG_��U�MV�@���Ą��Rܲ��4�mچ�n�t�H]?c|`o�87���˖hV
8�0�E�;Ϩ5G:�2� 
��W~|�P��U�I Oɠ��h`�I��֘�P����
�j�G7�?�'r�퇢����Ժ�l�El��u瑝yPT��9nDc�;!]t? ��X]�ٖ�@�D��O
�p*����&0�r����h.��v|��E�,0V9�FOt#ag�s�3�qh���F�߽�z�B�9�s��3���׉������>2ȍ?u���n4S!�6���S��|����h+�����n�)�Z=�J��
ȧ�����,����3�G7&,����7P�M���8�o��徦	�S¡�Ѝ	e��v�f�-���V��Rq��� �B��U�L�*j��B�U˃"9�	����`ޥ)���4��N��:9n��R�	��e��՟������_κj�qHݿ��z���rE,�w��y�& U�[���o/>�o=�..V�X:��F��¨�{ǒ>�kc��6�*�4���������!9pq�1��n�9AE�+"ܐ��>����;���\�$�����0O�dd�V���s��u�7�Ս�e�l�5�f�S�>�Q���;�9F�m�K������ ��~�I��Ɇ��r䛧vk�'��z�$�N��q1du��es�Y/����@��AJ��n��u�=!1"r�\i��tx�@�ɾW�g��@4ÍH7��}C7]tjg���S�{���u�_in��pO�X�vf>�)qs;mFl�IGߝ7b ���nn�֏I�:�)���5_�8=�M�]r����6i�qn.o$F�ƣ���`���`���_��rm���Q��({<�|�.U~��
\c?��L@��N��<�[_c���uU�H���/���୾�	�4��"��۴��k��Df�u��A�1.�q����.?v��\������o���9�� ��Y�[�Ɲ����M�M;ͻ�{�c	 3�}�Ô�Q�,ǔ�0q�܎���as,l��Y|-�3�D%.�fQ+Lm2�%��6sx=�.���Z�����y?ḍ��r˶~}����:J�	�m�]���t�8zX�7Z,�L~^�^� ��R:�N����7e�����%�"2�[�#69�׋�(�/���ё��NFk��v�l�_�9$R�y�kP�S�7�n&�΋�Th��b�ʎhj��~�S) �����9F}\_��ȸ\y�X�{��]v.�~�r� �r	��y��4�������sz]�J�u%3�	�/�[��Bwӵ�N�LX+�M�gw�T��<b�,�:d�c$��TkA�����Cc[�����́R�-�ڞ����(>t��
<�su�4��7f���0��˂ֺ���vc��
u0�����^#������׊��V�P��e�m�ӥ�{�S�v�蛏R�c�T��q2����#�6�*R H���i�{F�Z�?}S�Mf�$��C��j�]+9w�J����{�䄈�Ǣbvşn<�nZPsI�&oe/1&m�U�J��1r�U�UA.)���qf?�7
�y��3B�VuJaQN�r�݈�O�1mX\��R=��7���0G���^�>���ѡ���bU@e�$�E[uNҭ;�ܪ��˃�_�5V����Z�Tia�O'W�۠D�IWeS�����[�Qk�*�ˑ��s�W�HXk��T���WNU4��N��K$|��{�ĝ�5�u݌='qIۈ�0���`[�^��}$^r��@æ�,�7��V͈����K5҆��l@�#Ɔn `[��9�}��Ǎ�0ԑ��>}���;�07Sn0m�C[���=�����['��͵ΐߵxMs�`��J˼T�)fe^񄃅+���I;�ze��!���#@<������3t���H8�(q,�� �'*������u�عs���Ε<��P���Q�vKH���v|���ɩ�S'�	_cٳ\�냅��2��������C�N��'�ʙ;��w^� P�I�e���%����5�m�����0?-�D����,0�&P��U�%.#֭]��;��T	ߠĢ]�ޘ���o*�*U��K��6R�)������	RZ��Q�و��Ib�Bڈ��D،��-^��l���#�@7���og� ��	�g���s*"x����dÕ���m5�	���ﴯ`#�������B,d�tlWj�:ȹ��=���p�s�W���+L3��
�p�������X��O*_͘,!Y��nB�\C�2,�C2� �NH���M�M!o�]Zm��WW��2w&~O�X}�HNO��~9<���F��6hxB&$�z�Ǧ	�� �ۊU��m��k�7���18�}���A�W �ɼ��H���-J�.��ܫKJK�x�+TH�1���i^��ڹ�&��F����ޜ����C@ش��S���m�R�ѥ���z�!�eL�������6��8�k*�n� "Fi�a�8.mm��(�E��Z����؆�Y_���4���:	^>���%��dr�@�ˎ�1� +�L��$[�3�K�@�H�5i������S�{����+[W�mG�#�IXSzz�B	N^����5�]GPY���.�\�79���@�6$��b���7b��+��@G/piK�����J��+��ۓK��![4�1S|b~��M��ro�:ʛr���A����{?����H��8iPd�93���[��ԵB�J*��y�`�CM�/���/SJ��peo�?P�Ԋ����6wt���?�
�z�8z4��r*o��C.5�>qcH(���<�ZP�wwi�E.�m�w��,s�
a	�����9o.-~��>rM��a��rU �^�`ܣ1�?�(�?���
'{k��c��jm��G�[������\q���O4�dL}o��H	�
�W<ߒ&sf�l���4�,_rv9	8���
��������D��Jֺ���Z��a�PK   �X�XA��5�)  �)  /   images/f5d8cbe5-36a4-4687-b22e-186957e3c304.png�);։PNG

   IHDR   d   O   �`�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  )QIDATx��]t�նޙ̤��� Ҥ7iR�\Q�k�+z��U�U�\A���PDD��H/�$$�RI%�N������Of&�0���z�u������9��%�a�����sY�e<�b.p�V����EY���sY�e$�B.���N��VpY��y.N\�qy�K���U\>����o��%���Z��1 �����^\��r���g� �ɳIBޟ�l�U./��F?�p�a�ٷ��3�}��\�� �*���Fb��3Ԕ wS#1dp��4�� xw����O;.�&װz���T.�\���'Hee%����N�krρ���L<���$���s$0� {ߎ����H��4DEE�,ok���ԅ�����\b�����I���	��`/A��x�Ăl���R}UUUCppp���c; �� ���֞+//��.��&�n;��@�Fch�d��������c�qqqdq/�e�;���!V�\G3��g��] �"Q\"_�@���0�Hb�6�-	!I ��v��nk��wLL�>''G���M<+	D��P��H��F8͋cˑ�{w.X;_�@o��;r�7m�о��-((�;;;�����L �I2�I��&�s�� I�����D��#���ؾC��e��IRh���|�#�VF����EO�GJGG��C���i�t�B�1B\w4�7�0W�z�#�H6�F��I�p-ȽJ��@��2,2R����$rqv�!��2�u�-W��4��(8$����EC���J5���\֑�:1��5�s��xxW;��'%��`�K�����流ʚ�P��e�W���ess�D�E��m''%ujJJ��$�D�����Po֓�:�Z�$I�0�,�ӓ*۵�:���D����A�Tgn7�|:�v��è�^K
n�F��Ҳ�4|�Xrvv��e���3�	����ᩤ�6���	����U�m��P��ҁˇ�h� `#6C cG�ՓB�3�U��-ӭ�B�Hu�:��
F�D��� ��z�N,37���
!D�� �DЊ6D{$~��j�`�$��f`� =�:��\rI$i��2�������	RϿe�`�=�R}�zR�Kqs��2�UP��:�N�]]���nW�r���Z�6�tu"�R�I.1$-�~$� ˧>%I��0�h� ���lq�*��q9aq��\ܱ|+��:c�:n, �@'X���-䬘��|��Fg跻m�WQ��	a��l�`��R.sI�p��\ژ\���Ir������Z��$�XK�@�j�I��w�� �Md�2��;ݾ)�ŧy[�����v��\��d���.��K�� �(� {�1d�����C��(��Yb�{�;{�:1d8��'.�M��5;(A�`I�p+���Q.�Ē�	�4��-ףPج���6��M�=lC���A�`c��Rv �lh���EY�?|��01��� :t�M�5577�bbb�����OQQQV�0� *xBB�?^ԇ2~�x��A}�ڃ�����F�F�j�Z�9Xå�m��{�d��}������l�W٣�@]Ż2TWWۭ-����*7���� ���&@��׆*o��-��M���� �Ė�)�F�=,����k�{߷�ݙ$�ך�W�5���� ]I�$<���? �54-W��J%���Ю��B�;��Y�Y!55k��M�{��5m�z{�k���$�A$D��Z|9璯��o[fS����	�J�*���\���/�3��֬r{�t\�p� �8��$�f"`<Ol���;��˛�YQYG*�`^���� X7o**Q�J�'�ʅ�����JE.��L�æ��Ⱦ��ܶ �Dtt/JKK��
tL���@
		����PZ#k�(+hg����q��V��8q"]�r��^�js�v�ot{jLg�/SNn�ðA8�Z��*���_͍�筷�"D$~�a�qcAzv����N��A����E?QU�-���?�ի�iӆ:t�@��ϧe˖���]	�#'g%���y����_J��Z귣={��۷/���
�+d�ƍ�8���ƍ�����=��p���La�t��E��/!{�5,ﴖ����s���$�mk��777���ڵk@�~�-u��]ԃ{_}��`iM�$;��������<]��䦖��X�������צ��,b�ݺu3�Nul��a	x��G�� (P�o6�e�ݩS'cp��ϯ��&M�D3g�+���_��c�����o
��A�p�,Y��j=vu�Fk1dA��й���I#��$3�^@@���g�@0������ܹ3M�<Y<B���Sbb"͙3����O1}�焐��ש��:w��yY2�@�Md�®�^T�R%l���8��*]�Xޗg�Y<�䷌D��\P�\���R-;B�C�����Q�N�p���eX�b� ���K;v4�l�-<7k�,��Ƞ^x�.\��,�nA�8ZQQ!:�e�Y Ǟ!�G��ŉB����k)=��S#� L�����'�ii��}ԍA�999Զm[�{�:kkk�(//mBp�5�5�7��	���B�;tD/�ˤ�WŻ Th�?��՛�URU�:�G%��]u��E���b�x�!x�e8r�M�6�ƌC���pL�����B'N�,����oAЁ��:{6��hO}z%]�;-�[B��z�R�
\2�r��ѱ�g(>1]��ŋQ=��߿�._�lV��!��MKAm�RmU!=3w6?�"�9;;ҷ_.�acd�h��w�ҥK���ʕ+i��ʹt�RJII�`�	.{Ȍ��h�|:*�~1[�����ӧK��M�8�~h!)�nt��1Z��Zʺ^"&ÂD�PgG�!�	��h
�W8�V����Eϟ�G ʚ5k����>�t��������i��)T�Ճ��.�^~�~4+�qJ�s���L�kf���G��cǊ�H�ۿ�ڸ�s���� ���F ">���S�g
2{K��Y�n�̲��y���u�lG����⺃Vd��{�?]BӦN���ѣb�!EՔZV0 44Tx.01�x���N#G���[��GP�_��贤�O�R�A���kZ����A�z�"�� <�JJNNA"��g�T��{�#++�~��G�B�j׮]"�Ԓp�=�����+X�Ē��_�o��*���W��<=h���`�`Y-�E��8u�?~\L&�4���Y�`�a������-G��t"ogһJ3']�N��M���}=_H\.r�|��u#[u0�:b���믴g�7n��K�MV�!��%ؓ0�z���4�j8p }���6�l�� ��~���kb5@��۷��☛�!����'�vf�y�p�;hn���dU�&~���꣜�.����2����ڿe0�'�m �;�
�����U~������j6�����M&�tݲ6MDX �y��
��0�Q�O?n=B.e[�;4,�u�A���lLï�
�^�ӧO� ��z��)�{zzұc�n[�Жd�\+X�!v_A.�F^5�ܺt�1û��N#8�p?}��~��-�eb`Sҭ�A$q�>n���D)�Qa�)��cǎ��f��44a`���90����I��m�￷��~��V�!l��ׯ[��W_c��{�G̼��2UA׳/S\B�N�|S������Q�ߟ�|u)I[�� cIʭ
�+�|5����n�������l�N`
2A�����#�-�as 	�(�I�΋\��[�� 8l�[a�V+z���Q�o�7 ��c��Jw�+���� <ɥAи� +��2�
ֲy50�dC�9��$[��A���j�K�����	����=l�K����������z�(KZ��:*cE��h�L�;��,��$g�o-hr �������BEA!`�Mb$�A�P�+�z-��\�l���)Ҝ�m��ZLqtTR���t��q� `����޸F��6��um���%Y!�[���J8�#��u�ņqJ����(9~��� ����^L�5q�:4����D�jO�E�7>/_A'��?�v�9d�#��˝�;PWW#f8�W���U����*�j)>��BQ(.i�U|�/���{�p��gJJV�3�<#�n�^�\K��� RRR)�� ���t�4Z)a��Ƙ� �����U�5TUY��1��r���6�]\�TT2����=�p!U�b���z�[ ���!K�����Ud�|�:yР��Ot��e���TY^@�%y�d�oTX$����B�l�.�p��ܝ������~���KƝ4S�C�hQ����pYd���~�q�����D��m�饿��ޮ/yy���DG�6�R��e��%X8�1��㏉v��{f�Z����,�(ْP����5,Lz��i.i�Z�2r����X�T��3��*J�r�t���3M=�4�j�Km"���JK�GO���TU[A�Ǐ��ԓ��։�b�Ӯ��6���d#�V�@ o/w�T���+LK5ubśz�m����SJJzuAR�� ub��g)GK�>��:bg}[�R��@rr2�5�ut����� /�bSځ|��E�g� �*SS����w�"�<��C5�ר�����)nu'Tk�z^1���f�&����E����+.�#Ȱ_�#>ƈ��bd��y��<��M��ꩩ�&7���4�UT��2���Cc����LC���JU��t��ڀ|� �Q�i��w��^B�P���s`m���J��2��l�X��1�qŪV��v�ډqDx�� !��)�j"����k���Pq,�3�<�܅b���P�C�δ���Y�GE���-�m�f Y3�E^��)rҳnP@@��BЯ�]�-�+!$ȗ톩ԣ�D

��+EG��u��/��س���AI���U�q����@��+q<K����{Ba�"�B��c�~/F�5��ɣzM��Oi�֏�Y���B�b��ŋ2
nP���]��Q�B���WPF�L|Gb���E<㇌��M�L~�yy��Ҝ�O����P]M%���o��*�5��ʃ��/�Ȅ���v-�,��hhPq�I:��,��ȾÕj*�������|a�>��O�v���%Hvv�p5�`q<X��F�d�Yi7/�x'��M�CnXVј`G�]�R,��A�	%Fz2yh�Dt��XNl�wh�o�SP�+e�<B#��Y�� �M����Ӽ���@��}�O��"�Q��%��+ �oVR��4vs:�N�<)x8���?�<����eѩ�4� L����MW�D =!�(]��c-��^?���1(/�PX���
����&O�`�#<E��ʵ<�eB�:uR�ֶ�����L�dX7��á2Fґ�X!H2�����߸�ɾ�A"��𪇇�в��f^=C�����0A�ЯM�ԟ�5��F��J��I�&R�6j�r�%�Ϣںz1{�!t�]-F���5���+�"�߉k���c\²`��[#q_'˛���R�>($��0���p�=A:���J�o~�-���!/�^���s�+�&``�������׋|}��خ��,I����8:|,�&O-���
��][˶�W_Ӟ�۩�����C���Ơ[ D���`�8$�Mnn>�����j��mx�
o�R�*h��GI��i�bե�f�
�!r��n߭�����	i
�S�3�9uJ|g�P��:����`ƥ�$�� Z�F�:�:-�X*���;av�x��sӄ-Խ�8���I����Dq�ɓ�N��;�^]K�]���.TT���ɆX�^��:u���(yPI���T?�[�e;D���Plg�������q��S��Wl�q�����d�6*(l�Y�F������#�o��F�����e�]�%�%�b��Jo-�(X֝ Y��� ��5�z
�������r���(w��0M�N��Č��/�q��{�^(��LQ��YM���N�C��z��ч�:4������hޞ%sҲ�ܮ��%$�����
���D�3��$�� >Y��{�\�1�\��J��TVZb�.�N@oT*��88 ��DH1GGqM�R���<9)��[ȉ�3�^�SC�9�Ú�s�k�I�"�uQB���c�0's��B��?�Ȭ��j�B�ԣ��-Ģ{u��C��?��V�F���<�/*�9���d�
�"�_t��u�;î М�����'��"g
�=��RjJUW�	�Oi����B�����̬LM�=6�~ٶ������֤p�r<f�|+�h&�"|(��=z�u��X~�)s�(��e3F����]X�����h��A̲�o�m�m�$��(Ғw
���{�˂����fKir���n�����&�۫�#}*�l�3�{y��jD���­o��\z�W��;v���p�(t[�P	D]�V�x�M��X�V�Ȳ���v�h۞�|�V�XM�T$�7^S2/�
t[`�>�q��ɀ�be�F��f���O�%%fKd@��ƊtU�FdV"���!C�>���04�<r{�Ǿ$��	��Νك�D�Ok ��ڡ���NM=�������v�`�� �cu0�E�vRue�8�M �dި'gWo���3��'4$lTA%N@h	�L@���E#�=I6��۷	¸����o�E�M�FW��҇K�Uf����!�h����h|B�1233i�ܹ�o�>�)�s�NJJJI�gϞ����ׯ_�	���^zILum)UVVQ~a����P]�O���$��]dx ��n ��qT-��� D���g�S4��!����м9��좡?����j�&bΚ�3���OZf+Z��l|�&�~��!2I�(8(��"�Def���/�b԰��Y�U�� �h�=�x����z��LB����
����ݛZ�qƔ�4c�`�mL��?��� ���ww��3�	�����T/H��!Y����l����"��G��t �����e�6r�p�%&]��G3f�0����8���`��J�4>�� ��ٳg�Wˋ/�(f)�� �
�V�gp�́h���b��ƀ�$�����[]ػW��#Ƅ��-�~?��K�3�cR(�,4[��)"y�w*-&�
���H;��"�[W'�Y�4rޖ���-o �u Y��~ ?�����{6����<�]w�'`r�Oɤ�A�a�����ht�����]Aj �)��@N�ڵk[��)o��e��5Hw���@�ĥ+9�r�-&�%>�'{40��=<�E��g�8�X�ŋ�M�?��
@��2�x<:ku��ٰ�Hږ��rr�O��Vhs�"A`|��Gb�ɩP�ţ䤔؊F�(���>[E{��/V��{0�'�`R��=A`��/����
�w�u�`U@���5��P�!s�����/$�a�ىsK����5>|8�8~����,U:��^˫�'������`2sZR��%4�o���2�/Ӂ�_Qt�(rwkg��F�*[1��q�?���������c��hy�Pm����&[ DV:��,��{�Ȇ֒�D���2e� |[�k�� ��f!k���/fܸ�/�WP����%*�17��Bմ����-�Z��K�7��f��,A@���t*�?KC�@��yu�v5/�Dn�I��0����1#z=����)�n۶md+ H�ƀcbN����էO_&D��� �uH;^�}��b�LiY9�޽�ڷo�"AD���CS��d@�yy��˫��ٰ��o��ׇN�B���D�9��^�J�מD�0�ӟ��!=;�%��=��j�'}��V�b� �-�k�k�j1��2�\RZ9��ϳnu�E6n��֪78;;�:�k��w�@O<�,#`�@�)t�І�t
�[|�U*��-����
��%��t-��.��7�G��t$_���O�2���}.+;�j�C��I��^��_Lg�.�ΊL�:ݻF��!�G�P��`9*U���Jw��@.�,��('��\2��g̤�?���C�bҞ������ũ@�� ��'+�j�sws�үo�	��陵ϧ7o��99����).�8����ZeU�\/O�:�>T�������_��Kz����`'�����:���#�|7M�8�R�k�=��W��%������<��	�m��@�L��M[��߸}����>*���z�A�;t�<}��qW��g���t!��"��3"Z�r�N�3�a��>���a<�U�C�N�0�닯w�mF�E��s'����:Y;�^�����`Bc=���մTj��j�C%s��N*e,q�'N��rg��*��x��'t��t.��L�B_~��6�t�ԙ�b�R���h����
,�+W���?�g>x�	�o�6$�g���`�q��D�G&�n��G�7>��q�����{"���ҬF������������^�Ќa�#D*'G̜:�:���jfn^IR�Ƞy���3��9�:t绻�jj�s���~�gw����I����x&4�W�ūauv�7x����xl~􁑃?��'�?Bg=8��zLIi�#55u%�A��U�"V��cv��y�:F�B�����z�s�P���?���돈ď���|�V�����I�R��et�Y�M�e+��5h�~�)��(.)7����㷯�Ӏ��%''ոښ

o<M�C�P�9�����ž>�5NΪ��͚�6��x5�Նl�~^�Kx��C��S�������� ��f	�yV�2Q��V�\�ł:w�,�K'��6!8��;����tD���ֱ}�Sr��F��������z{�U2�+�Ԛ��`�a?_O���׬tqQe�����	�tۨ`W� ^̲�y� ��"dQ�v!��_��.�L�ޟ�+��O�N��r�X��1u_֣�ņJ���(����}�2"l^zvQ�̎ث����'��.*'�i7'f��^H^P���* `�tTD3r��|(������Z��>�Z̏���h㲏�����Ľ��mҮ�yz�Ν�(��bK'��'����(=�J�lD��h���� ���p���������WS֧e�AxD\H���ף	�E�@>��0��f.�%�)	����K8�Xk����ymEe5-�h.�b���O������v�5�����;ҕ��SR�%�Sfv��g�O�j�׌�N*��GN$a
@"vl�e;���j�6�e���˼��4������C��)�%�[y����y>Qt��7&���Ȝ჻�	
���+c˺�?�`$?x$��L*[�Ȩ��5rO��|?������/2q���/�}���2ԗ'J>��y��SM6�ffe2B�>)"OO�1����E���z����3�?~F�їH���&�����/o����L�[޶�#���0ae^9H�;E������H\�����S\�jx��YJ;hF�Πo�mܐ�hߪ/w҃3�E��
Y�Uq�d
���Y����Wר]����ԝr1� @M��gRI��}ܨ>������rD<�ڟ�������~�r��3������.�/���B}h��c��f���k֧m;NR�Z�ba���R��ۏ� �ٚ�|O��DG�h���J�+l�BpI���ܜ�)�����U�L��I��Ϡ����	hv��%A�ضgϞ�|r��8PxX��<SB����O/(,f��?�ΪY9���]�e�����=��M3�6�^��=1�c9������@��0,����DBa��6��7���v��~���+�I��c�i������J�+q�[���/�I�����P�b8Y&y)�e<}TV^A�j/n�]8=�p1�5��T��>�������Bڰn�������ҽΈHe��ĳ�y��Ff�9�����?F́-�qy�TK 6GS���:�b���|�w�+���׈��&�m�ϰ��6���k7&hxQQ	��XB��L���|��˸^e�FiB~ �\�nٲ���+�Ҟ]?�D�m|��Qؗ�Y��WAm�i3��K�_4�M.�����q��t [ .�����vP䓂���9�Wº�$����a��?_�O-�cG���GD�w���[0Ԫ*�G9ye��۞����?�E����&ۉ��!��w�����p��q0����QYy�ذB}�⁜�Y�>bvX=�>8����@$Ykǣ��7N���"[Cx!P�?!�d��"���S��آϠ��B�HC�H����l�ʟ��$|az&�<�g�Г������T��������CCۈ4��1���М�Ȃ'3���Pjk �(X!Hh@���0�[:�`�9sF8�bQ��b+� ���o����#""�hB
~��<��^abi������^��(>������S,ozt4b$H��M�U&��[���,D�Nt��֜`}萴�[>�P�~� 8e t��P+71.�0.[n��K&�����    IEND�B`�PK   $��XK숤u  �x  /   images/f8feb36c-29ce-4e87-9091-184ea2b3473b.jpg��eP@%:8,0������:�n��[p� ����;�-�m����j�ի��n��u�G�����Tu�-�m��HHK ��� ��m�� ���/�u$T$$DD�w((Ȩ�00�ߡ�cb�����BGO��>>>6!.>¿�HhHHhx��x����	�A�#�3F�����!������ pHp�5 �W����2
*�;�� x8xD����_��_������M��7C*<v��Tj��.|��#� �w�D�$�hh?��sprq��򉊉KHJI˨���k|��26153���rrvqu��{�
	�O����������_PXT\RZS[�ohlj����������_X\Z������?�sxtyu�������� �����?>����(�����$"�G6d\�o(����Q�D�r��Ш�(_�9N�# ql}�������P����F��y[` ��[0��E%7�3���p<����%�B���[a.����@:�)��t4y�\u��r�ƅ�i��<�f������\�����C����	��������/6v|��i�����%gΪ�<����]彩Ց���������Nr�P(�~O��1I~vs��jԵ �8J�_�B�y!س��_���[u��#F6$4�!���e0�� �4iN�6�\�ۢ��fTT@���T�L�fw��C�,;'�����S?������wd���;d�b�l�klI��*O�
�d���7 X��
���|�A��CM�}���G�H�k�|�&��^�N�~�}e��[�_��t�K��"�	��0N���Ss�x1>�#f6�}jd 0����r�𔏼�p�c(5�k��NJ �rh�Q���8����,�x���J������O(�����F���C�Z��Oc�s��em����R'��p�C.`��i}�ZG�����'�L�e��� �{��M�bmb���nU�����B>$������Xc|w'�W�)�:�2��[z)�D��|�ZS����Q-���o���U�������:��zri�iٟڍL�Prex�y�c�t*�Ҝ�Y��	{���6>��������͋m�2c��ja(���7q�yJl�m��� ����?�F�d-�������Vʹ)��qjqGq�|��Kr\Q!���T~:����ˤG<���{�%���/�^[�$P*lQ�p�炘c6��"\�C�Q� �m�P�	L1�cp�i�>>0�\�˿��0�K	�2�1A�~���ܞ�\=sVI��!w!�슬����-Ȩ72��@��j]�m�&�x!gu�|��cb�kJ�|��0B\��fZs��K��	�IB�o\�J�5�*f�H�E�}�{�w7t�lS5		��R�����޴����d�/����A� Dv�D?��A,�����U�ٚ���ś%E��`����N�åŔ~��AD�+�V��˼i��G(u͒�f�ӡ�f0�UCts�6��h:_K�y�\�^�+q�E��/x����#c���)ψ��������]l#�q�ʡ�����~C�u������W����Z���j�8B�/�MR��q����V�
]���!���%+�����)m��¨��j3|ʽUx3�X8��C}l ��R$��6�����{%6�Nb�Aa}A���Os�C���`B-V ϫ T;�p�w�s?`��=ݙ�Y��>ю�w�x���\l�Q��-�h2d��m�[�2^A��y�G�6�qz�I[>(`��d���e���� �Q�PFTɠ�p�Y��28�19Ӭ�F�a�(�}wR'�iv�@(�P?<���.����B��a�d��4E��/2�:@rP-��h�:�G��#2M�L�r[�[�ٮa0[�-�8ҹ*��g����]�����s��|8 Qb�L/��<pH�;j��j�-�4��/�YlyY ۴FZˁK����H���J^$;#:�k�m��%`�z�N�B��_�?v��c
A8.����T'��;`��T@O�zL
՟���J1-�k��·U�Qw��i������Pe�3B)�J�����d�;!H�3�"7�7DVIi�K�-�j
�� �8j)��5���^*�)v���s�=��x܊OɴB�
<�w~��6�ڴi�(��� u�b�7q ���E5�*���_���D�F>v��.Gݴ��
��N��tG^�R#�)�K��¿8?E{Q���l�-7#m�D��T4g ��̎��c�fۇ���3w�[��į�N=E�Lp[]In6��3Aێ�0R_g�T;r��a�{��<i�_�lBŖJ��	����s�G���&���C�2bZl�a�4�ԃr�E��%�n��oj��ncj�� ��/o������3�5A��1��}Ɗ���D�E��j�zE��� 
h����c���� �+���i�@�U��a�=�Gc�I���Da��;��Sހq�fW���	����m����({28����:D����Y(�ʢ�����l��K����o���T2��]�F@��=���9%P����,��G��8?bQV�>Ʌޱ*M�q�W��}����Zd�����p������\mj��&c_Zc�!-�p=o���]q\sSk����df<7sA��f����ŧ�e�氳e�<.ܭǬi�l��	Ŷ��(�i�EB~ȡ<��չ�A�:�ӫ�2mm��/�۽��H�h�fL�+��7�E>����  ��+��
S.�L���d�dF�q���O�l�Y��C䛿6�q���nϱ����+�g9�q�n�	Sm(A�޿�G���y��Zis 5�c[L��8/r>�u�Fv�8������q�����,�Bu� ءd�|��f�7v^���\镭����W&��~��(J3	k����Q��~�O .��e|)+�X�8��
y���S������@=����,{4+�i�X��ɤͶ`�S������*�&�f-/ŗ]t�6��\��O9k�I�6�(P�����{֩���
+�%��X�L�̜�֘����A�J����(�L�Gi��S�>�S��Bf�/+l9�ڻ��;���� �t�-Y&�*�Ǌ�����Ȉ�5�a���1�8��n	�ȚнL �6�7/U2Si�D��gL�S�����4�a��S�z��n�Ӷ�"��M����r��kJ����7��uf޼�oW8$/ߌeLo��o�|6^L����.���� ���M�Cr%Fo_Z�Ej�UT}��5�R;�^wX�]��ne��O3��@-�|��ޚ�h��9�8B�-����(�b�k��㘑�����M�I:C��Wj��9�^���ޝI)�u�ݯFƕ��:�ͦ��ҽ���#f�Y���f��O�b�͉B�L��v���,�{w[F�[K͖V�M�"Wt�ӕ�R���m�!['sk�7dl.�|&lږ���e�j�I"�g<K����C�|y�`OUŒ{��#�b�F�tawk����q�;�]0F-�A�c�ZtG�\v�~��/��m�-�3���5�g�d;ʗM~'�sƠfE�v���ߦ��|[v!���u��S#U�����Ȼ�v�Oٶ}C�;9l_�c�����~d��#K�Vb���^S�ć?$o	�Vm��,�ǳ�KVq휾�U�rHy�E�����˂#�E��%%T�)

̋Q�D�!���m��]zf���ͺ��sL3~�Jr'���ʟ^����ZYBBg�ʣ�PB�2~����Hxx%�ܿrN�8?C�1��rv�W�g��6J>�x��ߡ;��Kc�цԉ=$�g��2{���z��S{�57M�Y\ʗ�v�e��+��ԏ���g�J�ER&�T�_$	"\o�3ْ\���hz��\!s�c�)�0��@P����9󭴕c� �м��Ǩf�T*Q�/�ev������-��I����4���r	rR$ȟ\�`��eq������_{�Qh/�����WTb��FĊk���LM��mw�Eg$��SE�{в�t�]�P��H-Fs&[�i����͌�]����z��,F��sk�,��ɷHW{�pj������	��dǲJ��P\�j��<\��(��v&W�v�ļEy�i�H�
{��l:>��z.�a&�b$�i���س��RG֫:j^�м�:��׊4��5���oj`#{�ճ�ה��oG|�æ�������-�p=�
s#b�k�P���_�v.�?�g�o�%�H��/��|FW�H�� �;J[+�+������V��p��K���䣣��e*~��2���R��M��'�#����ȋC%PO���'l�}ٯ[
�o �������'.�_�\��g�Q`����gyR��>�K6 r��G�J�W  �	9,_�D�*y���9��� |�����
3�g` }���k�pw�����HS|w|9v��t~*A�Z����wh�xM�?�R�%ט�|��>|��$�f^�B�c��B�^b��%�r9�뢠Oיr	U����ͯ�T�(����+6�A%e���C��a����	ko�v��{�RX�&[�G��J�QG��񋼐�N꨺�h�_�;�b(8�V���4~��z���zC��j���O�]~U����Uz:�m+��H�X���S=�뉰qc����uU��/6�E*� �Y9�t�r�D`�/R���=��5k��v��;���$H��}E=��Ys�X+c�v��+��^[PM���J��%�vD�!��Չb(�Z�}/B,���[po�����9�
"��i.�Ӈ>B\_�%��1f����\�݌���H�O�s���"\'$9��I�:Ps5>�?.qΙFR�_���ى��,11cz 1_L��d�e;�$�-���9�1dDu��5.6���7�h��ȶ��"{���c��OG�F�>1��� ��4j!�h�dMj�ɨ:ϰ}ʆ*��u��?Rz5�!�������u4�/~�1s;�Z���=Q���޳A�N�Ā�+6�~w}_A�{�o5�|?��q��B�6|�|�?�/klƤ*�f��g��R��m��yA,�*&w��-����s��u��L��-�����:0�9�����\�꒗��ќ,8�:���y��!��p�d.����Qpu~c�9)���<%`���#�e��?wN��,��xTq���b_��RD�G���]�i�9yG�E!=���Zp#�fM�{����g�C�C[vhӉ.�v�n�F��<��k:�-쁍^�Ȋ^Fy���܌V䔳��@l�Cs�$��#�
��N\�n�G�N�Wb�dX3q+Ks!��D��/m� �eMfz_��5�(UG]���1���[to��`��'	�3�6w<~ c ]ldUlά92��3�6��a�@Om�������m��/Ⱦ�׊���jI�݋o�lye�p����`��$]�5��>�t�:D����N46�s�{c��W.�tҥ����5��������\��(m����O2�o�<�V G��K�=�l���'�%��"�����xyAS�H�� wn��_
^%l�p� �\f��/=�OSfSiIǴ�+y�������URJw����������;�D�q�iS�S�^K��m��x����8;ZU��v�zo���t���0��a�G��D�[��.d!��y޳<��,�n��$�Ք�j� 7�ڐ}{��
�Ⱦ�����ڴ�Z��F�g�t��	w��Q�Hx�ſ�k@�#��`@o�iu�&B�n�L� 5J�0JNy�͔<f�M�߻Ϲ��x��"WM����H�\����%�x��R@���~o����/��g\,���hf6����R|Đ�f8�.���E��b#���sμ�=ƶC�ԑ�c����8E��Գ�5/c�\EU�p��tCò�΀��׮%lc��}E����fV�=�9�(�{KX�{��0H�m7I?�-�8��L�s��j�j���{ �sX�S�8�e�k(��˞-��+q>����d�� 7�֯SW��qPsC�؜�>���.^��1��Ep��3)+���!A�u��gn2�BG@��}��g��������߭��g�D�߲
m�V��3�X}���ѻ�Y��=�����$�5@�����(E2�E{%��m	�.�u�D���_iC��� �g�ޜ��:�H�n};ǴyS������D�k6[���'Ix뤓���e�<K+�٢Yj��RI�F�J����O�\�}��#,����y0oъ%�Y6�MHl��@�ן�$�@E7k�X�kŨI�k<���ZR�����E]��ӿ+M���8wdޯ��V?+��bQ�p�ٽ0�0��Y��j,��� 
��~�5��p�Z� ,1�q����L��N�zm��c_3�Ě��a����y�*vz�K�X�	�;�Y�_i�Mq�%l#�+�q�x�?�g���6Qv��� �$�֗�O�hi��M��djCdFVӶ(�4v����枆!ޒR�"6��_$Rx_f"����jl�,UsdR�)k�����C����������JjIaڟ_c7�a!��MU���z�\�}��'�_A!�r)�RD1�����/n�ZC���0o��k�������/��(�8,�H6��A�!a�!����,��
%�g7�0��y�y��7�?7�2IZd/mk��kz�[&�4���g�ߝL ��"[X�8����������M��5��Ҁ�h� `'���Y��0IL���aܨ�ӓ����Q����'�L�&�L��g��m��ì�6���h�C@���F!_�<RCy:�]�Ȧ�J5���_S����4to��f���k��{�C�4��O�?W���"�P�p���Id35mab�����;��UE����ݭ �^�^y��Mb����>F�3�ïJ���9���-��5+�P~ %?�
����۫h����]}����̹W�a�ozP�9H[�7�9{ر�s�h~�=���yE�'e!.�C\��$��J������zXh<�Q�}I�Cj�:�݇�^���ޭ��y�@�w~���U�Kr�5AP��ܪ��2�x1����Q�쎮<(d$��k�St��I�����W!��!GR�_Dj �U��5L����/�w�lг��fĸ?���S�8�:�<��DV"L���U�@,,N;e%i�#Zr��`��������y�T�Lߥ�Bd� ا�ԭ����5�_|� �>�^!�\R��CK���:�����Xw����͓��;��Q��+~�1���]�+���U�2�2�[1X9G�q�J�%��%��!�l����³���ˋ�i3�ӈS�h>n���OW��l��rld��*J�E���f����n�9VJ���/ty�4�_A������1���U.�8�_ʧ�;4�@!F�H�VS�����Bc���J�&���F�0��y��QW��<S�	tg�_캫G�-�"I*��,ǒh��)��?��K�1�m+Zz����Z9�w��&A���v���}$��v���u�u��jI�����������tm)�;�Yu�˘��&�
#d�gCo�>�r�#�O�mb��\5i����Z'�����L*��W����;w�N�whCG-�r���$],T��^��ʇ\<}�����TW�m�7B�H?�WO&,+��B=�.�p۟����dg�L�>g�h�nq"� 4�ӳN��2V}1��;0�M�j��B��6����oL��lXiŷ|�'��t��lr=I [��1$%����q�W�KR�u�R1׫��iwҀ�v���TG�ǵf���%�Xz���ͪ·�":kZ�p֋�VK����JɻJG>dJ�J��K��3&�f%���;�$��?�"�.27�zB�R�.Mm7c�i*����>����M�� �U?X#q4�4�+��>:pه�u�9;�ƂQ�\����L����:5��VrV��(�����'�^E����q���i+Dz�Z{y5�ƩU�� �N[c�u6RD����}�H	tIAD���kkn �#$������7��{�7 \C��)b���$���e�Y�3Z������l'
a�CƊ�¦d�70�΄6��F����Շ6Ar�|sʲ������$�K�Cҡ�`�黜�uᚃ���1sn�`}���x�3�h�B<��r��)��ظPkA�b���|�3~���Oz@�T��8!�Y5�
푹������ ��M�R>1�D��Q9h���s[�>�P�]���YAx��m,+��G�7�^L��M���4�"�_�x2��Z��O鞤%������&}�^����?�k���.�
��_�_B�:��uT��V��[
�g�j-=t�k� �cO|�)�y(��b@�H��a���W�bh��}b90J���NE�QO����HYK#�i�x	-�^xF��":҄tfhY�rE~Q$�T�f?Y��7����\�����%Y�T-�Ū��՗���	�P�%������������J.��A[�è�}�t�qWq3z���Wأ�
̈��vH"��-��:�a7#��0;���2�`l���hZ8��z��T��ќK-�k��$Ϙ�)1�Q{�*��t���'����(U�!r�vW�=�#	3�IéE�j�ϲ�u�d$��fa���)/�Bi�[nU�m;Oܘ-�T��]��b����d�_���س��҆!�4Sr����g��GW��9L2��V����C��4���_�.�� ��k�+�ﻄ�+�*���j��য]@(��4XL��V���s{@�yi�G6�А��t�ԭ@��- ��}$� uRm��JV��	��)�*�`",��N���ˎY��Ҫ�����N�U!|F��� /�3"ME�^˃y�~M�j֩�Yf�Ɋ�f�-�2[WM����t�����;�8B��/ʃ�Ӛ,?��� =K�������aB`�o��A+�נ]��@�3v�y�\Z��@�o"غb����c
��+�F���h:�,��y��,W���J��=�6��R�vEe(8��@Sb�sӧgS��OĖoܯ*̾@�-�$��f��E]g�j�]�Բ�t՞-��q��ĉ;���p��E[�r{��M���oU �|���I����7@E�!�(<��۬��s����T�Y�Ʒz��W��%ĝ0ܯ����.�=�rY8��̅W�Z�W.�?Kփ)��\�b<�]3�ad�o=t�g�s �ga[c�߸^�G�������wê�ZDK:���VC`��{��縠���}����ؔ������4��pid���
Ia��Y����+�5a��2q��L��pN]��Leu���A�"lY�D$'	�I�����!�+��D\[�x��=���즂C�jY���~�Ǐumqj1�37���H^6?^��Y�g�������$�x��JԷT���������� ��,�t�,|��g��޻��j[�h���:~�R: '�����}@Ŀ�,�f���n�R��b�m�%���" �	�6��L�I.�j	�����a�
pD���%��|�#�N*�/E��C�hu�Q\W=ݏ6�L�2����1
���Z�'�rW�dk�]&�G;�8�������S��l����9�j1;4���(�{Wo�]���U̖��F�Y��q>d�~J HDD�[Kg̛�`���u]���ȏ�L�ۄֆ#r\�����a���Qb7S��g�h������`�&�VS�t�A�e/'D��z���
g���8t�.O�,9�t �XFA�c���*�˖��x���|jo*J����6�'��u�e/aFފ�����L?m�x��6�.~XYT[�[K�&�Hqs����9�6�ģ���WX�ȟp	p����%NC�U,]љ��e�T� ����,#cd�{���x��������ڲ�[���=�˫y��2l̂�h�q��z�>���z1��R�2W|+�m�Ȑ�j����B4RB%8�}��ԥY8e]9"'kd�W��kZE�뿬�s�}OY�:��m<����2r�ƞ�b%̒���B�.�f�Ȍ'�j��t�&��:<��_Ż�p�}z���N��ɵ�9����@`�'IJ��l��x��B�w'6�G�V���#��%���`p?#\��<����K�`�t��z���Q�ӱʆ�����}z`�e`��]��d� y�9hL]��w�<���d�E��$���Mۏ��suc�W߽���	����-�UG�h�'������Uw/
�����xpz�^�+��b֜?��H�ۺg�UP� ��"[`6�0�sƴ���]�V�8���㮼�̊kj��Ԓ(x��՚õlƪ�ta���W�����%��j�Xy��C�$_����p'��*^j-��ɑn~�|�x.��i�'z�%��uU����1���b(���O�1�C�V���B� Y��,�NGIͳ�d�=_�z��3;��q]�#m��[���]���ͫ�o6�'�8�H��q��ծv��e{�d�����}���n2�j#�����d�>KjpR�"B�A��q��b@^�^Hu�\�,Ѓ��^�G٩ނ��^Ҳ�[�&A�Å]O��P�WD��)Lq��GR�1Z}Қ�3=!� ?u��6,_�C\]DS�{����E%��#��]8�?@�ڙ,�).^�=�TS��՗7�>��:���ţ	��Nfkl%�ו��7��~��5�NU���A�$u�b��pA�~9�� C�蘫�W����(ؿz��1vw��JW�����8� &Kn��Kv��dW䓶��k[x��$�.^*��6[�B^	�*�=����N#��d!��Q�?�?�_��_�qZjp�y��wn�U�ah�5���[he�y���Ƽv��^���I�/B�XEc�q+e� ���v�-H0+&3�jj�ƽ�QN2قy�V2N�Z���εP(VQo�[%Mj�y��EQ9���%����*�|q�l�<���i�\*Ih�8D��chk�{�� �=f�Qd�~a�䮛K�.�uJ\�;�Au&�	���p����(r+� rj�������������B�v(��x6�K�1wh3��7Ib�%�i�cgu0�~����]��RK2�I_2�#1�ODY�V����d�Ð}�����.�0!�xYm��)d{��t�E���OU����t���i�b���c�m,=FT��<�p2�]��؈���JiSe%sL9ڜz��5��W=
��q�����L��c��84��إL�2R7�����e,AU+V�+{��{�!<`#�q��}��J/�K�_����nM��F�JV$&^@���nA��%�>�r�"ӑ�B�a�3

�TW
���ߙd��,���Cd-��K�����s'�s����?B�S+
TR���B�F�Ǘ'Bz��Z�~��I�Ŝ�I���2�ɱ{�����S0�� �)�η�����1/�D�|�V���m(m�$�Je���*��v!��� �C
�S���E�L��uH�Wh#^	 B�6��7@l�t/�ֶNݣ[�Ia�Q�r��r�����^2��u8�Qq�<���Q,��gvE�w�4(����7��(K�ىە�8.ҵj�q!H��$?ze���9��]c�ctb��\�1����*��!��S(��R -)�R֫D�ω��8��A��v*)@-�g�XbG�EN����t~��^ܤ�A�Vp�8]�Քy{R���3�2,��o��^㛤�~UP%�-�:]�@v�*��~w��v��J2�8	����3^����E��=]Y��Y�_H��ࢤU�d��ԺL�n���;{9E�'�FX���`���b�W�8JF��,����Ґ��b�����*n�7
"//*�}7~z�E*��Y�2.O��v�c��	u�э��ڐYh�j�ke���ݱRX�B=b�Q9��K��ȿ��0X#+R�Vɡ]9ǘW����߄~�׬���k`ڒW�P#��ݪ`�������Y��U�m�gvo�����..��tC�=�Vy6:X������-6��d��D��.Kqٷv�$���I(�n/�sɨ������9�,ձ���ך�����gX��򷍡OP0��"-�H���.�DjK �HfīJ_p��ڀ���8��>c_t���&��%δ�Űi� ��!e3��50���5�����5u�Ne��n��	��C��#z��V����u������W��ϔ�)�����8�B[?��tC=��կ��%��?)+�c��G�f�;��Z�}\ĭ�6�.^�/�j�#��m��7�ޚ�M��`qU��(]�E�����R�5�瑋��k�؞��ɋ��_g��d�Ar�s��,b�=,�Mk���Pv�%��v1�Ĥ�%�a�AU/�f�V�8S�z�O���s��Y����8x�缭����DsqV81��_c�����M)AD��"m>���y�t��9�K/3�R4_�L+�܃k-�D����vY���I5�t)O������ڲ��R���i
 ��E�F�������i��Jf���bܭ�I������e
���q�݄W}o��-|I�Z7R0üH���I���ϟ SuD��Di`�4��l[�%�$��n��zg��.$�J ����p3n#0S�sv}\��\]��4��\��A�'m_�X%�.����@��,�cs��@m�vg��aQC�r�4\���+1t�Jm��D5̃\<�S&ﳧҷ���ƀ�$�nG���/�9��^������I[u*i��EaMR)Aҁ�y�jx������^�����~��a�����k�-�?G�Æ9��n�q��)�>��/P8���zI��.].��W�Z0ݠ����ֱ�a�Frs`U�9B��ȫA��I*�p_K��c6��{�(����c������&8�}��T�������M��Mⲩ��f��7*�\V�V�bYZ��~C�r�۳�9\�D�럅O_�㄁=� ��ga��#�b�(Z���Y`c��[�1D��Gu���i�@�ƎiJ���1Ϙ���{[��E�wo�8T�Z�<�����.�B�J�5c�Կo�H�eR����|9��.��h<D�_���6Z����궬�:�fG��B��D�aܭ��0�sk=�i}���&�1��aJ��+vc˥I���K��Wg��!'��� #,��p%!�g��\/�����(�Y&�E�L?���途�W�Ɗ��<�H���6��Хm���a L)��*�0;�%䯞��ﹷ�H���?H����MP�%��$��� Q:Pԙ���hQ_*W�O���ۮ�6�U��3�r��ݏ]�l������ܷI���D��E��+p�'.|����MU���7��ھ���Xy;V�h�s��}`����հ�^a8�N�d��l�G���A���y�" �q ��I#-�w���p�p2������T�jG��%粙t~�Y�j̡S�K�W��7@M�Ɂ�f�F��\���&e��@b��e4֗:_l���"��F��CYq����u�<%F�O\���e�ۈ�����:`P�~���+Bm ��E�x�	wt����Xf^�%�"9�ֵ�>�6�t�7̳x����"$lj�#�b���=�f=Lg�zo�����%=��,�?r����@vz��$�T(ђ9��HZ���l�$r�O�ItǶ�XWO��i>յ/Y�5»�C�_�A�a��s�G��xF��S� ��㕮��\4l�M�[b�ׂ#�`����76�'�@�v�]�+V�u���s������U�PZ{&��z�2��W��3b#٦!�Ez�7��v�$�g&�z�+^�y�)�ңn�ʼ�>J�8]�B��:�ҳ˜�~��$1��hͲD�!�����UK��`��(9������T����rk��d{<"��#�࢏�p%�p�ԧ�5 ���x�xeB��	=�_~2�R���`����X4;id��Q�#��H�
y�6��|1i��_#��/
���\qt�ֽ�����#�U���Z�(�
]9����"5��פ�K|��!"�[�w�ըx�{�ɫ��hM�%ǎQ�n�-�T��V?s����"��'*|p@���8�AP���֋�&�	���G���I߼Q�fz��`z⻨��׈��k�dl�K��s|I�sǏ�������é��e���Z��鍭ŃG!2�{f�N�$�y����h o�
��\�Y�����٫9R	D����0�#9�
�aH��@�n֥��,NʹQaS�Ej�D�×GZ�p����H�w:��z���k�M�et5��}�!����F�ݜ�].dU'N�U�W��[tt3����`����SF�秪e����^�,�����M����$�O�*���+��6��S�T�����LK���9�{���+��2�z�[!4u�+��)ޑ¸�����&(�	��u�a<4>�e�Ϡm�ɔ�-=K�fu҃�Վ|�&���`�T/���O�W�:\q>{jZ�؉�nL�[�"���
�_�����µ�ړ/Ǔ|=����ڧ��L��W�	7��P�N9�DE�l�z�J��!���Gʠ�=h������)ةQZ��MUS�jv]�֕��}t�t��!1��71!f!ó�d%�n�4��I+�>DDDb���F� ���7���Y�º7B�}b{�k�l7e��\�%��x�}��o������K��%A�w���4�uR�ŷ�}4�H�:I�J����"���0��U�i[��B�Ȳ�
�~m�jn�M�1����̊�!G}���ˡv�{)�|	�K��%Q<�*���Bu�o
s����D7O�=�E_v�[�`��O�^z�j7~�_�h�x�J9�ѭ���Y��`WC��Z�lwպ��0����㐰��$jM�R��|��`:��{D&��@�w��A�,B@E����Օ�xM�3ƃ��k��5�p�(���?�v�9�нUěC9�ؙ��tb��M����>`�@v1�d��7=d���k-Te�������@�$ftZ��Ի$ǈ�$�{�q�p�6���>ס'�5̶���}�4$(��h���M�ݣຏ�Fo]#���"� �Z ʚ�w4!eC�n�Ny`m B���U ��p�9P^ƒ�g�M�tE��ٳ�9϶k�X��n�T��9��@��ܶ�����^�0�P��Q�M���|F>�Z���� %.Z��9��qa��{���;ٶ�7�DSll�v:��t4�N���k�j&�=#��½J��6��P��є�lIvb���:M���KE�K��/�(�؊҄y~������O=��G�����V?��<�7�� 3M�N���^�+ٮy�ݵ�� �Fq��nmL�Y�輽�p-1�+��<��WѶ�P�F�o�T��9���o�Ҕ��B؛ӰR�7�a98f=6�q{?-�����\�V�ZeLN���Id.gF�1*WJ��x%���3�^|�~���-�f��W!<�3��x�8i���h��>j������*��=��Ea�f�ι
�R�w�����/
������vJ�t:�Y�v����ۚ���4�F�|h��ģ���FJ!$�L��˾�Q�6i���F��j��S��Y��rvA��S2�G���όܥɔ�v��]z������o�tb 3+
��ǡ��;$�z�U���.�V��K]�$Jӻ�>�Z	���IQ�@��v��Y�+�X�{5j�t�S:�Y�ںQ,ٕ_���B4VA/)m"&�i[�rJa����d���� ����]���h����b�l1�ny?fq�J��޴_�]䴻/i���"�-�t ԖC�A$���{ErB�*.l�3/��d�sv�����B����z)=7��+�]�<�Ґӿ�^D�h�L���҆��p<�Y���o���O*����77B���8V�XGBY���X� ^�ퟟUk�E�Rl�� 4�R������OTH7��Zv�I-��/�֫�G�����?�$�A^ʞ��wJ�A�B؄Ba^���F#^�I��MB-����U�.;I*�*�"S7��Y�v����31c�&#�yB�����[h;��
��N�����\�h�F�����g��j���ȘsR�H�'�O�B�ޚ`�J���n.��Ϡ���,�~�*���N),-1��c��9��������~B�;?ӹiŗ������4q)���[�o#^r+|��C�pV��.]��jg�Sm(��?A�'?�B���e�������q�m^�xu��:e���k�C} 4��aMGO�b�]��Cƃq�CF-�믽��y��(s�F����;i�#̀hY�2�?���_�A��^�;����j����l	.B�
w)<��]www�[�����

�@�P�s���}q��t_̟����b�%�Q�eӞ;�'q��+�_B�Ē�Q�\>�0��o3��{����|���|�.`x�N^������S�V]����<��R��������	
�`dqe��<O�i �dOSVV���!v�
@A���)HZ�8��B?�T�zY
�$P%�m�)k
���ӂ��lx�	eT�M(r�g�n�5ﾯ��|���'��%C��y�Σ�`����ے�ړ����OB�j�]6^*+��d�a9�VU]h�`��-Nv-�e���C%��Z1�2 T���sQ�ٱ�z��k[� ��`��6x.r�V���<����3��.G��S��(�)	>O�.�������s���Wן�o��;��>}!)�I����F�r��A�HC|����&��G����`�|����w�J�̱�V����Ĺ3�X��&�x=�e�igÛ��#a<(�Y�����������H��=�C�\���8�����3KoC��N����(m��	��&_Ȳ�V6u^E=ۄH�dj�T�}��Q��1�+���,6�d�'�1�e����]����0����LiX�> i	Qv�Z	��%sbq�¾ɮW{Z��>qo$8ْ��f{)dA"'���ϽD}�3���7t��߯4����Qӯ�/�^�겋��D;��pf��2���SE�a�����bV�\��(DV߸\O���B'6Z)���-����u�P��_U�yeL�d���5I�q�#r<DQ�'��^�`�=���������@GB���:�$FC�T7���b�1W.�4F�)'Z�	����沧N�*T��Ó��7��py�L�ԭ(�����8��-8N�N��.�GU�瞿���M���>j�]6�������*��y�����Y={�˸S��_"T=֛��i�K����/@6&�>�v�!}��L/|퐬���Y�qq�H�4 �f=
�9.S�� �q�nH�ޔn�ԟn���=Ŏ�������-J[+_�v�A�����}�R~�'����|��gUnhn~H���i��MgF5S��vVK-HT��m�<i�ހ��۬�,e}.�:7��OM�H��MF��h󉨓����яٻG��/)���P�=�z8�%�V��*��MCFU��ed?-�5�k9��.e\��E��#ΰ��(߹N@(���E���o��[.�ڽ>̍��ց���Z{Y��:��s���5��r�EK���R�|9����}�A� ���BXe�m&Ξ�?N�б�U�ܸ�4�/�N�h���d���b1�xQ�c7*�6.6�̽�q�e� �^�z�PX��*a5�|�J@�:����W�g�h���R!ƻ�X�>>�U?��G?�K����[-�n'�J��1�`�m.���w�;�H����g0�֡��5��M]hsMZ �֔��ju���ah���������k�<+b�=�jq�� �X �k���<4�M�����-�pa�/+4�u)O����K��X�)9a�6� `�$+���~On��RI��N[Ɉ��"���+�gq3y��r%�S`+�����zD�E�a�y�Y�t���C�S� ̽}i�q���֤�Y��ϫU�3���fD-�*�Ga��Ɏ�����ڔ���Mm���y�
BZs�ȣiu:S������^X�E @Gh(S MUȏb���6��'��8B���3������O�Z�';%e�z�������.�V�)�o��>>��4����D����s�҂��b֞�}9�>�u#���ե\�������|�'_1U(���D�t1�n�]� ^�s�d)�����p'�L9�Ad�r��L�q���P���9�O���~y�P�c���b��?���M�j�.������i�m��D���[\o�2- �$�[��L����|�Z)�ӥ�r�qTh�f$d<s''�{�Pj�IqvwR�A�Ƞ��7v����2�@�ջB������c~��Ui&�j��6�͝�h��P�@*�U����E���T"�V�4�y���z�vư~��==�(����i���a$-��G{�on�Y������)�n��G<�0�6
` ��Q�۔տÿ�$��U.%/��e��e��fv�7.d�'����"W)3?=-%���A����Մ�<�Y�#4��,�ZlZ=�	��Ϡm]�z�]A�B������}�1�<Yg͜��"A�!�SE��2�����m�(��'.��G�Lމ��?�͍��KC^ɠ�'��07��%�]�G�F��<��|�{�L��TSu'�������`#�������1˾ZY�&8In0�r�V������^�O�+�`�!���|� c���岄b���撃2&\�6��xe�S�?)y.5�$ZS�-�E&�ǅ,"��#�0�}��X�v<	���뎰To��7Ga��j��[EX���"�2��'�[�S��A�����X�as#煮,f���v
x��Y��>�Y���\i]��J(�i���.<�,���M�śd����!/N�G�	&�F�D�]y����.�n=Y��� �����.n'��;�k�	6��]&#h���8���X^���/����i����g�>\;�v���,�����_��U�Ř��XpN}bHV������Cvq���m��YIra��9��.'*����[���Ӕٻ;�\�D�(�uޒ�N��?!���P6^{��ynOOc*���6��.�H�uPT�I�d�e	w�m��Br>�X4���ə��k:���b�!v�w8I��$�z�4���.3���j|-Y�2˞�l�_���T����Ae�a��y�/%�~�r��u�v��
�f+`Py�.$�B��a��8i6��<ZLf��hƋ�,[�oe�<����:��//���&`��ڿ�e�+���"�Gɇ�1?�����C�=�K�j"k�,vg'�.k	���q8sWN������I��1V��� ��W�	��W����Ws:��m�{Җ}�9[4�\��y����_[x��C�������ǳ��F^�b�JF�|��3%0^��	 >�j�gB��I�X����dr�^8ka�īxr��E��Z`�y��(�L�ٔUq��Z���Nf�LN���[��#wݐޢ��%�r� ��'����N��.�9�ݩP\��[߈i�q���5p�������%=6�G��W�P�Y��L������勇����:�ߘ���&ˤ�^3�H/��������~�@i�v�y���$n��_�����6ǎ��Nb&Q��m;r8:�5�<�����>"v�\���_t�tT]q/��E[匀��q��5-K�c�Y�c�ㅙnRi�4�y����Y�s�;	>N��}�"��j�Lk�紴�QRm�3�}�ݳ�@��D��{z�G�V���Z׺x]Yv#���3�?&�n�*�\y'������vn����l����D�Q�9͊O������4�2���q��\�٩�j�+Q��F@�Y��������iL��C�}��
�f}�*�5�'��?�=đ�F���������jW��������f����~�t�2��K�������4)�gE����r]��k.��BAwS$�nr�S��s �e�o����u�/��pq?�+G;�&wv�����d�֨F>l���P�VV�S�6�؞��Gx�>��Hxּ�^err�'���lq/�����Y������I�X���he�e|��	�o�|}Z���� %j�����G`����ix���;�J\;��x�+�x�t��-���-����51V�j=�/���g���xo�G��<�%���9�C%��z��do�<w���0��']	�&M=�g��I��3�T_��X�Mww�*�Q�4�x�/�)ֺ?i�?U�P�_#�=�~Jo��sH�ypM��?�7 ���TMd9�?�2�� ��T=YJ�Bg�5z\���3c�v��=�y��t@�.�ގ�q�K�#��-WP颃���lT���� L�*EQ]x_�}�X04>`׺tEVGWڂ���c�ze�ۤ`IߵM,�8����'���@H�����t*m�^��mɖ�1�t�X� B�n�8���i�j�U�O�����m�Aq����ISH6�H��R߶�����#��OA�9Z��Fl1���b�(�ek3䛂)�c~5U&Ѕ�����~�ȓ�Q����2>��
���EZ䲺;~�����LE��ا�[�Q�̕�@��m-���0^	sH���󢹀+Оyns�Xh21p�B��p��Q�l��h�k��Y���;l���9_��|<x�Z�0t��%3�����|���)4x���q���+#хCzS4���b0D�%��B)?q�ϊ8I.!k��3�����a�WRo_DD�44�J���~E��.^�_�a��c�.l�jT�r֪�F��go�}Xlq$��g-j�-?��l�L g� ��&�Q�>8�|d�*159�y�c*��`��5V�T�ޣp�џ
��]�QB��o���4K���P�J!���q���d��qu�E�wU��N�rw�gI6ޖ�j}U��vvl�~�'��}�J9�����s��C&{�K�H����C��;�١�!�������y}iL�\��6�ī��E�`�1	T��p�h��,g�K�5p�0(����f�њ�M�wh;������+a�
�f��-ĿN�'zr�Q��*X�ˬ�J"1�3r@���ސl���޾��r<�֋:͛�>*��z��@b��v����z"Hom�qW�?$�UGԺ$q�ȱO` B���IY�B��_g�̩��L�1�R��8B �Q�U<�	گXt��8��.�3�<��N���҂�9���IFg\�4�W$Ò���<�����������T�5M�_ʎ�e1Vi�<���o/��y�H��.G�b������]�{`0��k/>�KYM�g��n}�xЪ����"E�{����E'��i�g=��I_���cs�p� u��q�	���%�2?���#� ����ĳ�'.�� 7�b`ǳ������6C��H	�;#���1,��C�(�=(`�w����-�++e1i���%��o�Y?��}���}?_�6�WS�fO��s��#2=^A��J��Ј� e����V�{rI�7�<~���
�����5����]Sm ;�^E=9���;J�5�M�|J�� ��cY`�Ie�C������(0�[Q�wnU����i2r0�	����G"��"�d_���gx�\k˒�*�#c�n�/s�D��#�H���Й>�j��&0'40�����L�aq��=�ץ[�3����[�䅶�q�+j���M��}Np)B�2��c-c�\,�b�F�i.�����-��WH
 >�.,�gQƭ-�	��Qs�Q�GךA�u�f6��$��e��Bm��wC�_~M�\��&��&�Hr�֠>�6�=��޿�:x��N]�mS�z/ҡz&}�i�?�7옷-���4Ys֮m�.�em�1�ś�L$�(Q2>����'�l�00W���\���4�>��,�p�X�\WK�<��w��0����&�z�b0F;;Ӊ�;���(������<�dv���U0&XR��6��;vF	��.��#<[d>&�֕��
.�8���"���̣�︴�u#�>Jr�^NYq�ۆ�"�k�h�v��N����r����~I�h@{��l/���u�򈽁�R
��p��mD}1�+M
K���HRJ���T�H���ڱ�)0�u�݁N�y$t��c��q� 99<1�Mb��3�k�N��NA�Mg���=���G�����G�4%�í�e0K��p�dS��K�5�L����qm�>r�����<��N޲�]`;L'Yq��{���\x@^�vy������pټ�D.U� ��0FM��Q�� },-�˷H_N5#4�}e�I
��]��kKY��k�v�a��|2гD[�/�⧮f?.��F�+�6mت�l�q��G`��F������z4Z��ʊS�Ĉ^n�6�y�uY��Jo�|6A�]��N�����%/e�&�6�R�4�ֈS�8i[���?&$!�Cp�"�${%?#�5Z��?�� ʠ�U�=��&��[���ȇf1#�c��x�M�	��*8��|[ົd���1�<e����#��1��r� Nq��fLH"�ݞK�W?�m��q��bX'�DG��K���}q�J)�e�]�B���oӸu�`�0���Òiӓ`����gHc=�N:��D҈�Q���Uה��Ʉ������x�}�R�-YָU���Aj�C�����rd&$��2�G�o�s�t�;�|�D�a�kG�r���7��,���)��-4nku��<���4n��� K�`R�&�?��䱢���\���U�3�doLB������P��8B��u��$Dl�OS�j�QK�b�[��^��=a��.�]/,$c�!�?���q%�������b�U3���"�=s�
�ԛ�Č������Ѵ�ኸN����iNo��~A.�s�6�C�l�Q���}����\�^g�b�6�=��D�4��U�j�j�vi���\��>��N�����O �+�</�F�?�Dz�}R`7�(.U���R�[���7�����us�eY�9�>��U0A�ϡXP�6�CW=/�8%��@��oqS��_\�|F�k��o��:~{��_0�Z��{����J� ��� �&��'Li/�������F�D�٪�U�,:w���Đ��B��X+�t�lE�=Z�\�=Ь����r�#`B�N7Ӷ����`m�3|�F�V�KB��k°|�� 1�>l�sTl��ڜNm�Ǵ`σ��A�[A����ƙ��Y.���7�����ܰg�l�"�V10×��T��^��+vϷ�o�3'�A�=��I�k�����ք3v�U
n����C�;1QX�0�.����\�H�?�W��$�n�U0�4�˸�:_S��1�5�f���%M��5ճ�x�$�z0��^�H^�7\T�uq�ӻG�5WX{��Nb���6�F�pʗ����A\1\8weO�k ߗDp�%�|`����S.���]݊��:�5�;����X�(����|u#�;�'�%�����G7�$
_2��,�2���l� �R��N���+�c�b���D��sj�5JI5P��k�$�n}�SJ�~��> ~�	
	R��K)Y�^�'wFьN��=�x��O�DD}�����Ig�v'F���q'��W���W�2E9j��-�>h��b�˩�;�葵����1��,�q��}#�.��A.G��.�"�1���^5t�G�a�r.�LE䫨�c��ecz_1� �òe:��}��a������C����$Q��N�b-ϑA��©�q���X�WN�;�cJ���!<:j�°�SNl�t�/�d�p#���;Ș��:"�~w�}��_������AG7��E#^j��82��e��`�h����I���t�*�"��`���P$������߬��a��W�{K?���"�QN3ul �?,3�s�Z�e0�'�������~+1�; �`3�H �n ������мU+����v�V�/��fX����EQ�^4�
��ƅ����T��K�^al}ϛv`:��5�yL�I(v�їt,v������l��8����/�Y^q������j�,�9��vڍÆ����C#'l��gk���/߮�� \�(P<�鋕V�A���~�7�<C��ʛ/rV�`i�ﻠF�c�j���xy|>m�J����e�g����ve�&��G<h�:f�}
�(����y�ׯ����'��4����:\C.6]˨T-Hw��y��-��K��	8�/��g�F�i�q=���.���+B1vn?�w�B�8&I^4�͔�S�c!s^*�`ӓ�5����tSx[Dm}B{uc�춾�P�P�^�Dy������wŮ���%�ӣ'A��φ�:}ϡ�1w�C���*�v�6��9�<#!e*�V*q�7>&r���6�
���qks#֒w�K�
ķC�`�g�O��|_7��Ļ[=��e��y7b�?�=��q�"$L�ߵ��`-0v��q�yARH+�*���ծ4Kső�;䕎1j;��p��7<LQ����(�5FW��*�޹.eb��RXk
@uXp8;�9�7%A^�����1|�;��E����3�s䢄�AЏ�>B��Vq�����]��q^��{���`C�y�\(?��k��j�аz4�(Ҥd� Ƶ��l%C�k�GY��]��H��&"J.��p{�pot^�@{�<�r=�n�a������jV����Ɋt�v�����!�[7�
�iH�;fc ����YV��Q�)����J�������?�iG��6cD�����7�����I:��㋸��X<��w��.P���+/[�Dz�qn=�j�X@�y�	u�LR�r���\��ڮbƯ�K�	�q�Xhw �IV@n�^�I�P��>]�nAi��I���a�t8Q"���SR�1 ��R�̤kaf��~�G.������IFhΰ�K���{��V&EW�%'�&ۼ�K�E(��[��!����G��N�M^<���.�⦵����.��+�7��&�kA�?���4�*�!�v/���i�$���K��v ��Z~|Z���荕�u�e�WU5�B��Qux�5?��+���%��@�VY�VP߱�-�e�ʆ�xR�ȗY�F����+�u$��N!�g�Ⴆj}�����}��5a���<rDyx�����~�k�l> ߴp����\(��Q1��� 0?����}�h���Ω���I6X3Eu_����#Q%�M+�<����\HED�Z?�`r��Y�eJ�2��?�3�Y}hp�߅��D��*X���>>���-XY
�CF�q�X�&l8�|�+i��Q��D��'�/Ŝ+ n��<��C�-��M� u����K�59�2�#��맦����)SF��	�g&�Wt}�I9sj�uV>�Q%[�9�V�3���$T�J��s�^�CXD���%�ڜ_�X7�q�<�N�Ѩ�	�q�]���z�btD]�YJ�zƟ��lna%Uف�� l��)���i]�'�}O�D������`M�lҶ'Q��:A:9���(A��A-�#���!�s{��7�e�����=F��Tؕ#T��u$�6�A�4^�,�=���n89F7�J�N�W�lے����wM���!*��>}����d�&I%z<_��e	N����	..� i���άuG�:!� ���M�tkQ�UjwdK�}��짦��P��F8������~bD"V��\	y����ݳe�Y> R~��A}6�Kr��7�㦗�Wr�s��~:��z�k9���g�;L'���=����a �x)��F$^-��.^�M�p�AP��r Н.����|�=ֳ��e�g-ym�
�ݼ�nK�jO!;��W����?:���ܶO��d��Om7zn�+G3�*k=C��n���y�o��h���{1��v�O�9#���Ô{������-�,hl�ڤ̉��t������M^��ֲrW�Vb�� ��~C*�䤤�qڶ�b|�]��_��%�Vh�Q����5��He,�}"ͤ�v���p%a{����ǣ���-�)J�jSb�*��f���I�z'�	�~w�n�h���b���n���H8���IH�{��R�E�t�ϾJ2U�f1���P��^��i��8� �dR�c�ɇ��z;o����-ǃZU�Cĩ#Dvy��X	��5I�,�/YL������ ˤQ	b\����e���n�%��f~}�\���=΁�S�4�$+�$����Nwz�����#4��o�����!q*�w�Q�B՞܍�1cN�u��־>;F�� p1�[��Ɗ�㳨�Ԅ�K�>�,�@����Z�yEu�~ڥ#� ,��5#���g�;�d�]�Z��"kn�]��`�M�W���SL��������&�)*/683��AG��q�����2�����4uXP����dM��a�O�1�d�4䡕��`���A�`�c����<���w�u��@��W&����/�(
�?��1���'�dQ�,���Y7e�܂ٸ����B�6W�*��6p��L�)v�y�ң�|����2"���g�\춽y��ܛ�N)�7�{):��i�nϣ*���h�K+T�,����~E��B�qA@L�:_Z�Tޛ8NbJj�}���>j�/�P��`m�i�&}q�(3�mc�<p��!s�F�s�+3�m�����\]f=9:�"��$�Ml�;�]�b��>��o4e���J����tZ�i6P�"�`���H��Zʹ��5�a/�U���W���3�bL�@��4�d}oJɋ��?&��M�õ�C����t��'x~��, ��r'v�Ab�'������1��^!m�ow�4e����Oa�JK,���I��-��	��1�>�ں΅�J��%&#�Y�}�0V1`����(��DV�Р����� 	;��!�FO~���S���~��֍y�X,��&�+#Dt�I_����g����s�Iĝ��(*�"��B��ٲ��|ù�}�2̟ ۠�sKX1t@�����џR�az(�8
�O���sS�`��ߜ�{0k�6D��5�ev�i��[6̎��RX�tڍI�pmͪ�C�Kbb�Ə@gv9�IA��m�����"F�~mw���֏�=mW'���>Z
L|���I� ���o��b�
^r�6}m��3����C!�ӡ�<�Դ���>H9G$/T��JDJ-�뚣�a�_�0�d� ����7 �u޻�����u��"c|��R�R�~���S��دh��_׃4�
�l���l>&@�;���H}�<�R _��-r�2M��3����8-�@���F����܋�la�u
���y��7��j�t����*5���*�����?_��է'���;�bW�a�2^�^�i��C뙢�"�n'�έPOq4.�c|��<AB8A�K`�; *��ty�s[����ٹ����\ ��3�ܨ`��Q��3t�C��F�I{�.�������Nh4��������g�W���F���]r�Ps�����]�EPl������d?t����yv����[~�J���s�Y�Y�����ʱ�D� �X�-/j�|���I�T��{�v����<~\r�s b;K�N� ���a#�)re�>��Dlghx��i�V�`\����m�<*��x5��$;��)���7Kx����h�]	��ᑥ��l,i�Ȕ�@��e��gӎ�d�<�0Z���iM
�TP�Eg���Fa q��:�62�4��v	��RA<��4��.N&ަ�����|��-1�P��Ix��>��V��K�Pƛn����}�H�/N�'{���鍭&#Xݡ��F���7�u8��vC��8�mWW��I[�P�ݩ|�0(���`ӭ�sjD��E�����X�������]-��=}o ��H�ݻ]Î1��a�����{�=����yȎ���n��{q5 2�ep!���"�f�Ч/�ҙDR3C��=�E����W�.Ŷ����䘒�ˣ�e�j�Ͽd�G���tc}�G$��5�����_�L_���,(A##�����	�a�:W�GC��}�^�;���pi�d���>��hLp�*�&�1�2���{��g��f{���,ݔ��K*�:5��V�"&���	���{�����+<=q����t�R����r��";ͺ����A}���Є�3g�|��X_6�arQ�|%��-Ϥ?��L^H�ȐcA��=l��9����sCF���R N��,�WՉ)Cy�A%��=��}��(��#��&�]{���y� W��o�(
��	�=�ޚ��h�?���xƾR�캏����� n��^X��i��T�����G�g�I	��O�9I���~�AU1����� ���qo���P.�s�X����A�M�� "�Г�����@��Ղ��=�f�5���c�+<I��� Pz���G��&t���&�]�����kaw�m�:/w�̀M 9HM�^[K$��;'�5Յ�o&|�k�Y���=M��P��O�#��;�mըl�b�
c�6ȟ�3e'�eSfo�X���}�p{��-c�%%����'������$�!�<{�Cۏ�ٔSv��mIx� � �g�u�KN�4�r���-�Y{#��Z�ᑨ�+C�F^��u�!s8�Q����q< E.H�cK��n#��uY�#�߹�G���"���O��
I�MV�����X�a��x�1��|�kC��6�w�͚��+	e��P�D���]}(4��3��o���k�'��n{��N5ÃK�$'-�ݗ�a���D�Y�ԑ������y�jH4XWm*X�����=��@��s�M�C��`�Ue�`�i�mI�Tu]��CDAk�KA���1�,�K���ސ���RQO3�臎aңg6��zڛJ�r�cF�ş�5q	y`�?ߐ!�:�4#�鱝������P��q�G�z��Ɨ9!	?(3����Q����sH9a��9��y����)yEs^�%+T�\��*�9ѯj�n���)��:�̯��v7��!	��[0	X�;p����FK�m���Me��֕y�
n�c#��]�r` 1�W�+�|�R�,2���G_���ƫ6���N��jJ��F ��W���`�q���%�V��pɓ*4&��n���'$�Wb>hi�=Pm�P1�T6��;��g��G�8L���{�w��..&�PvV��_�Z���ކ�Sp��Y�>d�0�o� ����,�P���A7o��H��u��~	 8��o���T����gA��/�Z��?���҃�8�%����� �~{0�_%�|�Ƚ#�\��<�Oo5w�C~��(d6���G�� ,P�߳71ŴI���7����7u��� v��YNߥDс����QXB��Y���z�H���I [��m[>u +UL�e�]��c>��i��X!S7�Ym�T�uo�<��~
�Ђ�aJ��<�s3�t��Բ,Z�{��iF��j��Ěi�y9蚻x=,��Eu��W{Z�$�G�F�g�����aNB�����`Ѷ��=N2���%�( �U��Fj���>|��<���F�'��|��@=�O�*�b��N�=PD�~���}��%o�vK� ��-~ĩ�S���qR�Y�m���l�-���:�Z-�����%���N��.'��n�?��4%��Q���7��'��Z[������+��T!�8�!�DN��{g�[�or�\S��5Ikk|q[�Ƚp�&U�ޯB�wz%(��cUྭ�?PK   �X�X�BI9�  �  /   images/fec15d42-0ad5-4a5a-b895-65211c19e81b.png�T�[��D6�E`"��"C��5��ب�%�!�N�c�tLB�A������'�{��{�~�.�X���� �XC]Y������?����3|uco�}�G�'���JZ#����>�V^v����Nn.�6Vv��^�g�td��
zy�f.�K���BlY&q�)��:*c�'�֯=8)�])�
����@�>b�Jj�WjE�Ő�T�IG�\�x��.{�q��T�t8�k�*ki��뀲L�dd^t	5y�'�KOQ�
Iy��N�O�,��S���� G��A'�ǽ��ĈL���_�A?@�6���dܐ��|������%������M?���P�3#����Hq�M��
\�ϗS�-������H^�?Ŏ6��v=0�������>5���*�R����J�y5�(B>�~�/�u�n���]����[>t���`D<9"3F�%��`�o����[-��bZ���T��$���A�3Y��-�.L���=k�4Ĺ}�M(,� ������k]@M�\J���}
yxi��W�p�� �Xp��̈����ߥ��ݏ6�j�OI�����R�c�M���*��wa�����ѭ[�]��G$��Hc���E���`��O�t[�h��5�aP���Q�4\�9����XMj�6��:�i���z0_��7��Yv~�۷xH��P%>�5q��]j�K(�O�R塗bd��]�I���B)��*fՍ��y��E�t���4���c��p%�6A\n��b��k�ut�G�!N�3�C	�}��2H[3ݮ����F>�lfg�6.�v���Z�ܔ��y}\V�?6Y�Z�Y���->�[|;B���~d}R�0F۷���C��K+P/>����?��Q�eaM�1Z#�s�K#�4�ޅR�m��Vl�݂0s�< 	*[��D:�pp�ar=A���g̍_b
���]<��g��3�����G����xܔ�)�����zP���mb�J�{-75�I�!��g�h�ZT9GLTP��
=��gk�a�����?f��P���s|�b���+�Ɍ�n:�X��~�P�>M��{L��L�˂��'2	�m��]�jJ0 )�LRL,�U_�l�M�q������:�oçS�u�zi�:FF �O�z�i���P}�
��_Qr���$҈�����F\0�@���m���$]8W�V���G>�\L*���S #Q�Z�R�٩�nt��V�H��J�[i� �I�fD�F�DD��ϑ�7K��B�H��[�5_�oS����K��'}�FG�~����Z�2t�om��N$c[�A�O����wG��$H����j�%4��*����@b<��6�Ոt$X��W���}GG�K�E��~��Ct/8z�
�+"4�;��y�[L.��r�Z��6�jJK}�rbuCxP�)�lZ$�[&k���\x����Ĝ
��im�QE�Pa�!���y� jWj$�[�ѴM��u+b2B6��l��K$`6&������r�j#^NxI_z�g��H[%�g��8���y�]����f�c��57����|�y�!��x�]���WZ-�YG�l�*��#?��Ι��F3��Y'�T5[�q��Ķ�r�+�6��	n�,��7<�)�r#e:�$"�������umn�ns�?R��y�Qs'�F��;���i��X��ic^f4�j�L�.��+oM��I�B[N������X�J��M9[��-�$z�[����V�6/�+txB���-�t����_���y˼D[J�T&c�;�t�o?c,��8W"����}x�$Ifa	d"W�("�#����eG��) 4��������{��b���)�)�M��*�:��A�v��*ݞ�E��Na���	E�ε`K�\tC~ep`L��My�B���kr72HM�E��oC �<DJ�'<���rOS�r�;�/%]fU���)/	�=mD A~p+ �5>5�����D	8Kz#q�w����ɤ[�Ŏ�j0�u!pGf`W^]f}��6X���$\�u�#}��<A=DĤo�uC���"�`�z��22���.Ö�L'��~�b}�0�S�-�뗅z���4{��0���}�
��}-샡���W��0�X���0>-2hټ-� �X&�}p�mL z�E��[@8��E��Nr��N��am�an`��s`����w�����(33�gE���[�����l�)(�T=Y�*��0��\�c�Н�dr!m��R�k	�������Fְ'�G��'Ϟޅ����� DJ�w``����meӊ������ਛ�`�W�*>4�So{�ܳ��C6i��n�+��:w{��w�8�ۯs/R>�����I$���9��I�����-����O�x������]�ZJ�v�(�"�\��9�W�C�h
��{-�.;��aI= �x1�����JvXH����3r�ܩ"�-hInC����1e���I��i7���S61T�U�.n�~{�� �&m>2'�)z����4W<��m�5�3�G�	:����4�����|wH�=��.�9k4v���?1m�m2��zV�(�$��| >�R��^��S�������^<��i�;���8�3 F����lS�^>����"-�|K'�@����oҝ�^���Z5)�v�l!b����|�J+��'Di�e>ʈK�x-���g-Mb�I�W(uvq�>��/�IqI����m���D-��=��Z�w�(����wq�>��\����Wz�ԧ�Q�<?�b�����{ICcc*��S��I.E���fz� pq�޵np6h-��bJ)h�z�j�-i��˶߉�ک�LJ��}Q5T�:���e�!j���d�7�}T���
������U�	��=1jѧ�I<�m+�T/�ѹ��M|�4�ru��R����6��v3���69S����u�B��=�C�L=Ό�j�;�Ɗ1톶#,M�|��-A�W�J��nVܪ���+�0���ju'�{W<�F����z��D;��3p|pA���0'Pِ��4v������p�[�S<^��A�M� ����eu�z�t��K�(�'銗&T
?�!�P��:A�z=,�S]�����8���yM|rC|��%LA����RX�ǆ	�;���C�>����e��}��қ�:�j�?1*����\E!Z�s��[4f�ѵ5��S��˭jqi�j�is�W��B�q��k�sn�)�a48��vZU����o>ũ���X._�����ǳ>����G���:���\�E�Ww�FOTk��\=S���,���'�"��on��4��gD�GQv��+��9������fͅ&)���`�����=$�V���� �����ؾ�t	r�D(��p������YX��@&�%uN/w��Н�#��d.�o_KjŖ#����c����$��U��/U����Ks�,�-I��yTM"E���}̿�
E�G��+C����Q`���]���i:�#���}�@��
u�-ǵ�M9q3�*5TB�TjP�'��i2���g�\�8�����3����n�Hhm���!`�9��L�N�JqBuVQe=fߡp��1!	���U)��B�l���&`%�~�b�Y�g�$��4��R�̩R��������Z�%Z����$�ux^�޾A�ϽG��*P����S7�If�n��u���\���Al�^�N���q}����Z�D�e��e�-?-s���������$,��a��/���3#..�f��9��njE�Iˌ��Mzc���N`�	��m �Bڝ��oI$����[�,���"�ʲ���`+�����C�l�3d�\s��,�,rbj�����9|%�`/���T�ks�KS��3�V�⵱δ�މ�(Z�1��X� ZI��=�pp�Nj����6}��r�dΰ�d�ZSK���ɮV�(&���li~�$͘���Ν���91A�e
ۜ�u(�
d�$o���1g��⛟i!lv5��#�b�t��i�qOw���`�舾E���G�ӌ8��u���Ú�Y��Te���C�d���ùw�ZW�}�Үf�N}<Q�Mj�$[m=2�'��T,��_����ochם�	�� ӯ=i�p�b�3K�3��|"%Y:��]���b����t	u�˻��v_�]Y6��R�S�F�|�,�O�̧�3�<�P�)A�y��'+�����uZ�_���1F���:�u�7��E��nd�4�n�������v�=#Ddr����t�8?I#0�"y�.;������>�!��z?���8\�˞�+v�O���#�[�ݔd�+H�}R�v�t�8��O���V�93P�W�r�%���Sy�Ca�0��1��)�4-`��������2z�"�h���B*�۳e��Þ����Y�V�R��MZ: ��B�QwD�̲J�1��?1�\qÂ[�Mtᗇ������h.�l<{\��p�Q-�uJ_EN�	&��A�n�"�ߔ?9���hf�v�i���1�c�h��SE�$u���"�n�45��X�z���'m-���e|��Vj�"q�rE��Ns�s׭!�ix�^2)�3�����@yra/h��vJ������9͔_�>Z��If���}Ϝ�g�� ���]r��F]4}f�i�a9���xx�7k%�0����4T��u���PK   �X�X0+p�  L     jsons/user_defined.json�\�nI����f1�BfF^�f��/ܲ`�=c�W��K�K�{�A�3�Mɋ.d�,R�]�d�Ȋ��<q"2ӿ���ݥ���l����)ף���/i<��~A+Z1�2����I���_}�p��^f����5�;zgn:M�����������y0W�f)��t<K�~����;�3(�e$G�s��\k��ߤI�wӅm�/�PlM�ef1!;"�P�9��4уrL������wW�ލr��{4�}SO���f����R_����>6��w��F)����٨��-��W�q��ђ�fRC��x��J
�� $��4�����/�o^���T~O��e��\H[Q-��.=��������<������81�qs���z>���:4����,;KC$��HDԔ�d��jH&�t9����I�D�b���v���T����5�4�~Z���g}
����L{�M��S0�F(�VX���Q��E+4��d"�t��(	�Y��t:�[a�	Z�%�'�AR"��ħ�H�IZ/U�Ru��JR�Z�e+L�á�@ˊ��@�45����z$��k��*�oH'\T�q���a����։��$��H�=��l�֖	 K\��~��l:����R�ο��>��a���K4��(�
Ć�AR����<��(����*""���(�0�sk����
����QJX��@6�zDrm��	��ev�!���T����v�ᦫhe+�87�D��~�n:�ְ�F��>�Q��K�B��oF'��jT�3-��ϰ�p�eȻ
�-��j�1v�%~l���	_�i'��i��ŝ-��YZ��s�°�g�sI�ԖL{�;K�S%t猩�)ԙ�c�&L�"n��1���X/<:1�Q�TF�t�ó�'GaFn�fQqɏ�kܲJIi�@h����f6��MI�{�����0M���-"�w�Fi�����	���^#���i��/���/�$��@��(�^+�є1T��rv#C�n�9kC&i�4$�2t!VH��qvN�;�����	V2v���_ �+}�ȶ�p���Qp��:�C썕DI�X`6�W��3��*���b�rn�F� t�Y�$u������\~i�}�c������S=�=2�յq��ln�|��m��F���t6�Cs�v�޻Q��{�����$����Ƌr��b<��Y��|uv�{a0s�DM��XGÈ�R���aE�RW��:�,�%���O1|#��x��O�C��䪘�R�P,\��[�������vOM������Fn���`?^�9����|�Y�ۋ�g�����R���ه��Z���$C�I��B����c$��U���B�1$��J
E�3@ɭ�V��s�v��#.�@��������|�2#X*#9L4��L���R�Y�o�� N�9��t놩�O�vb�Z��`G4�ON,Gs�T#3�ͩY��Yg�5:�o,�Kv�Y&R�T	e�hfYh�<���E����� ���S�l aZkfUV��֕R��+=`TUZQ��a��Z�K:�;�_ǚ�g7���8l'�-逭�Ȏj淗g9�ӿ ����y�no�?��X��b����~�]��m=r����:�;1j'��-ME�2Q�:�X��ZR�1H&�2j�)n��ϊ��&7T�,�3xf:2�"yg��� �᝼�׬Wۋ\����1E.^��qN!�)d/?\���Ҳ���`t���S(P��O'�BW�Ѝ{�i8�5��d��D���)��@�]A�������ԥV�f�*�%j���6Ix�id�?��� =�荭 Q��pD��$5��T�,������Dr+Wҙ�&��kT���A�Y�d}�1b�dj
� 4�� � [��g�w����W�sp��:��&ڂ!9 	-&�yNHr�k����F'�$"x��Eg���/��B�B���A��q�x	�4/���=��7۫ؖV�E<ȁ�e�D�}e�.�mLA�S���%Y�/ȿ�8��(���'e��1{|�y{�h�� J�K1`�,�i���0��
����`�`_�W�A1�,��Y8��Zh����^&�dϗպ�պ��պ��䋟M��h^Wwn�5�F;�&p����E��n�ئ��\���5i2m��BTbX�`&���BY��l���ǵ6ms.+i1�A�p&8����(�o��R�2����\����h`�MPQ)5;H�8A�J�4ѭcԢ@�����xMX���#������ԍk�^`He��!�t9�B�t�ڱ�5�����Mr3��X�o�9Y�`t�$���f�R`(7�D���ɶ�Ǐ�9	0�qd��eAGⅰ�'�$mvԸ��#��Q1G�������`$a aB���s̎�	��<�qB+á�n�|+	�l,==@�Gz�c|���a��^=kN��*��]�6��JQ7-���lF����E<}���):{����7����THÕ�8��D�E)��(����9��B�X�&�8�8/ۧu���α5�^�Q���Ѝ��rK��@�6���:��Y��i�u��ͯ�?�f��H��ko��R����$�n����+zte�i~`W0~*}�����|�p,�VO�\����G&<��.|�7�Q� �<N�������~�s��C�E��ް��b�A�r3�^���C��Ȑ�f��ָw���2�IF�^�Ȑ�Ri��Rô�k��t��yo��J)��׭����5RP�D�����`K�,����&�2!"�s$8�>�2qT%�����g�C�Q���I��&��uS1t�.��&Z���ޥ�j�������Xc��G���	{�/�z������]2N{���l<.�p߸��+���'�樽�>��)*�\`����C0�9��1ٺ�K�N1�xEbbr,{G��D���Y���v(��Re�Z�TŁ�cv�Ҋ��"""B�݈{��j�6���x٦F)�*~p�޿{~����%(�uU���w��o?���Z}W��G{� ��%��8�8��­)
��OG@>�V���(�<h)1!x�P�tHJ'Ib����麻&8QZ�X�����@�`9��I|ՙm��u��M�n<�|z�������f�4�k?��g;�m��/c�t3e�%�{W��{�F8k����5Ճ�,��F�m�����y�b��K#������UtPb
���=#�o����0�����?�f��bt�V|~�Vl�����=/�
���o;����z�Tr�̍���&�� 1��I��H�,"4��o�ky��j.�1',IV!�����)��0K�ޏnv�z�t�����#��
&&�r;!�!y'�&`qJ���ł�^�!�Y$�"1�l���5��.���F�V'1��Zs2 g�Z������g�ŧ��C�$-�k�]����s�;˿:ȩ��|)�����S�Vt���b�b{˩��| �,���o?�tȱ *�c)�`��)�#�=��Y%��[*v`�lS �����G�}�$�]
��T#�����mQ���h  �/�o�Ʈ)`m��P��v ZU�1؇��Q�����g��ٻx�kئ��/d�r��At��o�1`l�|i`0�Kf�����ǂ�����C�>����
1���f`��),D���lӏK�A3UΈuTp��=Bϡ�=�dYb�$���?M�<f��:A *N��^�8�q~9�|�o���PK
   �X�X�,�-�  [                  cirkitFile.jsonPK
   ��X �x  ��  /             �  images/0edaf19c-8cfa-4246-aa67-58db36a161f7.pngPK
   �X�X�R�� $� /             �  images/179c08ce-6e18-4019-8002-932a24469ad1.pngPK
   �X�X��_�  >  /             Rl images/17d126d1-8a97-48c5-9cdb-beb53ba7b71c.pngPK
   �X�X����7  �  /             &� images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   �X�X�z���o U� /             �� images/3076bb86-a585-4cba-b1e7-fb1a193624b4.pngPK
   �X�X(rҪ15  ,5  /             � images/48f3676a-8ce7-4f44-9cda-e384043a380e.pngPK
   ���XdOv� +  �+  /             K= images/4b55d61a-3afb-42cc-8f41-c8483e8c29c3.pngPK
   �X�Xh`Pҷ!  �!  /             �h images/4b60cb4e-ac73-4aba-afdc-1cf5937e57a1.pngPK
   �X�Xd���Z �d /             �� images/57fbf569-4147-4eab-87dd-5f8b4e7be3fc.pngPK
   ���XvnG> �? /             ��
 images/61f4766b-b131-4d1d-b591-12c82c44e54c.pngPK
   ���X0jF6'� �� /             #$ images/6462d580-1c26-43d5-8ea3-52797bde3c40.pngPK
   �X�X�l��A Ԥ /             � images/670050b8-4f2c-4603-900e-28b8075f4ca8.pngPK
   z�X����U  8  /             �N images/68cd571a-d128-4aaf-a06e-233b43cf9b16.jpgPK
   ���X�\�#W 2Y /             �] images/72f7f29c-ad5c-43c9-9f1f-56c5e6d4e935.pngPK
   �X�X��E!  d  /             � images/73d4fb58-19c4-4d70-ae00-297313ed457a.pngPK
   �X�X�W��,  �,  /             p� images/754cf6f1-779b-4e0d-9f61-aeee66719356.pngPK
   $��X�,͓�u  sx  /             D� images/7a575584-996f-4f1b-8f01-a278e4b2f0d1.jpgPK
   �X�Xd��  �   /             ,j images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   z�X���b�  �  /             B� images/84b07818-b924-472b-989c-78bd96a030b6.jpgPK
   �X�X�ԴØ+ �{ /             �� images/85110ed8-4773-4cfe-99cf-d6f3d0ce91f3.pngPK
   ��X��x  7�  /             n� images/865a90cd-818d-4d70-9e9e-0a073e8e8390.pngPK
   ���X8Ȋܸ� �� /             �? images/88c2329a-9b4b-47e1-bc90-005d0a7e43bc.pngPK
   �X�Xmb?�4 �R /             � images/9399b738-9a99-483d-8480-139b77408719.pngPK
   �X�X�&�}[  y`  /             �J images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   ���X̜l�T~ �} /             i� images/9a4dac29-fc17-4e8f-bf63-f97779143c33.pngPK
   �X�XW���Y�   /             
%  images/a615f73c-88fd-4a5c-a08d-6962f48a0070.pngPK
   �X�X	��#u } /             ��  images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   ���Xo�Z��  �% /              a" images/bf12b6e8-34f4-4879-8616-fd29946f5bfe.pngPK
   ���XZMZ��� d� /             5�$ images/c9083cab-aae4-4f9e-a621-fba1f0ef8f4d.pngPK
   ���Xͧ��
 ܡ
 /             _|& images/d1ea3d2e-b350-4687-bed1-c7e59b56e556.pngPK
   ���XL���kB  WW  /             _1 images/e3ae6286-4af8-4c7d-b449-b4e8e59fa08a.pngPK
   �X�XA��5�)  �)  /             b1 images/f5d8cbe5-36a4-4687-b22e-186957e3c304.pngPK
   $��XK숤u  �x  /             -�1 images/f8feb36c-29ce-4e87-9091-184ea2b3473b.jpgPK
   �X�X�BI9�  �  /             2 images/fec15d42-0ad5-4a5a-b895-65211c19e81b.pngPK
   �X�X0+p�  L               2 jsons/user_defined.jsonPK    $ $ �  �#2   